module Rob(
  input         clock,
  input         reset,
  input         io_enq_valids_0,
  input  [6:0]  io_enq_uops_0_uopc,
  input  [31:0] io_enq_uops_0_inst,
  input  [31:0] io_enq_uops_0_debug_inst,
  input         io_enq_uops_0_is_rvc,
  input  [39:0] io_enq_uops_0_debug_pc,
  input  [2:0]  io_enq_uops_0_iq_type,
  input  [9:0]  io_enq_uops_0_fu_code,
  input  [3:0]  io_enq_uops_0_ctrl_br_type,
  input  [1:0]  io_enq_uops_0_ctrl_op1_sel,
  input  [2:0]  io_enq_uops_0_ctrl_op2_sel,
  input  [2:0]  io_enq_uops_0_ctrl_imm_sel,
  input  [3:0]  io_enq_uops_0_ctrl_op_fcn,
  input         io_enq_uops_0_ctrl_fcn_dw,
  input  [2:0]  io_enq_uops_0_ctrl_csr_cmd,
  input         io_enq_uops_0_ctrl_is_load,
  input         io_enq_uops_0_ctrl_is_sta,
  input         io_enq_uops_0_ctrl_is_std,
  input  [1:0]  io_enq_uops_0_iw_state,
  input         io_enq_uops_0_iw_p1_poisoned,
  input         io_enq_uops_0_iw_p2_poisoned,
  input         io_enq_uops_0_is_br,
  input         io_enq_uops_0_is_jalr,
  input         io_enq_uops_0_is_jal,
  input         io_enq_uops_0_is_sfb,
  input  [7:0]  io_enq_uops_0_br_mask,
  input  [2:0]  io_enq_uops_0_br_tag,
  input  [3:0]  io_enq_uops_0_ftq_idx,
  input         io_enq_uops_0_edge_inst,
  input  [5:0]  io_enq_uops_0_pc_lob,
  input         io_enq_uops_0_taken,
  input  [19:0] io_enq_uops_0_imm_packed,
  input  [11:0] io_enq_uops_0_csr_addr,
  input  [4:0]  io_enq_uops_0_rob_idx,
  input  [2:0]  io_enq_uops_0_ldq_idx,
  input  [2:0]  io_enq_uops_0_stq_idx,
  input  [1:0]  io_enq_uops_0_rxq_idx,
  input  [5:0]  io_enq_uops_0_pdst,
  input  [5:0]  io_enq_uops_0_prs1,
  input  [5:0]  io_enq_uops_0_prs2,
  input  [5:0]  io_enq_uops_0_prs3,
  input  [3:0]  io_enq_uops_0_ppred,
  input         io_enq_uops_0_prs1_busy,
  input         io_enq_uops_0_prs2_busy,
  input         io_enq_uops_0_prs3_busy,
  input         io_enq_uops_0_ppred_busy,
  input  [5:0]  io_enq_uops_0_stale_pdst,
  input         io_enq_uops_0_exception,
  input  [63:0] io_enq_uops_0_exc_cause,
  input         io_enq_uops_0_bypassable,
  input  [4:0]  io_enq_uops_0_mem_cmd,
  input  [1:0]  io_enq_uops_0_mem_size,
  input         io_enq_uops_0_mem_signed,
  input         io_enq_uops_0_is_fence,
  input         io_enq_uops_0_is_fencei,
  input         io_enq_uops_0_is_amo,
  input         io_enq_uops_0_uses_ldq,
  input         io_enq_uops_0_uses_stq,
  input         io_enq_uops_0_is_sys_pc2epc,
  input         io_enq_uops_0_is_unique,
  input         io_enq_uops_0_flush_on_commit,
  input         io_enq_uops_0_ldst_is_rs1,
  input  [5:0]  io_enq_uops_0_ldst,
  input  [5:0]  io_enq_uops_0_lrs1,
  input  [5:0]  io_enq_uops_0_lrs2,
  input  [5:0]  io_enq_uops_0_lrs3,
  input         io_enq_uops_0_ldst_val,
  input  [1:0]  io_enq_uops_0_dst_rtype,
  input  [1:0]  io_enq_uops_0_lrs1_rtype,
  input  [1:0]  io_enq_uops_0_lrs2_rtype,
  input         io_enq_uops_0_frs3_en,
  input         io_enq_uops_0_fp_val,
  input         io_enq_uops_0_fp_single,
  input         io_enq_uops_0_xcpt_pf_if,
  input         io_enq_uops_0_xcpt_ae_if,
  input         io_enq_uops_0_xcpt_ma_if,
  input         io_enq_uops_0_bp_debug_if,
  input         io_enq_uops_0_bp_xcpt_if,
  input  [1:0]  io_enq_uops_0_debug_fsrc,
  input  [1:0]  io_enq_uops_0_debug_tsrc,
  input         io_enq_partial_stall,
  input  [39:0] io_xcpt_fetch_pc,
  output [4:0]  io_rob_tail_idx,
  output [4:0]  io_rob_pnr_idx,
  output [4:0]  io_rob_head_idx,
  input  [7:0]  io_brupdate_b1_resolve_mask,
  input  [7:0]  io_brupdate_b1_mispredict_mask,
  input  [6:0]  io_brupdate_b2_uop_uopc,
  input  [31:0] io_brupdate_b2_uop_inst,
  input  [31:0] io_brupdate_b2_uop_debug_inst,
  input         io_brupdate_b2_uop_is_rvc,
  input  [39:0] io_brupdate_b2_uop_debug_pc,
  input  [2:0]  io_brupdate_b2_uop_iq_type,
  input  [9:0]  io_brupdate_b2_uop_fu_code,
  input  [3:0]  io_brupdate_b2_uop_ctrl_br_type,
  input  [1:0]  io_brupdate_b2_uop_ctrl_op1_sel,
  input  [2:0]  io_brupdate_b2_uop_ctrl_op2_sel,
  input  [2:0]  io_brupdate_b2_uop_ctrl_imm_sel,
  input  [3:0]  io_brupdate_b2_uop_ctrl_op_fcn,
  input         io_brupdate_b2_uop_ctrl_fcn_dw,
  input  [2:0]  io_brupdate_b2_uop_ctrl_csr_cmd,
  input         io_brupdate_b2_uop_ctrl_is_load,
  input         io_brupdate_b2_uop_ctrl_is_sta,
  input         io_brupdate_b2_uop_ctrl_is_std,
  input  [1:0]  io_brupdate_b2_uop_iw_state,
  input         io_brupdate_b2_uop_iw_p1_poisoned,
  input         io_brupdate_b2_uop_iw_p2_poisoned,
  input         io_brupdate_b2_uop_is_br,
  input         io_brupdate_b2_uop_is_jalr,
  input         io_brupdate_b2_uop_is_jal,
  input         io_brupdate_b2_uop_is_sfb,
  input  [7:0]  io_brupdate_b2_uop_br_mask,
  input  [2:0]  io_brupdate_b2_uop_br_tag,
  input  [3:0]  io_brupdate_b2_uop_ftq_idx,
  input         io_brupdate_b2_uop_edge_inst,
  input  [5:0]  io_brupdate_b2_uop_pc_lob,
  input         io_brupdate_b2_uop_taken,
  input  [19:0] io_brupdate_b2_uop_imm_packed,
  input  [11:0] io_brupdate_b2_uop_csr_addr,
  input  [4:0]  io_brupdate_b2_uop_rob_idx,
  input  [2:0]  io_brupdate_b2_uop_ldq_idx,
  input  [2:0]  io_brupdate_b2_uop_stq_idx,
  input  [1:0]  io_brupdate_b2_uop_rxq_idx,
  input  [5:0]  io_brupdate_b2_uop_pdst,
  input  [5:0]  io_brupdate_b2_uop_prs1,
  input  [5:0]  io_brupdate_b2_uop_prs2,
  input  [5:0]  io_brupdate_b2_uop_prs3,
  input  [3:0]  io_brupdate_b2_uop_ppred,
  input         io_brupdate_b2_uop_prs1_busy,
  input         io_brupdate_b2_uop_prs2_busy,
  input         io_brupdate_b2_uop_prs3_busy,
  input         io_brupdate_b2_uop_ppred_busy,
  input  [5:0]  io_brupdate_b2_uop_stale_pdst,
  input         io_brupdate_b2_uop_exception,
  input  [63:0] io_brupdate_b2_uop_exc_cause,
  input         io_brupdate_b2_uop_bypassable,
  input  [4:0]  io_brupdate_b2_uop_mem_cmd,
  input  [1:0]  io_brupdate_b2_uop_mem_size,
  input         io_brupdate_b2_uop_mem_signed,
  input         io_brupdate_b2_uop_is_fence,
  input         io_brupdate_b2_uop_is_fencei,
  input         io_brupdate_b2_uop_is_amo,
  input         io_brupdate_b2_uop_uses_ldq,
  input         io_brupdate_b2_uop_uses_stq,
  input         io_brupdate_b2_uop_is_sys_pc2epc,
  input         io_brupdate_b2_uop_is_unique,
  input         io_brupdate_b2_uop_flush_on_commit,
  input         io_brupdate_b2_uop_ldst_is_rs1,
  input  [5:0]  io_brupdate_b2_uop_ldst,
  input  [5:0]  io_brupdate_b2_uop_lrs1,
  input  [5:0]  io_brupdate_b2_uop_lrs2,
  input  [5:0]  io_brupdate_b2_uop_lrs3,
  input         io_brupdate_b2_uop_ldst_val,
  input  [1:0]  io_brupdate_b2_uop_dst_rtype,
  input  [1:0]  io_brupdate_b2_uop_lrs1_rtype,
  input  [1:0]  io_brupdate_b2_uop_lrs2_rtype,
  input         io_brupdate_b2_uop_frs3_en,
  input         io_brupdate_b2_uop_fp_val,
  input         io_brupdate_b2_uop_fp_single,
  input         io_brupdate_b2_uop_xcpt_pf_if,
  input         io_brupdate_b2_uop_xcpt_ae_if,
  input         io_brupdate_b2_uop_xcpt_ma_if,
  input         io_brupdate_b2_uop_bp_debug_if,
  input         io_brupdate_b2_uop_bp_xcpt_if,
  input  [1:0]  io_brupdate_b2_uop_debug_fsrc,
  input  [1:0]  io_brupdate_b2_uop_debug_tsrc,
  input         io_brupdate_b2_valid,
  input         io_brupdate_b2_mispredict,
  input         io_brupdate_b2_taken,
  input  [2:0]  io_brupdate_b2_cfi_type,
  input  [1:0]  io_brupdate_b2_pc_sel,
  input  [39:0] io_brupdate_b2_jalr_target,
  input         io_brupdate_b2_target_offset,
  input         io_wb_resps_0_valid,
  input  [6:0]  io_wb_resps_0_bits_uop_uopc,
  input  [31:0] io_wb_resps_0_bits_uop_inst,
  input  [31:0] io_wb_resps_0_bits_uop_debug_inst,
  input         io_wb_resps_0_bits_uop_is_rvc,
  input  [39:0] io_wb_resps_0_bits_uop_debug_pc,
  input  [2:0]  io_wb_resps_0_bits_uop_iq_type,
  input  [9:0]  io_wb_resps_0_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_0_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_0_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_0_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_wb_resps_0_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_0_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_0_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_wb_resps_0_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_0_bits_uop_ctrl_is_load,
  input         io_wb_resps_0_bits_uop_ctrl_is_sta,
  input         io_wb_resps_0_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_0_bits_uop_iw_state,
  input         io_wb_resps_0_bits_uop_iw_p1_poisoned,
  input         io_wb_resps_0_bits_uop_iw_p2_poisoned,
  input         io_wb_resps_0_bits_uop_is_br,
  input         io_wb_resps_0_bits_uop_is_jalr,
  input         io_wb_resps_0_bits_uop_is_jal,
  input         io_wb_resps_0_bits_uop_is_sfb,
  input  [7:0]  io_wb_resps_0_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_0_bits_uop_br_tag,
  input  [3:0]  io_wb_resps_0_bits_uop_ftq_idx,
  input         io_wb_resps_0_bits_uop_edge_inst,
  input  [5:0]  io_wb_resps_0_bits_uop_pc_lob,
  input         io_wb_resps_0_bits_uop_taken,
  input  [19:0] io_wb_resps_0_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_0_bits_uop_csr_addr,
  input  [4:0]  io_wb_resps_0_bits_uop_rob_idx,
  input  [2:0]  io_wb_resps_0_bits_uop_ldq_idx,
  input  [2:0]  io_wb_resps_0_bits_uop_stq_idx,
  input  [1:0]  io_wb_resps_0_bits_uop_rxq_idx,
  input  [5:0]  io_wb_resps_0_bits_uop_pdst,
  input  [5:0]  io_wb_resps_0_bits_uop_prs1,
  input  [5:0]  io_wb_resps_0_bits_uop_prs2,
  input  [5:0]  io_wb_resps_0_bits_uop_prs3,
  input  [3:0]  io_wb_resps_0_bits_uop_ppred,
  input         io_wb_resps_0_bits_uop_prs1_busy,
  input         io_wb_resps_0_bits_uop_prs2_busy,
  input         io_wb_resps_0_bits_uop_prs3_busy,
  input         io_wb_resps_0_bits_uop_ppred_busy,
  input  [5:0]  io_wb_resps_0_bits_uop_stale_pdst,
  input         io_wb_resps_0_bits_uop_exception,
  input  [63:0] io_wb_resps_0_bits_uop_exc_cause,
  input         io_wb_resps_0_bits_uop_bypassable,
  input  [4:0]  io_wb_resps_0_bits_uop_mem_cmd,
  input  [1:0]  io_wb_resps_0_bits_uop_mem_size,
  input         io_wb_resps_0_bits_uop_mem_signed,
  input         io_wb_resps_0_bits_uop_is_fence,
  input         io_wb_resps_0_bits_uop_is_fencei,
  input         io_wb_resps_0_bits_uop_is_amo,
  input         io_wb_resps_0_bits_uop_uses_ldq,
  input         io_wb_resps_0_bits_uop_uses_stq,
  input         io_wb_resps_0_bits_uop_is_sys_pc2epc,
  input         io_wb_resps_0_bits_uop_is_unique,
  input         io_wb_resps_0_bits_uop_flush_on_commit,
  input         io_wb_resps_0_bits_uop_ldst_is_rs1,
  input  [5:0]  io_wb_resps_0_bits_uop_ldst,
  input  [5:0]  io_wb_resps_0_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_0_bits_uop_lrs2,
  input  [5:0]  io_wb_resps_0_bits_uop_lrs3,
  input         io_wb_resps_0_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_0_bits_uop_dst_rtype,
  input  [1:0]  io_wb_resps_0_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_0_bits_uop_lrs2_rtype,
  input         io_wb_resps_0_bits_uop_frs3_en,
  input         io_wb_resps_0_bits_uop_fp_val,
  input         io_wb_resps_0_bits_uop_fp_single,
  input         io_wb_resps_0_bits_uop_xcpt_pf_if,
  input         io_wb_resps_0_bits_uop_xcpt_ae_if,
  input         io_wb_resps_0_bits_uop_xcpt_ma_if,
  input         io_wb_resps_0_bits_uop_bp_debug_if,
  input         io_wb_resps_0_bits_uop_bp_xcpt_if,
  input  [1:0]  io_wb_resps_0_bits_uop_debug_fsrc,
  input  [1:0]  io_wb_resps_0_bits_uop_debug_tsrc,
  input  [64:0] io_wb_resps_0_bits_data,
  input         io_wb_resps_0_bits_predicated,
  input         io_wb_resps_0_bits_fflags_valid,
  input  [6:0]  io_wb_resps_0_bits_fflags_bits_uop_uopc,
  input  [31:0] io_wb_resps_0_bits_fflags_bits_uop_inst,
  input  [31:0] io_wb_resps_0_bits_fflags_bits_uop_debug_inst,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_rvc,
  input  [39:0] io_wb_resps_0_bits_fflags_bits_uop_debug_pc,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_iq_type,
  input  [9:0]  io_wb_resps_0_bits_fflags_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_0_bits_fflags_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_0_bits_fflags_bits_uop_ctrl_is_load,
  input         io_wb_resps_0_bits_fflags_bits_uop_ctrl_is_sta,
  input         io_wb_resps_0_bits_fflags_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_iw_state,
  input         io_wb_resps_0_bits_fflags_bits_uop_iw_p1_poisoned,
  input         io_wb_resps_0_bits_fflags_bits_uop_iw_p2_poisoned,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_br,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_jalr,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_jal,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_sfb,
  input  [7:0]  io_wb_resps_0_bits_fflags_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_br_tag,
  input  [3:0]  io_wb_resps_0_bits_fflags_bits_uop_ftq_idx,
  input         io_wb_resps_0_bits_fflags_bits_uop_edge_inst,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_pc_lob,
  input         io_wb_resps_0_bits_fflags_bits_uop_taken,
  input  [19:0] io_wb_resps_0_bits_fflags_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_0_bits_fflags_bits_uop_csr_addr,
  input  [4:0]  io_wb_resps_0_bits_fflags_bits_uop_rob_idx,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_ldq_idx,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_stq_idx,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_rxq_idx,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_pdst,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_prs1,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_prs2,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_prs3,
  input  [3:0]  io_wb_resps_0_bits_fflags_bits_uop_ppred,
  input         io_wb_resps_0_bits_fflags_bits_uop_prs1_busy,
  input         io_wb_resps_0_bits_fflags_bits_uop_prs2_busy,
  input         io_wb_resps_0_bits_fflags_bits_uop_prs3_busy,
  input         io_wb_resps_0_bits_fflags_bits_uop_ppred_busy,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_stale_pdst,
  input         io_wb_resps_0_bits_fflags_bits_uop_exception,
  input  [63:0] io_wb_resps_0_bits_fflags_bits_uop_exc_cause,
  input         io_wb_resps_0_bits_fflags_bits_uop_bypassable,
  input  [4:0]  io_wb_resps_0_bits_fflags_bits_uop_mem_cmd,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_mem_size,
  input         io_wb_resps_0_bits_fflags_bits_uop_mem_signed,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_fence,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_fencei,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_amo,
  input         io_wb_resps_0_bits_fflags_bits_uop_uses_ldq,
  input         io_wb_resps_0_bits_fflags_bits_uop_uses_stq,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_sys_pc2epc,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_unique,
  input         io_wb_resps_0_bits_fflags_bits_uop_flush_on_commit,
  input         io_wb_resps_0_bits_fflags_bits_uop_ldst_is_rs1,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_ldst,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_lrs2,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_lrs3,
  input         io_wb_resps_0_bits_fflags_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_dst_rtype,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_lrs2_rtype,
  input         io_wb_resps_0_bits_fflags_bits_uop_frs3_en,
  input         io_wb_resps_0_bits_fflags_bits_uop_fp_val,
  input         io_wb_resps_0_bits_fflags_bits_uop_fp_single,
  input         io_wb_resps_0_bits_fflags_bits_uop_xcpt_pf_if,
  input         io_wb_resps_0_bits_fflags_bits_uop_xcpt_ae_if,
  input         io_wb_resps_0_bits_fflags_bits_uop_xcpt_ma_if,
  input         io_wb_resps_0_bits_fflags_bits_uop_bp_debug_if,
  input         io_wb_resps_0_bits_fflags_bits_uop_bp_xcpt_if,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_debug_fsrc,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_debug_tsrc,
  input  [4:0]  io_wb_resps_0_bits_fflags_bits_flags,
  input         io_wb_resps_1_valid,
  input  [6:0]  io_wb_resps_1_bits_uop_uopc,
  input  [31:0] io_wb_resps_1_bits_uop_inst,
  input  [31:0] io_wb_resps_1_bits_uop_debug_inst,
  input         io_wb_resps_1_bits_uop_is_rvc,
  input  [39:0] io_wb_resps_1_bits_uop_debug_pc,
  input  [2:0]  io_wb_resps_1_bits_uop_iq_type,
  input  [9:0]  io_wb_resps_1_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_1_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_1_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_1_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_wb_resps_1_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_1_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_1_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_wb_resps_1_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_1_bits_uop_ctrl_is_load,
  input         io_wb_resps_1_bits_uop_ctrl_is_sta,
  input         io_wb_resps_1_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_1_bits_uop_iw_state,
  input         io_wb_resps_1_bits_uop_iw_p1_poisoned,
  input         io_wb_resps_1_bits_uop_iw_p2_poisoned,
  input         io_wb_resps_1_bits_uop_is_br,
  input         io_wb_resps_1_bits_uop_is_jalr,
  input         io_wb_resps_1_bits_uop_is_jal,
  input         io_wb_resps_1_bits_uop_is_sfb,
  input  [7:0]  io_wb_resps_1_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_1_bits_uop_br_tag,
  input  [3:0]  io_wb_resps_1_bits_uop_ftq_idx,
  input         io_wb_resps_1_bits_uop_edge_inst,
  input  [5:0]  io_wb_resps_1_bits_uop_pc_lob,
  input         io_wb_resps_1_bits_uop_taken,
  input  [19:0] io_wb_resps_1_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_1_bits_uop_csr_addr,
  input  [4:0]  io_wb_resps_1_bits_uop_rob_idx,
  input  [2:0]  io_wb_resps_1_bits_uop_ldq_idx,
  input  [2:0]  io_wb_resps_1_bits_uop_stq_idx,
  input  [1:0]  io_wb_resps_1_bits_uop_rxq_idx,
  input  [5:0]  io_wb_resps_1_bits_uop_pdst,
  input  [5:0]  io_wb_resps_1_bits_uop_prs1,
  input  [5:0]  io_wb_resps_1_bits_uop_prs2,
  input  [5:0]  io_wb_resps_1_bits_uop_prs3,
  input  [3:0]  io_wb_resps_1_bits_uop_ppred,
  input         io_wb_resps_1_bits_uop_prs1_busy,
  input         io_wb_resps_1_bits_uop_prs2_busy,
  input         io_wb_resps_1_bits_uop_prs3_busy,
  input         io_wb_resps_1_bits_uop_ppred_busy,
  input  [5:0]  io_wb_resps_1_bits_uop_stale_pdst,
  input         io_wb_resps_1_bits_uop_exception,
  input  [63:0] io_wb_resps_1_bits_uop_exc_cause,
  input         io_wb_resps_1_bits_uop_bypassable,
  input  [4:0]  io_wb_resps_1_bits_uop_mem_cmd,
  input  [1:0]  io_wb_resps_1_bits_uop_mem_size,
  input         io_wb_resps_1_bits_uop_mem_signed,
  input         io_wb_resps_1_bits_uop_is_fence,
  input         io_wb_resps_1_bits_uop_is_fencei,
  input         io_wb_resps_1_bits_uop_is_amo,
  input         io_wb_resps_1_bits_uop_uses_ldq,
  input         io_wb_resps_1_bits_uop_uses_stq,
  input         io_wb_resps_1_bits_uop_is_sys_pc2epc,
  input         io_wb_resps_1_bits_uop_is_unique,
  input         io_wb_resps_1_bits_uop_flush_on_commit,
  input         io_wb_resps_1_bits_uop_ldst_is_rs1,
  input  [5:0]  io_wb_resps_1_bits_uop_ldst,
  input  [5:0]  io_wb_resps_1_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_1_bits_uop_lrs2,
  input  [5:0]  io_wb_resps_1_bits_uop_lrs3,
  input         io_wb_resps_1_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_1_bits_uop_dst_rtype,
  input  [1:0]  io_wb_resps_1_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_1_bits_uop_lrs2_rtype,
  input         io_wb_resps_1_bits_uop_frs3_en,
  input         io_wb_resps_1_bits_uop_fp_val,
  input         io_wb_resps_1_bits_uop_fp_single,
  input         io_wb_resps_1_bits_uop_xcpt_pf_if,
  input         io_wb_resps_1_bits_uop_xcpt_ae_if,
  input         io_wb_resps_1_bits_uop_xcpt_ma_if,
  input         io_wb_resps_1_bits_uop_bp_debug_if,
  input         io_wb_resps_1_bits_uop_bp_xcpt_if,
  input  [1:0]  io_wb_resps_1_bits_uop_debug_fsrc,
  input  [1:0]  io_wb_resps_1_bits_uop_debug_tsrc,
  input  [64:0] io_wb_resps_1_bits_data,
  input         io_wb_resps_1_bits_predicated,
  input         io_wb_resps_1_bits_fflags_valid,
  input  [6:0]  io_wb_resps_1_bits_fflags_bits_uop_uopc,
  input  [31:0] io_wb_resps_1_bits_fflags_bits_uop_inst,
  input  [31:0] io_wb_resps_1_bits_fflags_bits_uop_debug_inst,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_rvc,
  input  [39:0] io_wb_resps_1_bits_fflags_bits_uop_debug_pc,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_iq_type,
  input  [9:0]  io_wb_resps_1_bits_fflags_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_1_bits_fflags_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_1_bits_fflags_bits_uop_ctrl_is_load,
  input         io_wb_resps_1_bits_fflags_bits_uop_ctrl_is_sta,
  input         io_wb_resps_1_bits_fflags_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_iw_state,
  input         io_wb_resps_1_bits_fflags_bits_uop_iw_p1_poisoned,
  input         io_wb_resps_1_bits_fflags_bits_uop_iw_p2_poisoned,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_br,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_jalr,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_jal,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_sfb,
  input  [7:0]  io_wb_resps_1_bits_fflags_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_br_tag,
  input  [3:0]  io_wb_resps_1_bits_fflags_bits_uop_ftq_idx,
  input         io_wb_resps_1_bits_fflags_bits_uop_edge_inst,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_pc_lob,
  input         io_wb_resps_1_bits_fflags_bits_uop_taken,
  input  [19:0] io_wb_resps_1_bits_fflags_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_1_bits_fflags_bits_uop_csr_addr,
  input  [4:0]  io_wb_resps_1_bits_fflags_bits_uop_rob_idx,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_ldq_idx,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_stq_idx,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_rxq_idx,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_pdst,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_prs1,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_prs2,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_prs3,
  input  [3:0]  io_wb_resps_1_bits_fflags_bits_uop_ppred,
  input         io_wb_resps_1_bits_fflags_bits_uop_prs1_busy,
  input         io_wb_resps_1_bits_fflags_bits_uop_prs2_busy,
  input         io_wb_resps_1_bits_fflags_bits_uop_prs3_busy,
  input         io_wb_resps_1_bits_fflags_bits_uop_ppred_busy,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_stale_pdst,
  input         io_wb_resps_1_bits_fflags_bits_uop_exception,
  input  [63:0] io_wb_resps_1_bits_fflags_bits_uop_exc_cause,
  input         io_wb_resps_1_bits_fflags_bits_uop_bypassable,
  input  [4:0]  io_wb_resps_1_bits_fflags_bits_uop_mem_cmd,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_mem_size,
  input         io_wb_resps_1_bits_fflags_bits_uop_mem_signed,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_fence,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_fencei,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_amo,
  input         io_wb_resps_1_bits_fflags_bits_uop_uses_ldq,
  input         io_wb_resps_1_bits_fflags_bits_uop_uses_stq,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_sys_pc2epc,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_unique,
  input         io_wb_resps_1_bits_fflags_bits_uop_flush_on_commit,
  input         io_wb_resps_1_bits_fflags_bits_uop_ldst_is_rs1,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_ldst,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_lrs2,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_lrs3,
  input         io_wb_resps_1_bits_fflags_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_dst_rtype,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_lrs2_rtype,
  input         io_wb_resps_1_bits_fflags_bits_uop_frs3_en,
  input         io_wb_resps_1_bits_fflags_bits_uop_fp_val,
  input         io_wb_resps_1_bits_fflags_bits_uop_fp_single,
  input         io_wb_resps_1_bits_fflags_bits_uop_xcpt_pf_if,
  input         io_wb_resps_1_bits_fflags_bits_uop_xcpt_ae_if,
  input         io_wb_resps_1_bits_fflags_bits_uop_xcpt_ma_if,
  input         io_wb_resps_1_bits_fflags_bits_uop_bp_debug_if,
  input         io_wb_resps_1_bits_fflags_bits_uop_bp_xcpt_if,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_debug_fsrc,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_debug_tsrc,
  input  [4:0]  io_wb_resps_1_bits_fflags_bits_flags,
  input         io_wb_resps_2_valid,
  input  [6:0]  io_wb_resps_2_bits_uop_uopc,
  input  [31:0] io_wb_resps_2_bits_uop_inst,
  input  [31:0] io_wb_resps_2_bits_uop_debug_inst,
  input         io_wb_resps_2_bits_uop_is_rvc,
  input  [39:0] io_wb_resps_2_bits_uop_debug_pc,
  input  [2:0]  io_wb_resps_2_bits_uop_iq_type,
  input  [9:0]  io_wb_resps_2_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_2_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_2_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_2_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_wb_resps_2_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_2_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_2_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_wb_resps_2_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_2_bits_uop_ctrl_is_load,
  input         io_wb_resps_2_bits_uop_ctrl_is_sta,
  input         io_wb_resps_2_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_2_bits_uop_iw_state,
  input         io_wb_resps_2_bits_uop_iw_p1_poisoned,
  input         io_wb_resps_2_bits_uop_iw_p2_poisoned,
  input         io_wb_resps_2_bits_uop_is_br,
  input         io_wb_resps_2_bits_uop_is_jalr,
  input         io_wb_resps_2_bits_uop_is_jal,
  input         io_wb_resps_2_bits_uop_is_sfb,
  input  [7:0]  io_wb_resps_2_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_2_bits_uop_br_tag,
  input  [3:0]  io_wb_resps_2_bits_uop_ftq_idx,
  input         io_wb_resps_2_bits_uop_edge_inst,
  input  [5:0]  io_wb_resps_2_bits_uop_pc_lob,
  input         io_wb_resps_2_bits_uop_taken,
  input  [19:0] io_wb_resps_2_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_2_bits_uop_csr_addr,
  input  [4:0]  io_wb_resps_2_bits_uop_rob_idx,
  input  [2:0]  io_wb_resps_2_bits_uop_ldq_idx,
  input  [2:0]  io_wb_resps_2_bits_uop_stq_idx,
  input  [1:0]  io_wb_resps_2_bits_uop_rxq_idx,
  input  [5:0]  io_wb_resps_2_bits_uop_pdst,
  input  [5:0]  io_wb_resps_2_bits_uop_prs1,
  input  [5:0]  io_wb_resps_2_bits_uop_prs2,
  input  [5:0]  io_wb_resps_2_bits_uop_prs3,
  input  [3:0]  io_wb_resps_2_bits_uop_ppred,
  input         io_wb_resps_2_bits_uop_prs1_busy,
  input         io_wb_resps_2_bits_uop_prs2_busy,
  input         io_wb_resps_2_bits_uop_prs3_busy,
  input         io_wb_resps_2_bits_uop_ppred_busy,
  input  [5:0]  io_wb_resps_2_bits_uop_stale_pdst,
  input         io_wb_resps_2_bits_uop_exception,
  input  [63:0] io_wb_resps_2_bits_uop_exc_cause,
  input         io_wb_resps_2_bits_uop_bypassable,
  input  [4:0]  io_wb_resps_2_bits_uop_mem_cmd,
  input  [1:0]  io_wb_resps_2_bits_uop_mem_size,
  input         io_wb_resps_2_bits_uop_mem_signed,
  input         io_wb_resps_2_bits_uop_is_fence,
  input         io_wb_resps_2_bits_uop_is_fencei,
  input         io_wb_resps_2_bits_uop_is_amo,
  input         io_wb_resps_2_bits_uop_uses_ldq,
  input         io_wb_resps_2_bits_uop_uses_stq,
  input         io_wb_resps_2_bits_uop_is_sys_pc2epc,
  input         io_wb_resps_2_bits_uop_is_unique,
  input         io_wb_resps_2_bits_uop_flush_on_commit,
  input         io_wb_resps_2_bits_uop_ldst_is_rs1,
  input  [5:0]  io_wb_resps_2_bits_uop_ldst,
  input  [5:0]  io_wb_resps_2_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_2_bits_uop_lrs2,
  input  [5:0]  io_wb_resps_2_bits_uop_lrs3,
  input         io_wb_resps_2_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_2_bits_uop_dst_rtype,
  input  [1:0]  io_wb_resps_2_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_2_bits_uop_lrs2_rtype,
  input         io_wb_resps_2_bits_uop_frs3_en,
  input         io_wb_resps_2_bits_uop_fp_val,
  input         io_wb_resps_2_bits_uop_fp_single,
  input         io_wb_resps_2_bits_uop_xcpt_pf_if,
  input         io_wb_resps_2_bits_uop_xcpt_ae_if,
  input         io_wb_resps_2_bits_uop_xcpt_ma_if,
  input         io_wb_resps_2_bits_uop_bp_debug_if,
  input         io_wb_resps_2_bits_uop_bp_xcpt_if,
  input  [1:0]  io_wb_resps_2_bits_uop_debug_fsrc,
  input  [1:0]  io_wb_resps_2_bits_uop_debug_tsrc,
  input  [64:0] io_wb_resps_2_bits_data,
  input         io_wb_resps_2_bits_predicated,
  input         io_wb_resps_2_bits_fflags_valid,
  input  [6:0]  io_wb_resps_2_bits_fflags_bits_uop_uopc,
  input  [31:0] io_wb_resps_2_bits_fflags_bits_uop_inst,
  input  [31:0] io_wb_resps_2_bits_fflags_bits_uop_debug_inst,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_rvc,
  input  [39:0] io_wb_resps_2_bits_fflags_bits_uop_debug_pc,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_iq_type,
  input  [9:0]  io_wb_resps_2_bits_fflags_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_2_bits_fflags_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_2_bits_fflags_bits_uop_ctrl_is_load,
  input         io_wb_resps_2_bits_fflags_bits_uop_ctrl_is_sta,
  input         io_wb_resps_2_bits_fflags_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_iw_state,
  input         io_wb_resps_2_bits_fflags_bits_uop_iw_p1_poisoned,
  input         io_wb_resps_2_bits_fflags_bits_uop_iw_p2_poisoned,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_br,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_jalr,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_jal,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_sfb,
  input  [7:0]  io_wb_resps_2_bits_fflags_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_br_tag,
  input  [3:0]  io_wb_resps_2_bits_fflags_bits_uop_ftq_idx,
  input         io_wb_resps_2_bits_fflags_bits_uop_edge_inst,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_pc_lob,
  input         io_wb_resps_2_bits_fflags_bits_uop_taken,
  input  [19:0] io_wb_resps_2_bits_fflags_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_2_bits_fflags_bits_uop_csr_addr,
  input  [4:0]  io_wb_resps_2_bits_fflags_bits_uop_rob_idx,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_ldq_idx,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_stq_idx,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_rxq_idx,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_pdst,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_prs1,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_prs2,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_prs3,
  input  [3:0]  io_wb_resps_2_bits_fflags_bits_uop_ppred,
  input         io_wb_resps_2_bits_fflags_bits_uop_prs1_busy,
  input         io_wb_resps_2_bits_fflags_bits_uop_prs2_busy,
  input         io_wb_resps_2_bits_fflags_bits_uop_prs3_busy,
  input         io_wb_resps_2_bits_fflags_bits_uop_ppred_busy,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_stale_pdst,
  input         io_wb_resps_2_bits_fflags_bits_uop_exception,
  input  [63:0] io_wb_resps_2_bits_fflags_bits_uop_exc_cause,
  input         io_wb_resps_2_bits_fflags_bits_uop_bypassable,
  input  [4:0]  io_wb_resps_2_bits_fflags_bits_uop_mem_cmd,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_mem_size,
  input         io_wb_resps_2_bits_fflags_bits_uop_mem_signed,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_fence,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_fencei,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_amo,
  input         io_wb_resps_2_bits_fflags_bits_uop_uses_ldq,
  input         io_wb_resps_2_bits_fflags_bits_uop_uses_stq,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_sys_pc2epc,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_unique,
  input         io_wb_resps_2_bits_fflags_bits_uop_flush_on_commit,
  input         io_wb_resps_2_bits_fflags_bits_uop_ldst_is_rs1,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_ldst,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_lrs2,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_lrs3,
  input         io_wb_resps_2_bits_fflags_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_dst_rtype,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_lrs2_rtype,
  input         io_wb_resps_2_bits_fflags_bits_uop_frs3_en,
  input         io_wb_resps_2_bits_fflags_bits_uop_fp_val,
  input         io_wb_resps_2_bits_fflags_bits_uop_fp_single,
  input         io_wb_resps_2_bits_fflags_bits_uop_xcpt_pf_if,
  input         io_wb_resps_2_bits_fflags_bits_uop_xcpt_ae_if,
  input         io_wb_resps_2_bits_fflags_bits_uop_xcpt_ma_if,
  input         io_wb_resps_2_bits_fflags_bits_uop_bp_debug_if,
  input         io_wb_resps_2_bits_fflags_bits_uop_bp_xcpt_if,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_debug_fsrc,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_debug_tsrc,
  input  [4:0]  io_wb_resps_2_bits_fflags_bits_flags,
  input         io_wb_resps_3_valid,
  input  [6:0]  io_wb_resps_3_bits_uop_uopc,
  input  [31:0] io_wb_resps_3_bits_uop_inst,
  input  [31:0] io_wb_resps_3_bits_uop_debug_inst,
  input         io_wb_resps_3_bits_uop_is_rvc,
  input  [39:0] io_wb_resps_3_bits_uop_debug_pc,
  input  [2:0]  io_wb_resps_3_bits_uop_iq_type,
  input  [9:0]  io_wb_resps_3_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_3_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_3_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_3_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_wb_resps_3_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_3_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_3_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_wb_resps_3_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_3_bits_uop_ctrl_is_load,
  input         io_wb_resps_3_bits_uop_ctrl_is_sta,
  input         io_wb_resps_3_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_3_bits_uop_iw_state,
  input         io_wb_resps_3_bits_uop_iw_p1_poisoned,
  input         io_wb_resps_3_bits_uop_iw_p2_poisoned,
  input         io_wb_resps_3_bits_uop_is_br,
  input         io_wb_resps_3_bits_uop_is_jalr,
  input         io_wb_resps_3_bits_uop_is_jal,
  input         io_wb_resps_3_bits_uop_is_sfb,
  input  [7:0]  io_wb_resps_3_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_3_bits_uop_br_tag,
  input  [3:0]  io_wb_resps_3_bits_uop_ftq_idx,
  input         io_wb_resps_3_bits_uop_edge_inst,
  input  [5:0]  io_wb_resps_3_bits_uop_pc_lob,
  input         io_wb_resps_3_bits_uop_taken,
  input  [19:0] io_wb_resps_3_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_3_bits_uop_csr_addr,
  input  [4:0]  io_wb_resps_3_bits_uop_rob_idx,
  input  [2:0]  io_wb_resps_3_bits_uop_ldq_idx,
  input  [2:0]  io_wb_resps_3_bits_uop_stq_idx,
  input  [1:0]  io_wb_resps_3_bits_uop_rxq_idx,
  input  [5:0]  io_wb_resps_3_bits_uop_pdst,
  input  [5:0]  io_wb_resps_3_bits_uop_prs1,
  input  [5:0]  io_wb_resps_3_bits_uop_prs2,
  input  [5:0]  io_wb_resps_3_bits_uop_prs3,
  input  [3:0]  io_wb_resps_3_bits_uop_ppred,
  input         io_wb_resps_3_bits_uop_prs1_busy,
  input         io_wb_resps_3_bits_uop_prs2_busy,
  input         io_wb_resps_3_bits_uop_prs3_busy,
  input         io_wb_resps_3_bits_uop_ppred_busy,
  input  [5:0]  io_wb_resps_3_bits_uop_stale_pdst,
  input         io_wb_resps_3_bits_uop_exception,
  input  [63:0] io_wb_resps_3_bits_uop_exc_cause,
  input         io_wb_resps_3_bits_uop_bypassable,
  input  [4:0]  io_wb_resps_3_bits_uop_mem_cmd,
  input  [1:0]  io_wb_resps_3_bits_uop_mem_size,
  input         io_wb_resps_3_bits_uop_mem_signed,
  input         io_wb_resps_3_bits_uop_is_fence,
  input         io_wb_resps_3_bits_uop_is_fencei,
  input         io_wb_resps_3_bits_uop_is_amo,
  input         io_wb_resps_3_bits_uop_uses_ldq,
  input         io_wb_resps_3_bits_uop_uses_stq,
  input         io_wb_resps_3_bits_uop_is_sys_pc2epc,
  input         io_wb_resps_3_bits_uop_is_unique,
  input         io_wb_resps_3_bits_uop_flush_on_commit,
  input         io_wb_resps_3_bits_uop_ldst_is_rs1,
  input  [5:0]  io_wb_resps_3_bits_uop_ldst,
  input  [5:0]  io_wb_resps_3_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_3_bits_uop_lrs2,
  input  [5:0]  io_wb_resps_3_bits_uop_lrs3,
  input         io_wb_resps_3_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_3_bits_uop_dst_rtype,
  input  [1:0]  io_wb_resps_3_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_3_bits_uop_lrs2_rtype,
  input         io_wb_resps_3_bits_uop_frs3_en,
  input         io_wb_resps_3_bits_uop_fp_val,
  input         io_wb_resps_3_bits_uop_fp_single,
  input         io_wb_resps_3_bits_uop_xcpt_pf_if,
  input         io_wb_resps_3_bits_uop_xcpt_ae_if,
  input         io_wb_resps_3_bits_uop_xcpt_ma_if,
  input         io_wb_resps_3_bits_uop_bp_debug_if,
  input         io_wb_resps_3_bits_uop_bp_xcpt_if,
  input  [1:0]  io_wb_resps_3_bits_uop_debug_fsrc,
  input  [1:0]  io_wb_resps_3_bits_uop_debug_tsrc,
  input  [64:0] io_wb_resps_3_bits_data,
  input         io_wb_resps_3_bits_predicated,
  input         io_wb_resps_3_bits_fflags_valid,
  input  [6:0]  io_wb_resps_3_bits_fflags_bits_uop_uopc,
  input  [31:0] io_wb_resps_3_bits_fflags_bits_uop_inst,
  input  [31:0] io_wb_resps_3_bits_fflags_bits_uop_debug_inst,
  input         io_wb_resps_3_bits_fflags_bits_uop_is_rvc,
  input  [39:0] io_wb_resps_3_bits_fflags_bits_uop_debug_pc,
  input  [2:0]  io_wb_resps_3_bits_fflags_bits_uop_iq_type,
  input  [9:0]  io_wb_resps_3_bits_fflags_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_3_bits_fflags_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_3_bits_fflags_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_3_bits_fflags_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_wb_resps_3_bits_fflags_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_3_bits_fflags_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_3_bits_fflags_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_wb_resps_3_bits_fflags_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_3_bits_fflags_bits_uop_ctrl_is_load,
  input         io_wb_resps_3_bits_fflags_bits_uop_ctrl_is_sta,
  input         io_wb_resps_3_bits_fflags_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_3_bits_fflags_bits_uop_iw_state,
  input         io_wb_resps_3_bits_fflags_bits_uop_iw_p1_poisoned,
  input         io_wb_resps_3_bits_fflags_bits_uop_iw_p2_poisoned,
  input         io_wb_resps_3_bits_fflags_bits_uop_is_br,
  input         io_wb_resps_3_bits_fflags_bits_uop_is_jalr,
  input         io_wb_resps_3_bits_fflags_bits_uop_is_jal,
  input         io_wb_resps_3_bits_fflags_bits_uop_is_sfb,
  input  [7:0]  io_wb_resps_3_bits_fflags_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_3_bits_fflags_bits_uop_br_tag,
  input  [3:0]  io_wb_resps_3_bits_fflags_bits_uop_ftq_idx,
  input         io_wb_resps_3_bits_fflags_bits_uop_edge_inst,
  input  [5:0]  io_wb_resps_3_bits_fflags_bits_uop_pc_lob,
  input         io_wb_resps_3_bits_fflags_bits_uop_taken,
  input  [19:0] io_wb_resps_3_bits_fflags_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_3_bits_fflags_bits_uop_csr_addr,
  input  [4:0]  io_wb_resps_3_bits_fflags_bits_uop_rob_idx,
  input  [2:0]  io_wb_resps_3_bits_fflags_bits_uop_ldq_idx,
  input  [2:0]  io_wb_resps_3_bits_fflags_bits_uop_stq_idx,
  input  [1:0]  io_wb_resps_3_bits_fflags_bits_uop_rxq_idx,
  input  [5:0]  io_wb_resps_3_bits_fflags_bits_uop_pdst,
  input  [5:0]  io_wb_resps_3_bits_fflags_bits_uop_prs1,
  input  [5:0]  io_wb_resps_3_bits_fflags_bits_uop_prs2,
  input  [5:0]  io_wb_resps_3_bits_fflags_bits_uop_prs3,
  input  [3:0]  io_wb_resps_3_bits_fflags_bits_uop_ppred,
  input         io_wb_resps_3_bits_fflags_bits_uop_prs1_busy,
  input         io_wb_resps_3_bits_fflags_bits_uop_prs2_busy,
  input         io_wb_resps_3_bits_fflags_bits_uop_prs3_busy,
  input         io_wb_resps_3_bits_fflags_bits_uop_ppred_busy,
  input  [5:0]  io_wb_resps_3_bits_fflags_bits_uop_stale_pdst,
  input         io_wb_resps_3_bits_fflags_bits_uop_exception,
  input  [63:0] io_wb_resps_3_bits_fflags_bits_uop_exc_cause,
  input         io_wb_resps_3_bits_fflags_bits_uop_bypassable,
  input  [4:0]  io_wb_resps_3_bits_fflags_bits_uop_mem_cmd,
  input  [1:0]  io_wb_resps_3_bits_fflags_bits_uop_mem_size,
  input         io_wb_resps_3_bits_fflags_bits_uop_mem_signed,
  input         io_wb_resps_3_bits_fflags_bits_uop_is_fence,
  input         io_wb_resps_3_bits_fflags_bits_uop_is_fencei,
  input         io_wb_resps_3_bits_fflags_bits_uop_is_amo,
  input         io_wb_resps_3_bits_fflags_bits_uop_uses_ldq,
  input         io_wb_resps_3_bits_fflags_bits_uop_uses_stq,
  input         io_wb_resps_3_bits_fflags_bits_uop_is_sys_pc2epc,
  input         io_wb_resps_3_bits_fflags_bits_uop_is_unique,
  input         io_wb_resps_3_bits_fflags_bits_uop_flush_on_commit,
  input         io_wb_resps_3_bits_fflags_bits_uop_ldst_is_rs1,
  input  [5:0]  io_wb_resps_3_bits_fflags_bits_uop_ldst,
  input  [5:0]  io_wb_resps_3_bits_fflags_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_3_bits_fflags_bits_uop_lrs2,
  input  [5:0]  io_wb_resps_3_bits_fflags_bits_uop_lrs3,
  input         io_wb_resps_3_bits_fflags_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_3_bits_fflags_bits_uop_dst_rtype,
  input  [1:0]  io_wb_resps_3_bits_fflags_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_3_bits_fflags_bits_uop_lrs2_rtype,
  input         io_wb_resps_3_bits_fflags_bits_uop_frs3_en,
  input         io_wb_resps_3_bits_fflags_bits_uop_fp_val,
  input         io_wb_resps_3_bits_fflags_bits_uop_fp_single,
  input         io_wb_resps_3_bits_fflags_bits_uop_xcpt_pf_if,
  input         io_wb_resps_3_bits_fflags_bits_uop_xcpt_ae_if,
  input         io_wb_resps_3_bits_fflags_bits_uop_xcpt_ma_if,
  input         io_wb_resps_3_bits_fflags_bits_uop_bp_debug_if,
  input         io_wb_resps_3_bits_fflags_bits_uop_bp_xcpt_if,
  input  [1:0]  io_wb_resps_3_bits_fflags_bits_uop_debug_fsrc,
  input  [1:0]  io_wb_resps_3_bits_fflags_bits_uop_debug_tsrc,
  input  [4:0]  io_wb_resps_3_bits_fflags_bits_flags,
  input         io_lsu_clr_bsy_0_valid,
  input  [4:0]  io_lsu_clr_bsy_0_bits,
  input         io_lsu_clr_bsy_1_valid,
  input  [4:0]  io_lsu_clr_bsy_1_bits,
  input         io_lsu_clr_unsafe_0_valid,
  input  [4:0]  io_lsu_clr_unsafe_0_bits,
  input         io_debug_wb_valids_0,
  input         io_debug_wb_valids_1,
  input         io_debug_wb_valids_2,
  input         io_debug_wb_valids_3,
  input  [63:0] io_debug_wb_wdata_0,
  input  [63:0] io_debug_wb_wdata_1,
  input  [63:0] io_debug_wb_wdata_2,
  input  [63:0] io_debug_wb_wdata_3,
  input         io_fflags_0_valid,
  input  [6:0]  io_fflags_0_bits_uop_uopc,
  input  [31:0] io_fflags_0_bits_uop_inst,
  input  [31:0] io_fflags_0_bits_uop_debug_inst,
  input         io_fflags_0_bits_uop_is_rvc,
  input  [39:0] io_fflags_0_bits_uop_debug_pc,
  input  [2:0]  io_fflags_0_bits_uop_iq_type,
  input  [9:0]  io_fflags_0_bits_uop_fu_code,
  input  [3:0]  io_fflags_0_bits_uop_ctrl_br_type,
  input  [1:0]  io_fflags_0_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_fflags_0_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_fflags_0_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_fflags_0_bits_uop_ctrl_op_fcn,
  input         io_fflags_0_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_fflags_0_bits_uop_ctrl_csr_cmd,
  input         io_fflags_0_bits_uop_ctrl_is_load,
  input         io_fflags_0_bits_uop_ctrl_is_sta,
  input         io_fflags_0_bits_uop_ctrl_is_std,
  input  [1:0]  io_fflags_0_bits_uop_iw_state,
  input         io_fflags_0_bits_uop_iw_p1_poisoned,
  input         io_fflags_0_bits_uop_iw_p2_poisoned,
  input         io_fflags_0_bits_uop_is_br,
  input         io_fflags_0_bits_uop_is_jalr,
  input         io_fflags_0_bits_uop_is_jal,
  input         io_fflags_0_bits_uop_is_sfb,
  input  [7:0]  io_fflags_0_bits_uop_br_mask,
  input  [2:0]  io_fflags_0_bits_uop_br_tag,
  input  [3:0]  io_fflags_0_bits_uop_ftq_idx,
  input         io_fflags_0_bits_uop_edge_inst,
  input  [5:0]  io_fflags_0_bits_uop_pc_lob,
  input         io_fflags_0_bits_uop_taken,
  input  [19:0] io_fflags_0_bits_uop_imm_packed,
  input  [11:0] io_fflags_0_bits_uop_csr_addr,
  input  [4:0]  io_fflags_0_bits_uop_rob_idx,
  input  [2:0]  io_fflags_0_bits_uop_ldq_idx,
  input  [2:0]  io_fflags_0_bits_uop_stq_idx,
  input  [1:0]  io_fflags_0_bits_uop_rxq_idx,
  input  [5:0]  io_fflags_0_bits_uop_pdst,
  input  [5:0]  io_fflags_0_bits_uop_prs1,
  input  [5:0]  io_fflags_0_bits_uop_prs2,
  input  [5:0]  io_fflags_0_bits_uop_prs3,
  input  [3:0]  io_fflags_0_bits_uop_ppred,
  input         io_fflags_0_bits_uop_prs1_busy,
  input         io_fflags_0_bits_uop_prs2_busy,
  input         io_fflags_0_bits_uop_prs3_busy,
  input         io_fflags_0_bits_uop_ppred_busy,
  input  [5:0]  io_fflags_0_bits_uop_stale_pdst,
  input         io_fflags_0_bits_uop_exception,
  input  [63:0] io_fflags_0_bits_uop_exc_cause,
  input         io_fflags_0_bits_uop_bypassable,
  input  [4:0]  io_fflags_0_bits_uop_mem_cmd,
  input  [1:0]  io_fflags_0_bits_uop_mem_size,
  input         io_fflags_0_bits_uop_mem_signed,
  input         io_fflags_0_bits_uop_is_fence,
  input         io_fflags_0_bits_uop_is_fencei,
  input         io_fflags_0_bits_uop_is_amo,
  input         io_fflags_0_bits_uop_uses_ldq,
  input         io_fflags_0_bits_uop_uses_stq,
  input         io_fflags_0_bits_uop_is_sys_pc2epc,
  input         io_fflags_0_bits_uop_is_unique,
  input         io_fflags_0_bits_uop_flush_on_commit,
  input         io_fflags_0_bits_uop_ldst_is_rs1,
  input  [5:0]  io_fflags_0_bits_uop_ldst,
  input  [5:0]  io_fflags_0_bits_uop_lrs1,
  input  [5:0]  io_fflags_0_bits_uop_lrs2,
  input  [5:0]  io_fflags_0_bits_uop_lrs3,
  input         io_fflags_0_bits_uop_ldst_val,
  input  [1:0]  io_fflags_0_bits_uop_dst_rtype,
  input  [1:0]  io_fflags_0_bits_uop_lrs1_rtype,
  input  [1:0]  io_fflags_0_bits_uop_lrs2_rtype,
  input         io_fflags_0_bits_uop_frs3_en,
  input         io_fflags_0_bits_uop_fp_val,
  input         io_fflags_0_bits_uop_fp_single,
  input         io_fflags_0_bits_uop_xcpt_pf_if,
  input         io_fflags_0_bits_uop_xcpt_ae_if,
  input         io_fflags_0_bits_uop_xcpt_ma_if,
  input         io_fflags_0_bits_uop_bp_debug_if,
  input         io_fflags_0_bits_uop_bp_xcpt_if,
  input  [1:0]  io_fflags_0_bits_uop_debug_fsrc,
  input  [1:0]  io_fflags_0_bits_uop_debug_tsrc,
  input  [4:0]  io_fflags_0_bits_flags,
  input         io_fflags_1_valid,
  input  [6:0]  io_fflags_1_bits_uop_uopc,
  input  [31:0] io_fflags_1_bits_uop_inst,
  input  [31:0] io_fflags_1_bits_uop_debug_inst,
  input         io_fflags_1_bits_uop_is_rvc,
  input  [39:0] io_fflags_1_bits_uop_debug_pc,
  input  [2:0]  io_fflags_1_bits_uop_iq_type,
  input  [9:0]  io_fflags_1_bits_uop_fu_code,
  input  [3:0]  io_fflags_1_bits_uop_ctrl_br_type,
  input  [1:0]  io_fflags_1_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_fflags_1_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_fflags_1_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_fflags_1_bits_uop_ctrl_op_fcn,
  input         io_fflags_1_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_fflags_1_bits_uop_ctrl_csr_cmd,
  input         io_fflags_1_bits_uop_ctrl_is_load,
  input         io_fflags_1_bits_uop_ctrl_is_sta,
  input         io_fflags_1_bits_uop_ctrl_is_std,
  input  [1:0]  io_fflags_1_bits_uop_iw_state,
  input         io_fflags_1_bits_uop_iw_p1_poisoned,
  input         io_fflags_1_bits_uop_iw_p2_poisoned,
  input         io_fflags_1_bits_uop_is_br,
  input         io_fflags_1_bits_uop_is_jalr,
  input         io_fflags_1_bits_uop_is_jal,
  input         io_fflags_1_bits_uop_is_sfb,
  input  [7:0]  io_fflags_1_bits_uop_br_mask,
  input  [2:0]  io_fflags_1_bits_uop_br_tag,
  input  [3:0]  io_fflags_1_bits_uop_ftq_idx,
  input         io_fflags_1_bits_uop_edge_inst,
  input  [5:0]  io_fflags_1_bits_uop_pc_lob,
  input         io_fflags_1_bits_uop_taken,
  input  [19:0] io_fflags_1_bits_uop_imm_packed,
  input  [11:0] io_fflags_1_bits_uop_csr_addr,
  input  [4:0]  io_fflags_1_bits_uop_rob_idx,
  input  [2:0]  io_fflags_1_bits_uop_ldq_idx,
  input  [2:0]  io_fflags_1_bits_uop_stq_idx,
  input  [1:0]  io_fflags_1_bits_uop_rxq_idx,
  input  [5:0]  io_fflags_1_bits_uop_pdst,
  input  [5:0]  io_fflags_1_bits_uop_prs1,
  input  [5:0]  io_fflags_1_bits_uop_prs2,
  input  [5:0]  io_fflags_1_bits_uop_prs3,
  input  [3:0]  io_fflags_1_bits_uop_ppred,
  input         io_fflags_1_bits_uop_prs1_busy,
  input         io_fflags_1_bits_uop_prs2_busy,
  input         io_fflags_1_bits_uop_prs3_busy,
  input         io_fflags_1_bits_uop_ppred_busy,
  input  [5:0]  io_fflags_1_bits_uop_stale_pdst,
  input         io_fflags_1_bits_uop_exception,
  input  [63:0] io_fflags_1_bits_uop_exc_cause,
  input         io_fflags_1_bits_uop_bypassable,
  input  [4:0]  io_fflags_1_bits_uop_mem_cmd,
  input  [1:0]  io_fflags_1_bits_uop_mem_size,
  input         io_fflags_1_bits_uop_mem_signed,
  input         io_fflags_1_bits_uop_is_fence,
  input         io_fflags_1_bits_uop_is_fencei,
  input         io_fflags_1_bits_uop_is_amo,
  input         io_fflags_1_bits_uop_uses_ldq,
  input         io_fflags_1_bits_uop_uses_stq,
  input         io_fflags_1_bits_uop_is_sys_pc2epc,
  input         io_fflags_1_bits_uop_is_unique,
  input         io_fflags_1_bits_uop_flush_on_commit,
  input         io_fflags_1_bits_uop_ldst_is_rs1,
  input  [5:0]  io_fflags_1_bits_uop_ldst,
  input  [5:0]  io_fflags_1_bits_uop_lrs1,
  input  [5:0]  io_fflags_1_bits_uop_lrs2,
  input  [5:0]  io_fflags_1_bits_uop_lrs3,
  input         io_fflags_1_bits_uop_ldst_val,
  input  [1:0]  io_fflags_1_bits_uop_dst_rtype,
  input  [1:0]  io_fflags_1_bits_uop_lrs1_rtype,
  input  [1:0]  io_fflags_1_bits_uop_lrs2_rtype,
  input         io_fflags_1_bits_uop_frs3_en,
  input         io_fflags_1_bits_uop_fp_val,
  input         io_fflags_1_bits_uop_fp_single,
  input         io_fflags_1_bits_uop_xcpt_pf_if,
  input         io_fflags_1_bits_uop_xcpt_ae_if,
  input         io_fflags_1_bits_uop_xcpt_ma_if,
  input         io_fflags_1_bits_uop_bp_debug_if,
  input         io_fflags_1_bits_uop_bp_xcpt_if,
  input  [1:0]  io_fflags_1_bits_uop_debug_fsrc,
  input  [1:0]  io_fflags_1_bits_uop_debug_tsrc,
  input  [4:0]  io_fflags_1_bits_flags,
  input         io_lxcpt_valid,
  input  [6:0]  io_lxcpt_bits_uop_uopc,
  input  [31:0] io_lxcpt_bits_uop_inst,
  input  [31:0] io_lxcpt_bits_uop_debug_inst,
  input         io_lxcpt_bits_uop_is_rvc,
  input  [39:0] io_lxcpt_bits_uop_debug_pc,
  input  [2:0]  io_lxcpt_bits_uop_iq_type,
  input  [9:0]  io_lxcpt_bits_uop_fu_code,
  input  [3:0]  io_lxcpt_bits_uop_ctrl_br_type,
  input  [1:0]  io_lxcpt_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_lxcpt_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_lxcpt_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_lxcpt_bits_uop_ctrl_op_fcn,
  input         io_lxcpt_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_lxcpt_bits_uop_ctrl_csr_cmd,
  input         io_lxcpt_bits_uop_ctrl_is_load,
  input         io_lxcpt_bits_uop_ctrl_is_sta,
  input         io_lxcpt_bits_uop_ctrl_is_std,
  input  [1:0]  io_lxcpt_bits_uop_iw_state,
  input         io_lxcpt_bits_uop_iw_p1_poisoned,
  input         io_lxcpt_bits_uop_iw_p2_poisoned,
  input         io_lxcpt_bits_uop_is_br,
  input         io_lxcpt_bits_uop_is_jalr,
  input         io_lxcpt_bits_uop_is_jal,
  input         io_lxcpt_bits_uop_is_sfb,
  input  [7:0]  io_lxcpt_bits_uop_br_mask,
  input  [2:0]  io_lxcpt_bits_uop_br_tag,
  input  [3:0]  io_lxcpt_bits_uop_ftq_idx,
  input         io_lxcpt_bits_uop_edge_inst,
  input  [5:0]  io_lxcpt_bits_uop_pc_lob,
  input         io_lxcpt_bits_uop_taken,
  input  [19:0] io_lxcpt_bits_uop_imm_packed,
  input  [11:0] io_lxcpt_bits_uop_csr_addr,
  input  [4:0]  io_lxcpt_bits_uop_rob_idx,
  input  [2:0]  io_lxcpt_bits_uop_ldq_idx,
  input  [2:0]  io_lxcpt_bits_uop_stq_idx,
  input  [1:0]  io_lxcpt_bits_uop_rxq_idx,
  input  [5:0]  io_lxcpt_bits_uop_pdst,
  input  [5:0]  io_lxcpt_bits_uop_prs1,
  input  [5:0]  io_lxcpt_bits_uop_prs2,
  input  [5:0]  io_lxcpt_bits_uop_prs3,
  input  [3:0]  io_lxcpt_bits_uop_ppred,
  input         io_lxcpt_bits_uop_prs1_busy,
  input         io_lxcpt_bits_uop_prs2_busy,
  input         io_lxcpt_bits_uop_prs3_busy,
  input         io_lxcpt_bits_uop_ppred_busy,
  input  [5:0]  io_lxcpt_bits_uop_stale_pdst,
  input         io_lxcpt_bits_uop_exception,
  input  [63:0] io_lxcpt_bits_uop_exc_cause,
  input         io_lxcpt_bits_uop_bypassable,
  input  [4:0]  io_lxcpt_bits_uop_mem_cmd,
  input  [1:0]  io_lxcpt_bits_uop_mem_size,
  input         io_lxcpt_bits_uop_mem_signed,
  input         io_lxcpt_bits_uop_is_fence,
  input         io_lxcpt_bits_uop_is_fencei,
  input         io_lxcpt_bits_uop_is_amo,
  input         io_lxcpt_bits_uop_uses_ldq,
  input         io_lxcpt_bits_uop_uses_stq,
  input         io_lxcpt_bits_uop_is_sys_pc2epc,
  input         io_lxcpt_bits_uop_is_unique,
  input         io_lxcpt_bits_uop_flush_on_commit,
  input         io_lxcpt_bits_uop_ldst_is_rs1,
  input  [5:0]  io_lxcpt_bits_uop_ldst,
  input  [5:0]  io_lxcpt_bits_uop_lrs1,
  input  [5:0]  io_lxcpt_bits_uop_lrs2,
  input  [5:0]  io_lxcpt_bits_uop_lrs3,
  input         io_lxcpt_bits_uop_ldst_val,
  input  [1:0]  io_lxcpt_bits_uop_dst_rtype,
  input  [1:0]  io_lxcpt_bits_uop_lrs1_rtype,
  input  [1:0]  io_lxcpt_bits_uop_lrs2_rtype,
  input         io_lxcpt_bits_uop_frs3_en,
  input         io_lxcpt_bits_uop_fp_val,
  input         io_lxcpt_bits_uop_fp_single,
  input         io_lxcpt_bits_uop_xcpt_pf_if,
  input         io_lxcpt_bits_uop_xcpt_ae_if,
  input         io_lxcpt_bits_uop_xcpt_ma_if,
  input         io_lxcpt_bits_uop_bp_debug_if,
  input         io_lxcpt_bits_uop_bp_xcpt_if,
  input  [1:0]  io_lxcpt_bits_uop_debug_fsrc,
  input  [1:0]  io_lxcpt_bits_uop_debug_tsrc,
  input  [4:0]  io_lxcpt_bits_cause,
  input  [39:0] io_lxcpt_bits_badvaddr,
  output        io_commit_valids_0,
  output        io_commit_arch_valids_0,
  output [6:0]  io_commit_uops_0_uopc,
  output [31:0] io_commit_uops_0_inst,
  output [31:0] io_commit_uops_0_debug_inst,
  output        io_commit_uops_0_is_rvc,
  output [39:0] io_commit_uops_0_debug_pc,
  output [2:0]  io_commit_uops_0_iq_type,
  output [9:0]  io_commit_uops_0_fu_code,
  output [3:0]  io_commit_uops_0_ctrl_br_type,
  output [1:0]  io_commit_uops_0_ctrl_op1_sel,
  output [2:0]  io_commit_uops_0_ctrl_op2_sel,
  output [2:0]  io_commit_uops_0_ctrl_imm_sel,
  output [3:0]  io_commit_uops_0_ctrl_op_fcn,
  output        io_commit_uops_0_ctrl_fcn_dw,
  output [2:0]  io_commit_uops_0_ctrl_csr_cmd,
  output        io_commit_uops_0_ctrl_is_load,
  output        io_commit_uops_0_ctrl_is_sta,
  output        io_commit_uops_0_ctrl_is_std,
  output [1:0]  io_commit_uops_0_iw_state,
  output        io_commit_uops_0_iw_p1_poisoned,
  output        io_commit_uops_0_iw_p2_poisoned,
  output        io_commit_uops_0_is_br,
  output        io_commit_uops_0_is_jalr,
  output        io_commit_uops_0_is_jal,
  output        io_commit_uops_0_is_sfb,
  output [7:0]  io_commit_uops_0_br_mask,
  output [2:0]  io_commit_uops_0_br_tag,
  output [3:0]  io_commit_uops_0_ftq_idx,
  output        io_commit_uops_0_edge_inst,
  output [5:0]  io_commit_uops_0_pc_lob,
  output        io_commit_uops_0_taken,
  output [19:0] io_commit_uops_0_imm_packed,
  output [11:0] io_commit_uops_0_csr_addr,
  output [4:0]  io_commit_uops_0_rob_idx,
  output [2:0]  io_commit_uops_0_ldq_idx,
  output [2:0]  io_commit_uops_0_stq_idx,
  output [1:0]  io_commit_uops_0_rxq_idx,
  output [5:0]  io_commit_uops_0_pdst,
  output [5:0]  io_commit_uops_0_prs1,
  output [5:0]  io_commit_uops_0_prs2,
  output [5:0]  io_commit_uops_0_prs3,
  output [3:0]  io_commit_uops_0_ppred,
  output        io_commit_uops_0_prs1_busy,
  output        io_commit_uops_0_prs2_busy,
  output        io_commit_uops_0_prs3_busy,
  output        io_commit_uops_0_ppred_busy,
  output [5:0]  io_commit_uops_0_stale_pdst,
  output        io_commit_uops_0_exception,
  output [63:0] io_commit_uops_0_exc_cause,
  output        io_commit_uops_0_bypassable,
  output [4:0]  io_commit_uops_0_mem_cmd,
  output [1:0]  io_commit_uops_0_mem_size,
  output        io_commit_uops_0_mem_signed,
  output        io_commit_uops_0_is_fence,
  output        io_commit_uops_0_is_fencei,
  output        io_commit_uops_0_is_amo,
  output        io_commit_uops_0_uses_ldq,
  output        io_commit_uops_0_uses_stq,
  output        io_commit_uops_0_is_sys_pc2epc,
  output        io_commit_uops_0_is_unique,
  output        io_commit_uops_0_flush_on_commit,
  output        io_commit_uops_0_ldst_is_rs1,
  output [5:0]  io_commit_uops_0_ldst,
  output [5:0]  io_commit_uops_0_lrs1,
  output [5:0]  io_commit_uops_0_lrs2,
  output [5:0]  io_commit_uops_0_lrs3,
  output        io_commit_uops_0_ldst_val,
  output [1:0]  io_commit_uops_0_dst_rtype,
  output [1:0]  io_commit_uops_0_lrs1_rtype,
  output [1:0]  io_commit_uops_0_lrs2_rtype,
  output        io_commit_uops_0_frs3_en,
  output        io_commit_uops_0_fp_val,
  output        io_commit_uops_0_fp_single,
  output        io_commit_uops_0_xcpt_pf_if,
  output        io_commit_uops_0_xcpt_ae_if,
  output        io_commit_uops_0_xcpt_ma_if,
  output        io_commit_uops_0_bp_debug_if,
  output        io_commit_uops_0_bp_xcpt_if,
  output [1:0]  io_commit_uops_0_debug_fsrc,
  output [1:0]  io_commit_uops_0_debug_tsrc,
  output        io_commit_fflags_valid,
  output [4:0]  io_commit_fflags_bits,
  output [31:0] io_commit_debug_insts_0,
  output        io_commit_rbk_valids_0,
  output        io_commit_rollback,
  output [63:0] io_commit_debug_wdata_0,
  output        io_com_load_is_at_rob_head,
  output        io_com_xcpt_valid,
  output [3:0]  io_com_xcpt_bits_ftq_idx,
  output        io_com_xcpt_bits_edge_inst,
  output        io_com_xcpt_bits_is_rvc,
  output [5:0]  io_com_xcpt_bits_pc_lob,
  output [63:0] io_com_xcpt_bits_cause,
  output [63:0] io_com_xcpt_bits_badvaddr,
  output [2:0]  io_com_xcpt_bits_flush_typ,
  input         io_csr_stall,
  output        io_flush_valid,
  output [3:0]  io_flush_bits_ftq_idx,
  output        io_flush_bits_edge_inst,
  output        io_flush_bits_is_rvc,
  output [5:0]  io_flush_bits_pc_lob,
  output [63:0] io_flush_bits_cause,
  output [63:0] io_flush_bits_badvaddr,
  output [2:0]  io_flush_bits_flush_typ,
  output        io_empty,
  output        io_ready,
  output        io_flush_frontend,
  input  [63:0] io_debug_tsc
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [63:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [63:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [63:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [63:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [63:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [63:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [63:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [63:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [63:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [63:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [63:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [63:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [63:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [63:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [63:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [63:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [63:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [63:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [63:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [63:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [63:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [63:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [63:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [63:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [63:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [63:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [63:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [63:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [63:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [63:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [63:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [63:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [63:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [63:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [63:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [63:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [63:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [31:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [63:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1725;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
  reg [63:0] _RAND_1729;
  reg [31:0] _RAND_1730;
  reg [31:0] _RAND_1731;
  reg [31:0] _RAND_1732;
  reg [31:0] _RAND_1733;
  reg [31:0] _RAND_1734;
  reg [31:0] _RAND_1735;
  reg [31:0] _RAND_1736;
  reg [31:0] _RAND_1737;
  reg [31:0] _RAND_1738;
  reg [31:0] _RAND_1739;
  reg [31:0] _RAND_1740;
  reg [31:0] _RAND_1741;
  reg [31:0] _RAND_1742;
  reg [31:0] _RAND_1743;
  reg [31:0] _RAND_1744;
  reg [31:0] _RAND_1745;
  reg [31:0] _RAND_1746;
  reg [31:0] _RAND_1747;
  reg [31:0] _RAND_1748;
  reg [31:0] _RAND_1749;
  reg [31:0] _RAND_1750;
  reg [31:0] _RAND_1751;
  reg [31:0] _RAND_1752;
  reg [31:0] _RAND_1753;
  reg [31:0] _RAND_1754;
  reg [31:0] _RAND_1755;
  reg [31:0] _RAND_1756;
  reg [31:0] _RAND_1757;
  reg [31:0] _RAND_1758;
  reg [31:0] _RAND_1759;
  reg [31:0] _RAND_1760;
  reg [31:0] _RAND_1761;
  reg [31:0] _RAND_1762;
  reg [31:0] _RAND_1763;
  reg [31:0] _RAND_1764;
  reg [31:0] _RAND_1765;
  reg [31:0] _RAND_1766;
  reg [31:0] _RAND_1767;
  reg [31:0] _RAND_1768;
  reg [31:0] _RAND_1769;
  reg [31:0] _RAND_1770;
  reg [31:0] _RAND_1771;
  reg [63:0] _RAND_1772;
  reg [31:0] _RAND_1773;
  reg [31:0] _RAND_1774;
  reg [31:0] _RAND_1775;
  reg [31:0] _RAND_1776;
  reg [31:0] _RAND_1777;
  reg [31:0] _RAND_1778;
  reg [31:0] _RAND_1779;
  reg [31:0] _RAND_1780;
  reg [31:0] _RAND_1781;
  reg [31:0] _RAND_1782;
  reg [31:0] _RAND_1783;
  reg [31:0] _RAND_1784;
  reg [31:0] _RAND_1785;
  reg [31:0] _RAND_1786;
  reg [31:0] _RAND_1787;
  reg [31:0] _RAND_1788;
  reg [31:0] _RAND_1789;
  reg [31:0] _RAND_1790;
  reg [31:0] _RAND_1791;
  reg [31:0] _RAND_1792;
  reg [31:0] _RAND_1793;
  reg [31:0] _RAND_1794;
  reg [31:0] _RAND_1795;
  reg [31:0] _RAND_1796;
  reg [31:0] _RAND_1797;
  reg [31:0] _RAND_1798;
  reg [31:0] _RAND_1799;
  reg [31:0] _RAND_1800;
  reg [31:0] _RAND_1801;
  reg [31:0] _RAND_1802;
  reg [31:0] _RAND_1803;
  reg [31:0] _RAND_1804;
  reg [31:0] _RAND_1805;
  reg [31:0] _RAND_1806;
  reg [31:0] _RAND_1807;
  reg [63:0] _RAND_1808;
  reg [31:0] _RAND_1809;
  reg [31:0] _RAND_1810;
  reg [31:0] _RAND_1811;
  reg [31:0] _RAND_1812;
  reg [31:0] _RAND_1813;
  reg [31:0] _RAND_1814;
  reg [31:0] _RAND_1815;
  reg [31:0] _RAND_1816;
  reg [31:0] _RAND_1817;
  reg [31:0] _RAND_1818;
  reg [31:0] _RAND_1819;
  reg [31:0] _RAND_1820;
  reg [31:0] _RAND_1821;
  reg [31:0] _RAND_1822;
  reg [31:0] _RAND_1823;
  reg [31:0] _RAND_1824;
  reg [31:0] _RAND_1825;
  reg [31:0] _RAND_1826;
  reg [31:0] _RAND_1827;
  reg [31:0] _RAND_1828;
  reg [31:0] _RAND_1829;
  reg [31:0] _RAND_1830;
  reg [31:0] _RAND_1831;
  reg [31:0] _RAND_1832;
  reg [31:0] _RAND_1833;
  reg [31:0] _RAND_1834;
  reg [31:0] _RAND_1835;
  reg [31:0] _RAND_1836;
  reg [31:0] _RAND_1837;
  reg [31:0] _RAND_1838;
  reg [31:0] _RAND_1839;
  reg [31:0] _RAND_1840;
  reg [31:0] _RAND_1841;
  reg [31:0] _RAND_1842;
  reg [31:0] _RAND_1843;
  reg [31:0] _RAND_1844;
  reg [31:0] _RAND_1845;
  reg [31:0] _RAND_1846;
  reg [31:0] _RAND_1847;
  reg [31:0] _RAND_1848;
  reg [31:0] _RAND_1849;
  reg [31:0] _RAND_1850;
  reg [63:0] _RAND_1851;
  reg [31:0] _RAND_1852;
  reg [31:0] _RAND_1853;
  reg [31:0] _RAND_1854;
  reg [31:0] _RAND_1855;
  reg [31:0] _RAND_1856;
  reg [31:0] _RAND_1857;
  reg [31:0] _RAND_1858;
  reg [31:0] _RAND_1859;
  reg [31:0] _RAND_1860;
  reg [31:0] _RAND_1861;
  reg [31:0] _RAND_1862;
  reg [31:0] _RAND_1863;
  reg [31:0] _RAND_1864;
  reg [31:0] _RAND_1865;
  reg [31:0] _RAND_1866;
  reg [31:0] _RAND_1867;
  reg [31:0] _RAND_1868;
  reg [31:0] _RAND_1869;
  reg [31:0] _RAND_1870;
  reg [31:0] _RAND_1871;
  reg [31:0] _RAND_1872;
  reg [31:0] _RAND_1873;
  reg [31:0] _RAND_1874;
  reg [31:0] _RAND_1875;
  reg [31:0] _RAND_1876;
  reg [31:0] _RAND_1877;
  reg [31:0] _RAND_1878;
  reg [31:0] _RAND_1879;
  reg [31:0] _RAND_1880;
  reg [31:0] _RAND_1881;
  reg [31:0] _RAND_1882;
  reg [31:0] _RAND_1883;
  reg [31:0] _RAND_1884;
  reg [31:0] _RAND_1885;
  reg [31:0] _RAND_1886;
  reg [63:0] _RAND_1887;
  reg [31:0] _RAND_1888;
  reg [31:0] _RAND_1889;
  reg [31:0] _RAND_1890;
  reg [31:0] _RAND_1891;
  reg [31:0] _RAND_1892;
  reg [31:0] _RAND_1893;
  reg [31:0] _RAND_1894;
  reg [31:0] _RAND_1895;
  reg [31:0] _RAND_1896;
  reg [31:0] _RAND_1897;
  reg [31:0] _RAND_1898;
  reg [31:0] _RAND_1899;
  reg [31:0] _RAND_1900;
  reg [31:0] _RAND_1901;
  reg [31:0] _RAND_1902;
  reg [31:0] _RAND_1903;
  reg [31:0] _RAND_1904;
  reg [31:0] _RAND_1905;
  reg [31:0] _RAND_1906;
  reg [31:0] _RAND_1907;
  reg [31:0] _RAND_1908;
  reg [31:0] _RAND_1909;
  reg [31:0] _RAND_1910;
  reg [31:0] _RAND_1911;
  reg [31:0] _RAND_1912;
  reg [31:0] _RAND_1913;
  reg [31:0] _RAND_1914;
  reg [31:0] _RAND_1915;
  reg [31:0] _RAND_1916;
  reg [31:0] _RAND_1917;
  reg [31:0] _RAND_1918;
  reg [31:0] _RAND_1919;
  reg [31:0] _RAND_1920;
  reg [31:0] _RAND_1921;
  reg [31:0] _RAND_1922;
  reg [31:0] _RAND_1923;
  reg [31:0] _RAND_1924;
  reg [31:0] _RAND_1925;
  reg [31:0] _RAND_1926;
  reg [31:0] _RAND_1927;
  reg [31:0] _RAND_1928;
  reg [31:0] _RAND_1929;
  reg [63:0] _RAND_1930;
  reg [31:0] _RAND_1931;
  reg [31:0] _RAND_1932;
  reg [31:0] _RAND_1933;
  reg [31:0] _RAND_1934;
  reg [31:0] _RAND_1935;
  reg [31:0] _RAND_1936;
  reg [31:0] _RAND_1937;
  reg [31:0] _RAND_1938;
  reg [31:0] _RAND_1939;
  reg [31:0] _RAND_1940;
  reg [31:0] _RAND_1941;
  reg [31:0] _RAND_1942;
  reg [31:0] _RAND_1943;
  reg [31:0] _RAND_1944;
  reg [31:0] _RAND_1945;
  reg [31:0] _RAND_1946;
  reg [31:0] _RAND_1947;
  reg [31:0] _RAND_1948;
  reg [31:0] _RAND_1949;
  reg [31:0] _RAND_1950;
  reg [31:0] _RAND_1951;
  reg [31:0] _RAND_1952;
  reg [31:0] _RAND_1953;
  reg [31:0] _RAND_1954;
  reg [31:0] _RAND_1955;
  reg [31:0] _RAND_1956;
  reg [31:0] _RAND_1957;
  reg [31:0] _RAND_1958;
  reg [31:0] _RAND_1959;
  reg [31:0] _RAND_1960;
  reg [31:0] _RAND_1961;
  reg [31:0] _RAND_1962;
  reg [31:0] _RAND_1963;
  reg [31:0] _RAND_1964;
  reg [31:0] _RAND_1965;
  reg [63:0] _RAND_1966;
  reg [31:0] _RAND_1967;
  reg [31:0] _RAND_1968;
  reg [31:0] _RAND_1969;
  reg [31:0] _RAND_1970;
  reg [31:0] _RAND_1971;
  reg [31:0] _RAND_1972;
  reg [31:0] _RAND_1973;
  reg [31:0] _RAND_1974;
  reg [31:0] _RAND_1975;
  reg [31:0] _RAND_1976;
  reg [31:0] _RAND_1977;
  reg [31:0] _RAND_1978;
  reg [31:0] _RAND_1979;
  reg [31:0] _RAND_1980;
  reg [31:0] _RAND_1981;
  reg [31:0] _RAND_1982;
  reg [31:0] _RAND_1983;
  reg [31:0] _RAND_1984;
  reg [31:0] _RAND_1985;
  reg [31:0] _RAND_1986;
  reg [31:0] _RAND_1987;
  reg [31:0] _RAND_1988;
  reg [31:0] _RAND_1989;
  reg [31:0] _RAND_1990;
  reg [31:0] _RAND_1991;
  reg [31:0] _RAND_1992;
  reg [31:0] _RAND_1993;
  reg [31:0] _RAND_1994;
  reg [31:0] _RAND_1995;
  reg [31:0] _RAND_1996;
  reg [31:0] _RAND_1997;
  reg [31:0] _RAND_1998;
  reg [31:0] _RAND_1999;
  reg [31:0] _RAND_2000;
  reg [31:0] _RAND_2001;
  reg [31:0] _RAND_2002;
  reg [31:0] _RAND_2003;
  reg [31:0] _RAND_2004;
  reg [31:0] _RAND_2005;
  reg [31:0] _RAND_2006;
  reg [31:0] _RAND_2007;
  reg [31:0] _RAND_2008;
  reg [63:0] _RAND_2009;
  reg [31:0] _RAND_2010;
  reg [31:0] _RAND_2011;
  reg [31:0] _RAND_2012;
  reg [31:0] _RAND_2013;
  reg [31:0] _RAND_2014;
  reg [31:0] _RAND_2015;
  reg [31:0] _RAND_2016;
  reg [31:0] _RAND_2017;
  reg [31:0] _RAND_2018;
  reg [31:0] _RAND_2019;
  reg [31:0] _RAND_2020;
  reg [31:0] _RAND_2021;
  reg [31:0] _RAND_2022;
  reg [31:0] _RAND_2023;
  reg [31:0] _RAND_2024;
  reg [31:0] _RAND_2025;
  reg [31:0] _RAND_2026;
  reg [31:0] _RAND_2027;
  reg [31:0] _RAND_2028;
  reg [31:0] _RAND_2029;
  reg [31:0] _RAND_2030;
  reg [31:0] _RAND_2031;
  reg [31:0] _RAND_2032;
  reg [31:0] _RAND_2033;
  reg [31:0] _RAND_2034;
  reg [31:0] _RAND_2035;
  reg [31:0] _RAND_2036;
  reg [31:0] _RAND_2037;
  reg [31:0] _RAND_2038;
  reg [31:0] _RAND_2039;
  reg [31:0] _RAND_2040;
  reg [31:0] _RAND_2041;
  reg [31:0] _RAND_2042;
  reg [31:0] _RAND_2043;
  reg [31:0] _RAND_2044;
  reg [63:0] _RAND_2045;
  reg [31:0] _RAND_2046;
  reg [31:0] _RAND_2047;
  reg [31:0] _RAND_2048;
  reg [31:0] _RAND_2049;
  reg [31:0] _RAND_2050;
  reg [31:0] _RAND_2051;
  reg [31:0] _RAND_2052;
  reg [31:0] _RAND_2053;
  reg [31:0] _RAND_2054;
  reg [31:0] _RAND_2055;
  reg [31:0] _RAND_2056;
  reg [31:0] _RAND_2057;
  reg [31:0] _RAND_2058;
  reg [31:0] _RAND_2059;
  reg [31:0] _RAND_2060;
  reg [31:0] _RAND_2061;
  reg [31:0] _RAND_2062;
  reg [31:0] _RAND_2063;
  reg [31:0] _RAND_2064;
  reg [31:0] _RAND_2065;
  reg [31:0] _RAND_2066;
  reg [31:0] _RAND_2067;
  reg [31:0] _RAND_2068;
  reg [31:0] _RAND_2069;
  reg [31:0] _RAND_2070;
  reg [31:0] _RAND_2071;
  reg [31:0] _RAND_2072;
  reg [31:0] _RAND_2073;
  reg [31:0] _RAND_2074;
  reg [31:0] _RAND_2075;
  reg [31:0] _RAND_2076;
  reg [31:0] _RAND_2077;
  reg [31:0] _RAND_2078;
  reg [31:0] _RAND_2079;
  reg [31:0] _RAND_2080;
  reg [31:0] _RAND_2081;
  reg [31:0] _RAND_2082;
  reg [31:0] _RAND_2083;
  reg [31:0] _RAND_2084;
  reg [31:0] _RAND_2085;
  reg [31:0] _RAND_2086;
  reg [31:0] _RAND_2087;
  reg [63:0] _RAND_2088;
  reg [31:0] _RAND_2089;
  reg [31:0] _RAND_2090;
  reg [31:0] _RAND_2091;
  reg [31:0] _RAND_2092;
  reg [31:0] _RAND_2093;
  reg [31:0] _RAND_2094;
  reg [31:0] _RAND_2095;
  reg [31:0] _RAND_2096;
  reg [31:0] _RAND_2097;
  reg [31:0] _RAND_2098;
  reg [31:0] _RAND_2099;
  reg [31:0] _RAND_2100;
  reg [31:0] _RAND_2101;
  reg [31:0] _RAND_2102;
  reg [31:0] _RAND_2103;
  reg [31:0] _RAND_2104;
  reg [31:0] _RAND_2105;
  reg [31:0] _RAND_2106;
  reg [31:0] _RAND_2107;
  reg [31:0] _RAND_2108;
  reg [31:0] _RAND_2109;
  reg [31:0] _RAND_2110;
  reg [31:0] _RAND_2111;
  reg [31:0] _RAND_2112;
  reg [31:0] _RAND_2113;
  reg [31:0] _RAND_2114;
  reg [31:0] _RAND_2115;
  reg [31:0] _RAND_2116;
  reg [31:0] _RAND_2117;
  reg [31:0] _RAND_2118;
  reg [31:0] _RAND_2119;
  reg [31:0] _RAND_2120;
  reg [31:0] _RAND_2121;
  reg [31:0] _RAND_2122;
  reg [31:0] _RAND_2123;
  reg [63:0] _RAND_2124;
  reg [31:0] _RAND_2125;
  reg [31:0] _RAND_2126;
  reg [31:0] _RAND_2127;
  reg [31:0] _RAND_2128;
  reg [31:0] _RAND_2129;
  reg [31:0] _RAND_2130;
  reg [31:0] _RAND_2131;
  reg [31:0] _RAND_2132;
  reg [31:0] _RAND_2133;
  reg [31:0] _RAND_2134;
  reg [31:0] _RAND_2135;
  reg [31:0] _RAND_2136;
  reg [31:0] _RAND_2137;
  reg [31:0] _RAND_2138;
  reg [31:0] _RAND_2139;
  reg [31:0] _RAND_2140;
  reg [31:0] _RAND_2141;
  reg [31:0] _RAND_2142;
  reg [31:0] _RAND_2143;
  reg [31:0] _RAND_2144;
  reg [31:0] _RAND_2145;
  reg [31:0] _RAND_2146;
  reg [31:0] _RAND_2147;
  reg [31:0] _RAND_2148;
  reg [31:0] _RAND_2149;
  reg [31:0] _RAND_2150;
  reg [31:0] _RAND_2151;
  reg [31:0] _RAND_2152;
  reg [31:0] _RAND_2153;
  reg [31:0] _RAND_2154;
  reg [31:0] _RAND_2155;
  reg [31:0] _RAND_2156;
  reg [31:0] _RAND_2157;
  reg [31:0] _RAND_2158;
  reg [31:0] _RAND_2159;
  reg [31:0] _RAND_2160;
  reg [31:0] _RAND_2161;
  reg [31:0] _RAND_2162;
  reg [31:0] _RAND_2163;
  reg [31:0] _RAND_2164;
  reg [31:0] _RAND_2165;
  reg [31:0] _RAND_2166;
  reg [63:0] _RAND_2167;
  reg [31:0] _RAND_2168;
  reg [31:0] _RAND_2169;
  reg [31:0] _RAND_2170;
  reg [31:0] _RAND_2171;
  reg [31:0] _RAND_2172;
  reg [31:0] _RAND_2173;
  reg [31:0] _RAND_2174;
  reg [31:0] _RAND_2175;
  reg [31:0] _RAND_2176;
  reg [31:0] _RAND_2177;
  reg [31:0] _RAND_2178;
  reg [31:0] _RAND_2179;
  reg [31:0] _RAND_2180;
  reg [31:0] _RAND_2181;
  reg [31:0] _RAND_2182;
  reg [31:0] _RAND_2183;
  reg [31:0] _RAND_2184;
  reg [31:0] _RAND_2185;
  reg [31:0] _RAND_2186;
  reg [31:0] _RAND_2187;
  reg [31:0] _RAND_2188;
  reg [31:0] _RAND_2189;
  reg [31:0] _RAND_2190;
  reg [31:0] _RAND_2191;
  reg [31:0] _RAND_2192;
  reg [31:0] _RAND_2193;
  reg [31:0] _RAND_2194;
  reg [31:0] _RAND_2195;
  reg [31:0] _RAND_2196;
  reg [31:0] _RAND_2197;
  reg [31:0] _RAND_2198;
  reg [31:0] _RAND_2199;
  reg [31:0] _RAND_2200;
  reg [31:0] _RAND_2201;
  reg [31:0] _RAND_2202;
  reg [63:0] _RAND_2203;
  reg [31:0] _RAND_2204;
  reg [31:0] _RAND_2205;
  reg [31:0] _RAND_2206;
  reg [31:0] _RAND_2207;
  reg [31:0] _RAND_2208;
  reg [31:0] _RAND_2209;
  reg [31:0] _RAND_2210;
  reg [31:0] _RAND_2211;
  reg [31:0] _RAND_2212;
  reg [31:0] _RAND_2213;
  reg [31:0] _RAND_2214;
  reg [31:0] _RAND_2215;
  reg [31:0] _RAND_2216;
  reg [31:0] _RAND_2217;
  reg [31:0] _RAND_2218;
  reg [31:0] _RAND_2219;
  reg [31:0] _RAND_2220;
  reg [31:0] _RAND_2221;
  reg [31:0] _RAND_2222;
  reg [31:0] _RAND_2223;
  reg [31:0] _RAND_2224;
  reg [31:0] _RAND_2225;
  reg [31:0] _RAND_2226;
  reg [31:0] _RAND_2227;
  reg [31:0] _RAND_2228;
  reg [31:0] _RAND_2229;
  reg [31:0] _RAND_2230;
  reg [31:0] _RAND_2231;
  reg [31:0] _RAND_2232;
  reg [31:0] _RAND_2233;
  reg [31:0] _RAND_2234;
  reg [31:0] _RAND_2235;
  reg [31:0] _RAND_2236;
  reg [31:0] _RAND_2237;
  reg [31:0] _RAND_2238;
  reg [31:0] _RAND_2239;
  reg [31:0] _RAND_2240;
  reg [31:0] _RAND_2241;
  reg [31:0] _RAND_2242;
  reg [31:0] _RAND_2243;
  reg [31:0] _RAND_2244;
  reg [31:0] _RAND_2245;
  reg [63:0] _RAND_2246;
  reg [31:0] _RAND_2247;
  reg [31:0] _RAND_2248;
  reg [31:0] _RAND_2249;
  reg [31:0] _RAND_2250;
  reg [31:0] _RAND_2251;
  reg [31:0] _RAND_2252;
  reg [31:0] _RAND_2253;
  reg [31:0] _RAND_2254;
  reg [31:0] _RAND_2255;
  reg [31:0] _RAND_2256;
  reg [31:0] _RAND_2257;
  reg [31:0] _RAND_2258;
  reg [31:0] _RAND_2259;
  reg [31:0] _RAND_2260;
  reg [31:0] _RAND_2261;
  reg [31:0] _RAND_2262;
  reg [31:0] _RAND_2263;
  reg [31:0] _RAND_2264;
  reg [31:0] _RAND_2265;
  reg [31:0] _RAND_2266;
  reg [31:0] _RAND_2267;
  reg [31:0] _RAND_2268;
  reg [31:0] _RAND_2269;
  reg [31:0] _RAND_2270;
  reg [31:0] _RAND_2271;
  reg [31:0] _RAND_2272;
  reg [31:0] _RAND_2273;
  reg [31:0] _RAND_2274;
  reg [31:0] _RAND_2275;
  reg [31:0] _RAND_2276;
  reg [31:0] _RAND_2277;
  reg [31:0] _RAND_2278;
  reg [31:0] _RAND_2279;
  reg [31:0] _RAND_2280;
  reg [31:0] _RAND_2281;
  reg [63:0] _RAND_2282;
  reg [31:0] _RAND_2283;
  reg [31:0] _RAND_2284;
  reg [31:0] _RAND_2285;
  reg [31:0] _RAND_2286;
  reg [31:0] _RAND_2287;
  reg [31:0] _RAND_2288;
  reg [31:0] _RAND_2289;
  reg [31:0] _RAND_2290;
  reg [31:0] _RAND_2291;
  reg [31:0] _RAND_2292;
  reg [31:0] _RAND_2293;
  reg [31:0] _RAND_2294;
  reg [31:0] _RAND_2295;
  reg [31:0] _RAND_2296;
  reg [31:0] _RAND_2297;
  reg [31:0] _RAND_2298;
  reg [31:0] _RAND_2299;
  reg [31:0] _RAND_2300;
  reg [31:0] _RAND_2301;
  reg [31:0] _RAND_2302;
  reg [31:0] _RAND_2303;
  reg [31:0] _RAND_2304;
  reg [31:0] _RAND_2305;
  reg [31:0] _RAND_2306;
  reg [31:0] _RAND_2307;
  reg [31:0] _RAND_2308;
  reg [31:0] _RAND_2309;
  reg [31:0] _RAND_2310;
  reg [31:0] _RAND_2311;
  reg [31:0] _RAND_2312;
  reg [31:0] _RAND_2313;
  reg [31:0] _RAND_2314;
  reg [31:0] _RAND_2315;
  reg [31:0] _RAND_2316;
  reg [31:0] _RAND_2317;
  reg [31:0] _RAND_2318;
  reg [31:0] _RAND_2319;
  reg [31:0] _RAND_2320;
  reg [31:0] _RAND_2321;
  reg [31:0] _RAND_2322;
  reg [31:0] _RAND_2323;
  reg [31:0] _RAND_2324;
  reg [63:0] _RAND_2325;
  reg [31:0] _RAND_2326;
  reg [31:0] _RAND_2327;
  reg [31:0] _RAND_2328;
  reg [31:0] _RAND_2329;
  reg [31:0] _RAND_2330;
  reg [31:0] _RAND_2331;
  reg [31:0] _RAND_2332;
  reg [31:0] _RAND_2333;
  reg [31:0] _RAND_2334;
  reg [31:0] _RAND_2335;
  reg [31:0] _RAND_2336;
  reg [31:0] _RAND_2337;
  reg [31:0] _RAND_2338;
  reg [31:0] _RAND_2339;
  reg [31:0] _RAND_2340;
  reg [31:0] _RAND_2341;
  reg [31:0] _RAND_2342;
  reg [31:0] _RAND_2343;
  reg [31:0] _RAND_2344;
  reg [31:0] _RAND_2345;
  reg [31:0] _RAND_2346;
  reg [31:0] _RAND_2347;
  reg [31:0] _RAND_2348;
  reg [31:0] _RAND_2349;
  reg [31:0] _RAND_2350;
  reg [31:0] _RAND_2351;
  reg [31:0] _RAND_2352;
  reg [31:0] _RAND_2353;
  reg [31:0] _RAND_2354;
  reg [31:0] _RAND_2355;
  reg [31:0] _RAND_2356;
  reg [31:0] _RAND_2357;
  reg [31:0] _RAND_2358;
  reg [31:0] _RAND_2359;
  reg [31:0] _RAND_2360;
  reg [63:0] _RAND_2361;
  reg [31:0] _RAND_2362;
  reg [31:0] _RAND_2363;
  reg [31:0] _RAND_2364;
  reg [31:0] _RAND_2365;
  reg [31:0] _RAND_2366;
  reg [31:0] _RAND_2367;
  reg [31:0] _RAND_2368;
  reg [31:0] _RAND_2369;
  reg [31:0] _RAND_2370;
  reg [31:0] _RAND_2371;
  reg [31:0] _RAND_2372;
  reg [31:0] _RAND_2373;
  reg [31:0] _RAND_2374;
  reg [31:0] _RAND_2375;
  reg [31:0] _RAND_2376;
  reg [31:0] _RAND_2377;
  reg [31:0] _RAND_2378;
  reg [31:0] _RAND_2379;
  reg [31:0] _RAND_2380;
  reg [31:0] _RAND_2381;
  reg [31:0] _RAND_2382;
  reg [31:0] _RAND_2383;
  reg [31:0] _RAND_2384;
  reg [31:0] _RAND_2385;
  reg [31:0] _RAND_2386;
  reg [31:0] _RAND_2387;
  reg [31:0] _RAND_2388;
  reg [31:0] _RAND_2389;
  reg [31:0] _RAND_2390;
  reg [31:0] _RAND_2391;
  reg [31:0] _RAND_2392;
  reg [31:0] _RAND_2393;
  reg [31:0] _RAND_2394;
  reg [31:0] _RAND_2395;
  reg [31:0] _RAND_2396;
  reg [31:0] _RAND_2397;
  reg [31:0] _RAND_2398;
  reg [31:0] _RAND_2399;
  reg [31:0] _RAND_2400;
  reg [31:0] _RAND_2401;
  reg [31:0] _RAND_2402;
  reg [31:0] _RAND_2403;
  reg [63:0] _RAND_2404;
  reg [31:0] _RAND_2405;
  reg [31:0] _RAND_2406;
  reg [31:0] _RAND_2407;
  reg [31:0] _RAND_2408;
  reg [31:0] _RAND_2409;
  reg [31:0] _RAND_2410;
  reg [31:0] _RAND_2411;
  reg [31:0] _RAND_2412;
  reg [31:0] _RAND_2413;
  reg [31:0] _RAND_2414;
  reg [31:0] _RAND_2415;
  reg [31:0] _RAND_2416;
  reg [31:0] _RAND_2417;
  reg [31:0] _RAND_2418;
  reg [31:0] _RAND_2419;
  reg [31:0] _RAND_2420;
  reg [31:0] _RAND_2421;
  reg [31:0] _RAND_2422;
  reg [31:0] _RAND_2423;
  reg [31:0] _RAND_2424;
  reg [31:0] _RAND_2425;
  reg [31:0] _RAND_2426;
  reg [31:0] _RAND_2427;
  reg [31:0] _RAND_2428;
  reg [31:0] _RAND_2429;
  reg [31:0] _RAND_2430;
  reg [31:0] _RAND_2431;
  reg [31:0] _RAND_2432;
  reg [31:0] _RAND_2433;
  reg [31:0] _RAND_2434;
  reg [31:0] _RAND_2435;
  reg [31:0] _RAND_2436;
  reg [31:0] _RAND_2437;
  reg [31:0] _RAND_2438;
  reg [31:0] _RAND_2439;
  reg [63:0] _RAND_2440;
  reg [31:0] _RAND_2441;
  reg [31:0] _RAND_2442;
  reg [31:0] _RAND_2443;
  reg [31:0] _RAND_2444;
  reg [31:0] _RAND_2445;
  reg [31:0] _RAND_2446;
  reg [31:0] _RAND_2447;
  reg [31:0] _RAND_2448;
  reg [31:0] _RAND_2449;
  reg [31:0] _RAND_2450;
  reg [31:0] _RAND_2451;
  reg [31:0] _RAND_2452;
  reg [31:0] _RAND_2453;
  reg [31:0] _RAND_2454;
  reg [31:0] _RAND_2455;
  reg [31:0] _RAND_2456;
  reg [31:0] _RAND_2457;
  reg [31:0] _RAND_2458;
  reg [31:0] _RAND_2459;
  reg [31:0] _RAND_2460;
  reg [31:0] _RAND_2461;
  reg [31:0] _RAND_2462;
  reg [31:0] _RAND_2463;
  reg [31:0] _RAND_2464;
  reg [31:0] _RAND_2465;
  reg [31:0] _RAND_2466;
  reg [31:0] _RAND_2467;
  reg [31:0] _RAND_2468;
  reg [31:0] _RAND_2469;
  reg [31:0] _RAND_2470;
  reg [31:0] _RAND_2471;
  reg [31:0] _RAND_2472;
  reg [31:0] _RAND_2473;
  reg [31:0] _RAND_2474;
  reg [31:0] _RAND_2475;
  reg [31:0] _RAND_2476;
  reg [31:0] _RAND_2477;
  reg [31:0] _RAND_2478;
  reg [31:0] _RAND_2479;
  reg [31:0] _RAND_2480;
  reg [31:0] _RAND_2481;
  reg [31:0] _RAND_2482;
  reg [63:0] _RAND_2483;
  reg [31:0] _RAND_2484;
  reg [31:0] _RAND_2485;
  reg [31:0] _RAND_2486;
  reg [31:0] _RAND_2487;
  reg [31:0] _RAND_2488;
  reg [31:0] _RAND_2489;
  reg [31:0] _RAND_2490;
  reg [31:0] _RAND_2491;
  reg [31:0] _RAND_2492;
  reg [31:0] _RAND_2493;
  reg [31:0] _RAND_2494;
  reg [31:0] _RAND_2495;
  reg [31:0] _RAND_2496;
  reg [31:0] _RAND_2497;
  reg [31:0] _RAND_2498;
  reg [31:0] _RAND_2499;
  reg [31:0] _RAND_2500;
  reg [31:0] _RAND_2501;
  reg [31:0] _RAND_2502;
  reg [31:0] _RAND_2503;
  reg [31:0] _RAND_2504;
  reg [31:0] _RAND_2505;
  reg [31:0] _RAND_2506;
  reg [31:0] _RAND_2507;
  reg [31:0] _RAND_2508;
  reg [31:0] _RAND_2509;
  reg [31:0] _RAND_2510;
  reg [31:0] _RAND_2511;
  reg [31:0] _RAND_2512;
  reg [31:0] _RAND_2513;
  reg [31:0] _RAND_2514;
  reg [31:0] _RAND_2515;
  reg [31:0] _RAND_2516;
  reg [31:0] _RAND_2517;
  reg [31:0] _RAND_2518;
  reg [63:0] _RAND_2519;
  reg [31:0] _RAND_2520;
  reg [31:0] _RAND_2521;
  reg [31:0] _RAND_2522;
  reg [31:0] _RAND_2523;
  reg [31:0] _RAND_2524;
  reg [31:0] _RAND_2525;
  reg [31:0] _RAND_2526;
  reg [31:0] _RAND_2527;
  reg [31:0] _RAND_2528;
  reg [31:0] _RAND_2529;
  reg [31:0] _RAND_2530;
  reg [31:0] _RAND_2531;
  reg [31:0] _RAND_2532;
  reg [31:0] _RAND_2533;
  reg [31:0] _RAND_2534;
  reg [31:0] _RAND_2535;
  reg [31:0] _RAND_2536;
  reg [31:0] _RAND_2537;
  reg [31:0] _RAND_2538;
  reg [31:0] _RAND_2539;
  reg [31:0] _RAND_2540;
  reg [31:0] _RAND_2541;
  reg [31:0] _RAND_2542;
  reg [31:0] _RAND_2543;
  reg [31:0] _RAND_2544;
  reg [31:0] _RAND_2545;
  reg [31:0] _RAND_2546;
  reg [31:0] _RAND_2547;
  reg [31:0] _RAND_2548;
  reg [31:0] _RAND_2549;
  reg [31:0] _RAND_2550;
  reg [31:0] _RAND_2551;
  reg [31:0] _RAND_2552;
  reg [31:0] _RAND_2553;
  reg [31:0] _RAND_2554;
  reg [31:0] _RAND_2555;
  reg [31:0] _RAND_2556;
  reg [31:0] _RAND_2557;
  reg [31:0] _RAND_2558;
  reg [31:0] _RAND_2559;
  reg [31:0] _RAND_2560;
  reg [31:0] _RAND_2561;
  reg [63:0] _RAND_2562;
  reg [31:0] _RAND_2563;
  reg [31:0] _RAND_2564;
  reg [31:0] _RAND_2565;
  reg [31:0] _RAND_2566;
  reg [31:0] _RAND_2567;
  reg [31:0] _RAND_2568;
  reg [31:0] _RAND_2569;
  reg [31:0] _RAND_2570;
  reg [31:0] _RAND_2571;
  reg [31:0] _RAND_2572;
  reg [31:0] _RAND_2573;
  reg [31:0] _RAND_2574;
  reg [31:0] _RAND_2575;
  reg [31:0] _RAND_2576;
  reg [31:0] _RAND_2577;
  reg [31:0] _RAND_2578;
  reg [31:0] _RAND_2579;
  reg [31:0] _RAND_2580;
  reg [31:0] _RAND_2581;
  reg [31:0] _RAND_2582;
  reg [31:0] _RAND_2583;
  reg [31:0] _RAND_2584;
  reg [31:0] _RAND_2585;
  reg [31:0] _RAND_2586;
  reg [31:0] _RAND_2587;
  reg [31:0] _RAND_2588;
  reg [31:0] _RAND_2589;
  reg [31:0] _RAND_2590;
  reg [31:0] _RAND_2591;
  reg [31:0] _RAND_2592;
  reg [31:0] _RAND_2593;
  reg [31:0] _RAND_2594;
  reg [31:0] _RAND_2595;
  reg [31:0] _RAND_2596;
  reg [31:0] _RAND_2597;
  reg [63:0] _RAND_2598;
  reg [31:0] _RAND_2599;
  reg [31:0] _RAND_2600;
  reg [31:0] _RAND_2601;
  reg [31:0] _RAND_2602;
  reg [31:0] _RAND_2603;
  reg [31:0] _RAND_2604;
  reg [31:0] _RAND_2605;
  reg [31:0] _RAND_2606;
  reg [31:0] _RAND_2607;
  reg [31:0] _RAND_2608;
  reg [31:0] _RAND_2609;
  reg [31:0] _RAND_2610;
  reg [31:0] _RAND_2611;
  reg [31:0] _RAND_2612;
  reg [31:0] _RAND_2613;
  reg [31:0] _RAND_2614;
  reg [31:0] _RAND_2615;
  reg [31:0] _RAND_2616;
  reg [31:0] _RAND_2617;
  reg [31:0] _RAND_2618;
  reg [31:0] _RAND_2619;
  reg [31:0] _RAND_2620;
  reg [31:0] _RAND_2621;
  reg [31:0] _RAND_2622;
  reg [31:0] _RAND_2623;
  reg [31:0] _RAND_2624;
  reg [31:0] _RAND_2625;
  reg [31:0] _RAND_2626;
  reg [31:0] _RAND_2627;
  reg [31:0] _RAND_2628;
  reg [31:0] _RAND_2629;
  reg [31:0] _RAND_2630;
  reg [31:0] _RAND_2631;
  reg [31:0] _RAND_2632;
  reg [31:0] _RAND_2633;
  reg [31:0] _RAND_2634;
  reg [31:0] _RAND_2635;
  reg [31:0] _RAND_2636;
  reg [31:0] _RAND_2637;
  reg [31:0] _RAND_2638;
  reg [31:0] _RAND_2639;
  reg [31:0] _RAND_2640;
  reg [63:0] _RAND_2641;
  reg [31:0] _RAND_2642;
  reg [31:0] _RAND_2643;
  reg [31:0] _RAND_2644;
  reg [31:0] _RAND_2645;
  reg [31:0] _RAND_2646;
  reg [31:0] _RAND_2647;
  reg [31:0] _RAND_2648;
  reg [31:0] _RAND_2649;
  reg [31:0] _RAND_2650;
  reg [31:0] _RAND_2651;
  reg [31:0] _RAND_2652;
  reg [31:0] _RAND_2653;
  reg [31:0] _RAND_2654;
  reg [31:0] _RAND_2655;
  reg [31:0] _RAND_2656;
  reg [31:0] _RAND_2657;
  reg [31:0] _RAND_2658;
  reg [31:0] _RAND_2659;
  reg [31:0] _RAND_2660;
  reg [31:0] _RAND_2661;
  reg [31:0] _RAND_2662;
  reg [31:0] _RAND_2663;
  reg [31:0] _RAND_2664;
  reg [31:0] _RAND_2665;
  reg [31:0] _RAND_2666;
  reg [31:0] _RAND_2667;
  reg [31:0] _RAND_2668;
  reg [31:0] _RAND_2669;
  reg [31:0] _RAND_2670;
  reg [31:0] _RAND_2671;
  reg [31:0] _RAND_2672;
  reg [31:0] _RAND_2673;
  reg [31:0] _RAND_2674;
  reg [31:0] _RAND_2675;
  reg [31:0] _RAND_2676;
  reg [31:0] _RAND_2677;
  reg [31:0] _RAND_2678;
  reg [31:0] _RAND_2679;
  reg [31:0] _RAND_2680;
  reg [31:0] _RAND_2681;
  reg [31:0] _RAND_2682;
  reg [31:0] _RAND_2683;
  reg [31:0] _RAND_2684;
  reg [31:0] _RAND_2685;
  reg [31:0] _RAND_2686;
  reg [31:0] _RAND_2687;
  reg [31:0] _RAND_2688;
  reg [31:0] _RAND_2689;
  reg [31:0] _RAND_2690;
  reg [31:0] _RAND_2691;
  reg [31:0] _RAND_2692;
  reg [31:0] _RAND_2693;
  reg [31:0] _RAND_2694;
  reg [31:0] _RAND_2695;
  reg [31:0] _RAND_2696;
  reg [31:0] _RAND_2697;
  reg [31:0] _RAND_2698;
  reg [31:0] _RAND_2699;
  reg [31:0] _RAND_2700;
  reg [31:0] _RAND_2701;
  reg [31:0] _RAND_2702;
  reg [31:0] _RAND_2703;
  reg [31:0] _RAND_2704;
  reg [31:0] _RAND_2705;
  reg [31:0] _RAND_2706;
  reg [31:0] _RAND_2707;
  reg [31:0] _RAND_2708;
  reg [31:0] _RAND_2709;
  reg [31:0] _RAND_2710;
  reg [31:0] _RAND_2711;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] rob_debug_inst_mem_0 [0:31]; // @[rob.scala 297:41]
  wire  rob_debug_inst_mem_0_rob_debug_inst_rdata_en; // @[rob.scala 297:41]
  wire [4:0] rob_debug_inst_mem_0_rob_debug_inst_rdata_addr; // @[rob.scala 297:41]
  wire [31:0] rob_debug_inst_mem_0_rob_debug_inst_rdata_data; // @[rob.scala 297:41]
  wire [31:0] rob_debug_inst_mem_0__T_3_data; // @[rob.scala 297:41]
  wire [4:0] rob_debug_inst_mem_0__T_3_addr; // @[rob.scala 297:41]
  wire  rob_debug_inst_mem_0__T_3_mask; // @[rob.scala 297:41]
  wire  rob_debug_inst_mem_0__T_3_en; // @[rob.scala 297:41]
  reg  rob_debug_inst_mem_0_rob_debug_inst_rdata_en_pipe_0;
  reg [4:0] rob_debug_inst_mem_0_rob_debug_inst_rdata_addr_pipe_0;
  reg [4:0] rob_fflags [0:31]; // @[rob.scala 313:28]
  wire  rob_fflags__T_221_en; // @[rob.scala 313:28]
  wire [4:0] rob_fflags__T_221_addr; // @[rob.scala 313:28]
  wire [4:0] rob_fflags__T_221_data; // @[rob.scala 313:28]
  wire [4:0] rob_fflags__T_15_data; // @[rob.scala 313:28]
  wire [4:0] rob_fflags__T_15_addr; // @[rob.scala 313:28]
  wire  rob_fflags__T_15_mask; // @[rob.scala 313:28]
  wire  rob_fflags__T_15_en; // @[rob.scala 313:28]
  wire [4:0] rob_fflags__T_59_data; // @[rob.scala 313:28]
  wire [4:0] rob_fflags__T_59_addr; // @[rob.scala 313:28]
  wire  rob_fflags__T_59_mask; // @[rob.scala 313:28]
  wire  rob_fflags__T_59_en; // @[rob.scala 313:28]
  wire [4:0] rob_fflags__T_62_data; // @[rob.scala 313:28]
  wire [4:0] rob_fflags__T_62_addr; // @[rob.scala 313:28]
  wire  rob_fflags__T_62_mask; // @[rob.scala 313:28]
  wire  rob_fflags__T_62_en; // @[rob.scala 313:28]
  reg [63:0] rob_debug_wdata [0:31]; // @[rob.scala 315:30]
  wire  rob_debug_wdata__T_400_en; // @[rob.scala 315:30]
  wire [4:0] rob_debug_wdata__T_400_addr; // @[rob.scala 315:30]
  wire [63:0] rob_debug_wdata__T_400_data; // @[rob.scala 315:30]
  wire [63:0] rob_debug_wdata__T_290_data; // @[rob.scala 315:30]
  wire [4:0] rob_debug_wdata__T_290_addr; // @[rob.scala 315:30]
  wire  rob_debug_wdata__T_290_mask; // @[rob.scala 315:30]
  wire  rob_debug_wdata__T_290_en; // @[rob.scala 315:30]
  wire [63:0] rob_debug_wdata__T_318_data; // @[rob.scala 315:30]
  wire [4:0] rob_debug_wdata__T_318_addr; // @[rob.scala 315:30]
  wire  rob_debug_wdata__T_318_mask; // @[rob.scala 315:30]
  wire  rob_debug_wdata__T_318_en; // @[rob.scala 315:30]
  wire [63:0] rob_debug_wdata__T_346_data; // @[rob.scala 315:30]
  wire [4:0] rob_debug_wdata__T_346_addr; // @[rob.scala 315:30]
  wire  rob_debug_wdata__T_346_mask; // @[rob.scala 315:30]
  wire  rob_debug_wdata__T_346_en; // @[rob.scala 315:30]
  wire [63:0] rob_debug_wdata__T_374_data; // @[rob.scala 315:30]
  wire [4:0] rob_debug_wdata__T_374_addr; // @[rob.scala 315:30]
  wire  rob_debug_wdata__T_374_mask; // @[rob.scala 315:30]
  wire  rob_debug_wdata__T_374_en; // @[rob.scala 315:30]
  reg [1:0] rob_state; // @[rob.scala 221:26]
  reg [4:0] rob_head; // @[rob.scala 224:29]
  reg [4:0] rob_tail; // @[rob.scala 228:29]
  reg [4:0] rob_pnr; // @[rob.scala 232:29]
  wire  _T = rob_state == 2'h2; // @[rob.scala 236:31]
  wire [4:0] com_idx = rob_state == 2'h2 ? rob_tail : rob_head; // @[rob.scala 236:20]
  reg  maybe_full; // @[rob.scala 239:29]
  reg  r_xcpt_val; // @[rob.scala 258:33]
  reg [7:0] r_xcpt_uop_br_mask; // @[rob.scala 259:29]
  reg [4:0] r_xcpt_uop_rob_idx; // @[rob.scala 259:29]
  reg [63:0] r_xcpt_uop_exc_cause; // @[rob.scala 259:29]
  reg [39:0] r_xcpt_badvaddr; // @[rob.scala 260:29]
  reg  rob_val_31; // @[rob.scala 307:32]
  reg  rob_val_30; // @[rob.scala 307:32]
  reg  rob_val_29; // @[rob.scala 307:32]
  reg  rob_val_28; // @[rob.scala 307:32]
  reg  rob_val_27; // @[rob.scala 307:32]
  reg  rob_val_26; // @[rob.scala 307:32]
  reg  rob_val_25; // @[rob.scala 307:32]
  reg  rob_val_24; // @[rob.scala 307:32]
  reg  rob_val_23; // @[rob.scala 307:32]
  reg  rob_val_22; // @[rob.scala 307:32]
  reg  rob_val_21; // @[rob.scala 307:32]
  reg  rob_val_20; // @[rob.scala 307:32]
  reg  rob_val_19; // @[rob.scala 307:32]
  reg  rob_val_18; // @[rob.scala 307:32]
  reg  rob_val_17; // @[rob.scala 307:32]
  reg  rob_val_16; // @[rob.scala 307:32]
  reg  rob_val_15; // @[rob.scala 307:32]
  reg  rob_val_14; // @[rob.scala 307:32]
  reg  rob_val_13; // @[rob.scala 307:32]
  reg  rob_val_12; // @[rob.scala 307:32]
  reg  rob_val_11; // @[rob.scala 307:32]
  reg  rob_val_10; // @[rob.scala 307:32]
  reg  rob_val_9; // @[rob.scala 307:32]
  reg  rob_val_8; // @[rob.scala 307:32]
  reg  rob_val_7; // @[rob.scala 307:32]
  reg  rob_val_6; // @[rob.scala 307:32]
  reg  rob_val_5; // @[rob.scala 307:32]
  reg  rob_val_4; // @[rob.scala 307:32]
  reg  rob_val_3; // @[rob.scala 307:32]
  reg  rob_val_2; // @[rob.scala 307:32]
  reg  rob_val_1; // @[rob.scala 307:32]
  reg  rob_val_0; // @[rob.scala 307:32]
  wire  _GEN_6806 = 5'h1 == rob_head ? rob_val_1 : rob_val_0; // @[rob.scala 398:{49,49}]
  wire  _GEN_6807 = 5'h2 == rob_head ? rob_val_2 : _GEN_6806; // @[rob.scala 398:{49,49}]
  wire  _GEN_6808 = 5'h3 == rob_head ? rob_val_3 : _GEN_6807; // @[rob.scala 398:{49,49}]
  wire  _GEN_6809 = 5'h4 == rob_head ? rob_val_4 : _GEN_6808; // @[rob.scala 398:{49,49}]
  wire  _GEN_6810 = 5'h5 == rob_head ? rob_val_5 : _GEN_6809; // @[rob.scala 398:{49,49}]
  wire  _GEN_6811 = 5'h6 == rob_head ? rob_val_6 : _GEN_6810; // @[rob.scala 398:{49,49}]
  wire  _GEN_6812 = 5'h7 == rob_head ? rob_val_7 : _GEN_6811; // @[rob.scala 398:{49,49}]
  wire  _GEN_6813 = 5'h8 == rob_head ? rob_val_8 : _GEN_6812; // @[rob.scala 398:{49,49}]
  wire  _GEN_6814 = 5'h9 == rob_head ? rob_val_9 : _GEN_6813; // @[rob.scala 398:{49,49}]
  wire  _GEN_6815 = 5'ha == rob_head ? rob_val_10 : _GEN_6814; // @[rob.scala 398:{49,49}]
  wire  _GEN_6816 = 5'hb == rob_head ? rob_val_11 : _GEN_6815; // @[rob.scala 398:{49,49}]
  wire  _GEN_6817 = 5'hc == rob_head ? rob_val_12 : _GEN_6816; // @[rob.scala 398:{49,49}]
  wire  _GEN_6818 = 5'hd == rob_head ? rob_val_13 : _GEN_6817; // @[rob.scala 398:{49,49}]
  wire  _GEN_6819 = 5'he == rob_head ? rob_val_14 : _GEN_6818; // @[rob.scala 398:{49,49}]
  wire  _GEN_6820 = 5'hf == rob_head ? rob_val_15 : _GEN_6819; // @[rob.scala 398:{49,49}]
  wire  _GEN_6821 = 5'h10 == rob_head ? rob_val_16 : _GEN_6820; // @[rob.scala 398:{49,49}]
  wire  _GEN_6822 = 5'h11 == rob_head ? rob_val_17 : _GEN_6821; // @[rob.scala 398:{49,49}]
  wire  _GEN_6823 = 5'h12 == rob_head ? rob_val_18 : _GEN_6822; // @[rob.scala 398:{49,49}]
  wire  _GEN_6824 = 5'h13 == rob_head ? rob_val_19 : _GEN_6823; // @[rob.scala 398:{49,49}]
  wire  _GEN_6825 = 5'h14 == rob_head ? rob_val_20 : _GEN_6824; // @[rob.scala 398:{49,49}]
  wire  _GEN_6826 = 5'h15 == rob_head ? rob_val_21 : _GEN_6825; // @[rob.scala 398:{49,49}]
  wire  _GEN_6827 = 5'h16 == rob_head ? rob_val_22 : _GEN_6826; // @[rob.scala 398:{49,49}]
  wire  _GEN_6828 = 5'h17 == rob_head ? rob_val_23 : _GEN_6827; // @[rob.scala 398:{49,49}]
  wire  _GEN_6829 = 5'h18 == rob_head ? rob_val_24 : _GEN_6828; // @[rob.scala 398:{49,49}]
  wire  _GEN_6830 = 5'h19 == rob_head ? rob_val_25 : _GEN_6829; // @[rob.scala 398:{49,49}]
  wire  _GEN_6831 = 5'h1a == rob_head ? rob_val_26 : _GEN_6830; // @[rob.scala 398:{49,49}]
  wire  _GEN_6832 = 5'h1b == rob_head ? rob_val_27 : _GEN_6831; // @[rob.scala 398:{49,49}]
  wire  _GEN_6833 = 5'h1c == rob_head ? rob_val_28 : _GEN_6832; // @[rob.scala 398:{49,49}]
  wire  _GEN_6834 = 5'h1d == rob_head ? rob_val_29 : _GEN_6833; // @[rob.scala 398:{49,49}]
  wire  _GEN_6835 = 5'h1e == rob_head ? rob_val_30 : _GEN_6834; // @[rob.scala 398:{49,49}]
  wire  rob_head_vals_0 = 5'h1f == rob_head ? rob_val_31 : _GEN_6835; // @[rob.scala 398:{49,49}]
  reg  rob_bsy_31; // @[rob.scala 308:28]
  reg  rob_bsy_30; // @[rob.scala 308:28]
  reg  rob_bsy_29; // @[rob.scala 308:28]
  reg  rob_bsy_28; // @[rob.scala 308:28]
  reg  rob_bsy_27; // @[rob.scala 308:28]
  reg  rob_bsy_26; // @[rob.scala 308:28]
  reg  rob_bsy_25; // @[rob.scala 308:28]
  reg  rob_bsy_24; // @[rob.scala 308:28]
  reg  rob_bsy_23; // @[rob.scala 308:28]
  reg  rob_bsy_22; // @[rob.scala 308:28]
  reg  rob_bsy_21; // @[rob.scala 308:28]
  reg  rob_bsy_20; // @[rob.scala 308:28]
  reg  rob_bsy_19; // @[rob.scala 308:28]
  reg  rob_bsy_18; // @[rob.scala 308:28]
  reg  rob_bsy_17; // @[rob.scala 308:28]
  reg  rob_bsy_16; // @[rob.scala 308:28]
  reg  rob_bsy_15; // @[rob.scala 308:28]
  reg  rob_bsy_14; // @[rob.scala 308:28]
  reg  rob_bsy_13; // @[rob.scala 308:28]
  reg  rob_bsy_12; // @[rob.scala 308:28]
  reg  rob_bsy_11; // @[rob.scala 308:28]
  reg  rob_bsy_10; // @[rob.scala 308:28]
  reg  rob_bsy_9; // @[rob.scala 308:28]
  reg  rob_bsy_8; // @[rob.scala 308:28]
  reg  rob_bsy_7; // @[rob.scala 308:28]
  reg  rob_bsy_6; // @[rob.scala 308:28]
  reg  rob_bsy_5; // @[rob.scala 308:28]
  reg  rob_bsy_4; // @[rob.scala 308:28]
  reg  rob_bsy_3; // @[rob.scala 308:28]
  reg  rob_bsy_2; // @[rob.scala 308:28]
  reg  rob_bsy_1; // @[rob.scala 308:28]
  reg  rob_bsy_0; // @[rob.scala 308:28]
  wire  _GEN_6870 = 5'h1 == rob_head ? rob_bsy_1 : rob_bsy_0; // @[rob.scala 404:{43,43}]
  wire  _GEN_6871 = 5'h2 == rob_head ? rob_bsy_2 : _GEN_6870; // @[rob.scala 404:{43,43}]
  wire  _GEN_6872 = 5'h3 == rob_head ? rob_bsy_3 : _GEN_6871; // @[rob.scala 404:{43,43}]
  wire  _GEN_6873 = 5'h4 == rob_head ? rob_bsy_4 : _GEN_6872; // @[rob.scala 404:{43,43}]
  wire  _GEN_6874 = 5'h5 == rob_head ? rob_bsy_5 : _GEN_6873; // @[rob.scala 404:{43,43}]
  wire  _GEN_6875 = 5'h6 == rob_head ? rob_bsy_6 : _GEN_6874; // @[rob.scala 404:{43,43}]
  wire  _GEN_6876 = 5'h7 == rob_head ? rob_bsy_7 : _GEN_6875; // @[rob.scala 404:{43,43}]
  wire  _GEN_6877 = 5'h8 == rob_head ? rob_bsy_8 : _GEN_6876; // @[rob.scala 404:{43,43}]
  wire  _GEN_6878 = 5'h9 == rob_head ? rob_bsy_9 : _GEN_6877; // @[rob.scala 404:{43,43}]
  wire  _GEN_6879 = 5'ha == rob_head ? rob_bsy_10 : _GEN_6878; // @[rob.scala 404:{43,43}]
  wire  _GEN_6880 = 5'hb == rob_head ? rob_bsy_11 : _GEN_6879; // @[rob.scala 404:{43,43}]
  wire  _GEN_6881 = 5'hc == rob_head ? rob_bsy_12 : _GEN_6880; // @[rob.scala 404:{43,43}]
  wire  _GEN_6882 = 5'hd == rob_head ? rob_bsy_13 : _GEN_6881; // @[rob.scala 404:{43,43}]
  wire  _GEN_6883 = 5'he == rob_head ? rob_bsy_14 : _GEN_6882; // @[rob.scala 404:{43,43}]
  wire  _GEN_6884 = 5'hf == rob_head ? rob_bsy_15 : _GEN_6883; // @[rob.scala 404:{43,43}]
  wire  _GEN_6885 = 5'h10 == rob_head ? rob_bsy_16 : _GEN_6884; // @[rob.scala 404:{43,43}]
  wire  _GEN_6886 = 5'h11 == rob_head ? rob_bsy_17 : _GEN_6885; // @[rob.scala 404:{43,43}]
  wire  _GEN_6887 = 5'h12 == rob_head ? rob_bsy_18 : _GEN_6886; // @[rob.scala 404:{43,43}]
  wire  _GEN_6888 = 5'h13 == rob_head ? rob_bsy_19 : _GEN_6887; // @[rob.scala 404:{43,43}]
  wire  _GEN_6889 = 5'h14 == rob_head ? rob_bsy_20 : _GEN_6888; // @[rob.scala 404:{43,43}]
  wire  _GEN_6890 = 5'h15 == rob_head ? rob_bsy_21 : _GEN_6889; // @[rob.scala 404:{43,43}]
  wire  _GEN_6891 = 5'h16 == rob_head ? rob_bsy_22 : _GEN_6890; // @[rob.scala 404:{43,43}]
  wire  _GEN_6892 = 5'h17 == rob_head ? rob_bsy_23 : _GEN_6891; // @[rob.scala 404:{43,43}]
  wire  _GEN_6893 = 5'h18 == rob_head ? rob_bsy_24 : _GEN_6892; // @[rob.scala 404:{43,43}]
  wire  _GEN_6894 = 5'h19 == rob_head ? rob_bsy_25 : _GEN_6893; // @[rob.scala 404:{43,43}]
  wire  _GEN_6895 = 5'h1a == rob_head ? rob_bsy_26 : _GEN_6894; // @[rob.scala 404:{43,43}]
  wire  _GEN_6896 = 5'h1b == rob_head ? rob_bsy_27 : _GEN_6895; // @[rob.scala 404:{43,43}]
  wire  _GEN_6897 = 5'h1c == rob_head ? rob_bsy_28 : _GEN_6896; // @[rob.scala 404:{43,43}]
  wire  _GEN_6898 = 5'h1d == rob_head ? rob_bsy_29 : _GEN_6897; // @[rob.scala 404:{43,43}]
  wire  _GEN_6899 = 5'h1e == rob_head ? rob_bsy_30 : _GEN_6898; // @[rob.scala 404:{43,43}]
  wire  _GEN_6900 = 5'h1f == rob_head ? rob_bsy_31 : _GEN_6899; // @[rob.scala 404:{43,43}]
  wire  can_commit_0 = rob_head_vals_0 & ~_GEN_6900 & ~io_csr_stall; // @[rob.scala 404:64]
  reg  rob_exception_31; // @[rob.scala 311:28]
  reg  rob_exception_30; // @[rob.scala 311:28]
  reg  rob_exception_29; // @[rob.scala 311:28]
  reg  rob_exception_28; // @[rob.scala 311:28]
  reg  rob_exception_27; // @[rob.scala 311:28]
  reg  rob_exception_26; // @[rob.scala 311:28]
  reg  rob_exception_25; // @[rob.scala 311:28]
  reg  rob_exception_24; // @[rob.scala 311:28]
  reg  rob_exception_23; // @[rob.scala 311:28]
  reg  rob_exception_22; // @[rob.scala 311:28]
  reg  rob_exception_21; // @[rob.scala 311:28]
  reg  rob_exception_20; // @[rob.scala 311:28]
  reg  rob_exception_19; // @[rob.scala 311:28]
  reg  rob_exception_18; // @[rob.scala 311:28]
  reg  rob_exception_17; // @[rob.scala 311:28]
  reg  rob_exception_16; // @[rob.scala 311:28]
  reg  rob_exception_15; // @[rob.scala 311:28]
  reg  rob_exception_14; // @[rob.scala 311:28]
  reg  rob_exception_13; // @[rob.scala 311:28]
  reg  rob_exception_12; // @[rob.scala 311:28]
  reg  rob_exception_11; // @[rob.scala 311:28]
  reg  rob_exception_10; // @[rob.scala 311:28]
  reg  rob_exception_9; // @[rob.scala 311:28]
  reg  rob_exception_8; // @[rob.scala 311:28]
  reg  rob_exception_7; // @[rob.scala 311:28]
  reg  rob_exception_6; // @[rob.scala 311:28]
  reg  rob_exception_5; // @[rob.scala 311:28]
  reg  rob_exception_4; // @[rob.scala 311:28]
  reg  rob_exception_3; // @[rob.scala 311:28]
  reg  rob_exception_2; // @[rob.scala 311:28]
  reg  rob_exception_1; // @[rob.scala 311:28]
  reg  rob_exception_0; // @[rob.scala 311:28]
  wire  _GEN_6838 = 5'h1 == rob_head ? rob_exception_1 : rob_exception_0; // @[rob.scala 398:{49,49}]
  wire  _GEN_6839 = 5'h2 == rob_head ? rob_exception_2 : _GEN_6838; // @[rob.scala 398:{49,49}]
  wire  _GEN_6840 = 5'h3 == rob_head ? rob_exception_3 : _GEN_6839; // @[rob.scala 398:{49,49}]
  wire  _GEN_6841 = 5'h4 == rob_head ? rob_exception_4 : _GEN_6840; // @[rob.scala 398:{49,49}]
  wire  _GEN_6842 = 5'h5 == rob_head ? rob_exception_5 : _GEN_6841; // @[rob.scala 398:{49,49}]
  wire  _GEN_6843 = 5'h6 == rob_head ? rob_exception_6 : _GEN_6842; // @[rob.scala 398:{49,49}]
  wire  _GEN_6844 = 5'h7 == rob_head ? rob_exception_7 : _GEN_6843; // @[rob.scala 398:{49,49}]
  wire  _GEN_6845 = 5'h8 == rob_head ? rob_exception_8 : _GEN_6844; // @[rob.scala 398:{49,49}]
  wire  _GEN_6846 = 5'h9 == rob_head ? rob_exception_9 : _GEN_6845; // @[rob.scala 398:{49,49}]
  wire  _GEN_6847 = 5'ha == rob_head ? rob_exception_10 : _GEN_6846; // @[rob.scala 398:{49,49}]
  wire  _GEN_6848 = 5'hb == rob_head ? rob_exception_11 : _GEN_6847; // @[rob.scala 398:{49,49}]
  wire  _GEN_6849 = 5'hc == rob_head ? rob_exception_12 : _GEN_6848; // @[rob.scala 398:{49,49}]
  wire  _GEN_6850 = 5'hd == rob_head ? rob_exception_13 : _GEN_6849; // @[rob.scala 398:{49,49}]
  wire  _GEN_6851 = 5'he == rob_head ? rob_exception_14 : _GEN_6850; // @[rob.scala 398:{49,49}]
  wire  _GEN_6852 = 5'hf == rob_head ? rob_exception_15 : _GEN_6851; // @[rob.scala 398:{49,49}]
  wire  _GEN_6853 = 5'h10 == rob_head ? rob_exception_16 : _GEN_6852; // @[rob.scala 398:{49,49}]
  wire  _GEN_6854 = 5'h11 == rob_head ? rob_exception_17 : _GEN_6853; // @[rob.scala 398:{49,49}]
  wire  _GEN_6855 = 5'h12 == rob_head ? rob_exception_18 : _GEN_6854; // @[rob.scala 398:{49,49}]
  wire  _GEN_6856 = 5'h13 == rob_head ? rob_exception_19 : _GEN_6855; // @[rob.scala 398:{49,49}]
  wire  _GEN_6857 = 5'h14 == rob_head ? rob_exception_20 : _GEN_6856; // @[rob.scala 398:{49,49}]
  wire  _GEN_6858 = 5'h15 == rob_head ? rob_exception_21 : _GEN_6857; // @[rob.scala 398:{49,49}]
  wire  _GEN_6859 = 5'h16 == rob_head ? rob_exception_22 : _GEN_6858; // @[rob.scala 398:{49,49}]
  wire  _GEN_6860 = 5'h17 == rob_head ? rob_exception_23 : _GEN_6859; // @[rob.scala 398:{49,49}]
  wire  _GEN_6861 = 5'h18 == rob_head ? rob_exception_24 : _GEN_6860; // @[rob.scala 398:{49,49}]
  wire  _GEN_6862 = 5'h19 == rob_head ? rob_exception_25 : _GEN_6861; // @[rob.scala 398:{49,49}]
  wire  _GEN_6863 = 5'h1a == rob_head ? rob_exception_26 : _GEN_6862; // @[rob.scala 398:{49,49}]
  wire  _GEN_6864 = 5'h1b == rob_head ? rob_exception_27 : _GEN_6863; // @[rob.scala 398:{49,49}]
  wire  _GEN_6865 = 5'h1c == rob_head ? rob_exception_28 : _GEN_6864; // @[rob.scala 398:{49,49}]
  wire  _GEN_6866 = 5'h1d == rob_head ? rob_exception_29 : _GEN_6865; // @[rob.scala 398:{49,49}]
  wire  _GEN_6867 = 5'h1e == rob_head ? rob_exception_30 : _GEN_6866; // @[rob.scala 398:{49,49}]
  wire  _GEN_6868 = 5'h1f == rob_head ? rob_exception_31 : _GEN_6867; // @[rob.scala 398:{49,49}]
  wire  can_throw_exception_0 = rob_head_vals_0 & _GEN_6868; // @[rob.scala 398:49]
  wire  _T_414 = can_commit_0 & ~can_throw_exception_0; // @[rob.scala 547:43]
  reg  _T_404; // @[rob.scala 540:94]
  reg  _T_407; // @[rob.scala 540:123]
  wire  _T_408 = rob_state != 2'h1 & rob_state != 2'h3 | _T_404 | _T_407; // @[rob.scala 540:113]
  wire  _T_415 = ~_T_408; // @[rob.scala 547:73]
  wire  will_commit_0 = can_commit_0 & ~can_throw_exception_0 & ~_T_408; // @[rob.scala 547:70]
  reg  rob_unsafe_0; // @[rob.scala 309:28]
  reg  rob_unsafe_1; // @[rob.scala 309:28]
  reg  rob_unsafe_2; // @[rob.scala 309:28]
  reg  rob_unsafe_3; // @[rob.scala 309:28]
  reg  rob_unsafe_4; // @[rob.scala 309:28]
  reg  rob_unsafe_5; // @[rob.scala 309:28]
  reg  rob_unsafe_6; // @[rob.scala 309:28]
  reg  rob_unsafe_7; // @[rob.scala 309:28]
  reg  rob_unsafe_8; // @[rob.scala 309:28]
  reg  rob_unsafe_9; // @[rob.scala 309:28]
  reg  rob_unsafe_10; // @[rob.scala 309:28]
  reg  rob_unsafe_11; // @[rob.scala 309:28]
  reg  rob_unsafe_12; // @[rob.scala 309:28]
  reg  rob_unsafe_13; // @[rob.scala 309:28]
  reg  rob_unsafe_14; // @[rob.scala 309:28]
  reg  rob_unsafe_15; // @[rob.scala 309:28]
  reg  rob_unsafe_16; // @[rob.scala 309:28]
  reg  rob_unsafe_17; // @[rob.scala 309:28]
  reg  rob_unsafe_18; // @[rob.scala 309:28]
  reg  rob_unsafe_19; // @[rob.scala 309:28]
  reg  rob_unsafe_20; // @[rob.scala 309:28]
  reg  rob_unsafe_21; // @[rob.scala 309:28]
  reg  rob_unsafe_22; // @[rob.scala 309:28]
  reg  rob_unsafe_23; // @[rob.scala 309:28]
  reg  rob_unsafe_24; // @[rob.scala 309:28]
  reg  rob_unsafe_25; // @[rob.scala 309:28]
  reg  rob_unsafe_26; // @[rob.scala 309:28]
  reg  rob_unsafe_27; // @[rob.scala 309:28]
  reg  rob_unsafe_28; // @[rob.scala 309:28]
  reg  rob_unsafe_29; // @[rob.scala 309:28]
  reg  rob_unsafe_30; // @[rob.scala 309:28]
  reg  rob_unsafe_31; // @[rob.scala 309:28]
  reg [6:0] rob_uop_0_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_0_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_0_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_0_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_0_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_0_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_0_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_0_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_0_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_0_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_0_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_0_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_0_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_0_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_0_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_0_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_0_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_0_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_0_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_0_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_0_is_br; // @[rob.scala 310:28]
  reg  rob_uop_0_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_0_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_0_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_0_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_0_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_0_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_0_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_0_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_0_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_0_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_0_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_0_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_0_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_0_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_0_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_0_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_0_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_0_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_0_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_0_ppred; // @[rob.scala 310:28]
  reg  rob_uop_0_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_0_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_0_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_0_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_0_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_0_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_0_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_0_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_0_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_0_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_0_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_0_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_0_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_0_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_0_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_0_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_0_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_0_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_0_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_0_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_0_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_0_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_0_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_0_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_0_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_0_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_0_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_0_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_0_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_0_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_0_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_0_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_0_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_0_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_0_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_0_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_0_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_0_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_1_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_1_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_1_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_1_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_1_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_1_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_1_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_1_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_1_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_1_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_1_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_1_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_1_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_1_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_1_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_1_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_1_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_1_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_1_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_1_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_1_is_br; // @[rob.scala 310:28]
  reg  rob_uop_1_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_1_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_1_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_1_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_1_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_1_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_1_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_1_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_1_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_1_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_1_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_1_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_1_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_1_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_1_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_1_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_1_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_1_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_1_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_1_ppred; // @[rob.scala 310:28]
  reg  rob_uop_1_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_1_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_1_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_1_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_1_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_1_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_1_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_1_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_1_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_1_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_1_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_1_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_1_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_1_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_1_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_1_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_1_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_1_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_1_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_1_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_1_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_1_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_1_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_1_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_1_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_1_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_1_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_1_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_1_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_1_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_1_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_1_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_1_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_1_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_1_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_1_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_1_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_1_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_2_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_2_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_2_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_2_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_2_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_2_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_2_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_2_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_2_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_2_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_2_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_2_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_2_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_2_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_2_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_2_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_2_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_2_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_2_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_2_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_2_is_br; // @[rob.scala 310:28]
  reg  rob_uop_2_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_2_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_2_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_2_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_2_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_2_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_2_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_2_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_2_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_2_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_2_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_2_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_2_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_2_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_2_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_2_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_2_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_2_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_2_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_2_ppred; // @[rob.scala 310:28]
  reg  rob_uop_2_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_2_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_2_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_2_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_2_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_2_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_2_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_2_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_2_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_2_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_2_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_2_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_2_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_2_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_2_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_2_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_2_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_2_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_2_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_2_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_2_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_2_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_2_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_2_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_2_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_2_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_2_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_2_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_2_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_2_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_2_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_2_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_2_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_2_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_2_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_2_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_2_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_2_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_3_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_3_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_3_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_3_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_3_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_3_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_3_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_3_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_3_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_3_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_3_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_3_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_3_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_3_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_3_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_3_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_3_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_3_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_3_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_3_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_3_is_br; // @[rob.scala 310:28]
  reg  rob_uop_3_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_3_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_3_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_3_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_3_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_3_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_3_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_3_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_3_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_3_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_3_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_3_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_3_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_3_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_3_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_3_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_3_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_3_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_3_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_3_ppred; // @[rob.scala 310:28]
  reg  rob_uop_3_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_3_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_3_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_3_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_3_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_3_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_3_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_3_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_3_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_3_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_3_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_3_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_3_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_3_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_3_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_3_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_3_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_3_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_3_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_3_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_3_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_3_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_3_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_3_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_3_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_3_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_3_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_3_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_3_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_3_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_3_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_3_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_3_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_3_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_3_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_3_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_3_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_3_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_4_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_4_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_4_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_4_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_4_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_4_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_4_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_4_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_4_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_4_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_4_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_4_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_4_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_4_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_4_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_4_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_4_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_4_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_4_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_4_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_4_is_br; // @[rob.scala 310:28]
  reg  rob_uop_4_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_4_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_4_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_4_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_4_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_4_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_4_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_4_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_4_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_4_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_4_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_4_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_4_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_4_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_4_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_4_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_4_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_4_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_4_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_4_ppred; // @[rob.scala 310:28]
  reg  rob_uop_4_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_4_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_4_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_4_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_4_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_4_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_4_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_4_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_4_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_4_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_4_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_4_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_4_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_4_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_4_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_4_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_4_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_4_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_4_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_4_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_4_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_4_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_4_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_4_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_4_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_4_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_4_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_4_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_4_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_4_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_4_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_4_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_4_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_4_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_4_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_4_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_4_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_4_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_5_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_5_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_5_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_5_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_5_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_5_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_5_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_5_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_5_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_5_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_5_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_5_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_5_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_5_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_5_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_5_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_5_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_5_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_5_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_5_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_5_is_br; // @[rob.scala 310:28]
  reg  rob_uop_5_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_5_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_5_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_5_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_5_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_5_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_5_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_5_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_5_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_5_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_5_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_5_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_5_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_5_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_5_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_5_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_5_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_5_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_5_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_5_ppred; // @[rob.scala 310:28]
  reg  rob_uop_5_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_5_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_5_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_5_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_5_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_5_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_5_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_5_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_5_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_5_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_5_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_5_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_5_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_5_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_5_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_5_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_5_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_5_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_5_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_5_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_5_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_5_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_5_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_5_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_5_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_5_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_5_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_5_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_5_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_5_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_5_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_5_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_5_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_5_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_5_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_5_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_5_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_5_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_6_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_6_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_6_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_6_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_6_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_6_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_6_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_6_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_6_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_6_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_6_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_6_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_6_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_6_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_6_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_6_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_6_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_6_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_6_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_6_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_6_is_br; // @[rob.scala 310:28]
  reg  rob_uop_6_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_6_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_6_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_6_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_6_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_6_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_6_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_6_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_6_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_6_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_6_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_6_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_6_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_6_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_6_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_6_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_6_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_6_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_6_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_6_ppred; // @[rob.scala 310:28]
  reg  rob_uop_6_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_6_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_6_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_6_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_6_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_6_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_6_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_6_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_6_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_6_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_6_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_6_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_6_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_6_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_6_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_6_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_6_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_6_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_6_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_6_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_6_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_6_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_6_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_6_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_6_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_6_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_6_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_6_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_6_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_6_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_6_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_6_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_6_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_6_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_6_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_6_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_6_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_6_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_7_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_7_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_7_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_7_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_7_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_7_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_7_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_7_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_7_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_7_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_7_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_7_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_7_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_7_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_7_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_7_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_7_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_7_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_7_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_7_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_7_is_br; // @[rob.scala 310:28]
  reg  rob_uop_7_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_7_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_7_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_7_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_7_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_7_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_7_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_7_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_7_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_7_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_7_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_7_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_7_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_7_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_7_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_7_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_7_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_7_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_7_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_7_ppred; // @[rob.scala 310:28]
  reg  rob_uop_7_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_7_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_7_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_7_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_7_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_7_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_7_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_7_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_7_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_7_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_7_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_7_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_7_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_7_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_7_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_7_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_7_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_7_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_7_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_7_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_7_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_7_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_7_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_7_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_7_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_7_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_7_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_7_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_7_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_7_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_7_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_7_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_7_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_7_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_7_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_7_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_7_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_7_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_8_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_8_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_8_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_8_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_8_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_8_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_8_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_8_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_8_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_8_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_8_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_8_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_8_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_8_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_8_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_8_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_8_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_8_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_8_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_8_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_8_is_br; // @[rob.scala 310:28]
  reg  rob_uop_8_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_8_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_8_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_8_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_8_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_8_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_8_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_8_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_8_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_8_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_8_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_8_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_8_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_8_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_8_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_8_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_8_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_8_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_8_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_8_ppred; // @[rob.scala 310:28]
  reg  rob_uop_8_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_8_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_8_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_8_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_8_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_8_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_8_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_8_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_8_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_8_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_8_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_8_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_8_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_8_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_8_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_8_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_8_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_8_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_8_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_8_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_8_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_8_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_8_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_8_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_8_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_8_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_8_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_8_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_8_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_8_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_8_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_8_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_8_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_8_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_8_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_8_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_8_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_8_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_9_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_9_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_9_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_9_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_9_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_9_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_9_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_9_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_9_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_9_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_9_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_9_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_9_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_9_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_9_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_9_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_9_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_9_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_9_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_9_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_9_is_br; // @[rob.scala 310:28]
  reg  rob_uop_9_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_9_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_9_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_9_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_9_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_9_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_9_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_9_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_9_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_9_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_9_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_9_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_9_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_9_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_9_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_9_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_9_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_9_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_9_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_9_ppred; // @[rob.scala 310:28]
  reg  rob_uop_9_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_9_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_9_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_9_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_9_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_9_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_9_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_9_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_9_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_9_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_9_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_9_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_9_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_9_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_9_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_9_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_9_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_9_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_9_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_9_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_9_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_9_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_9_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_9_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_9_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_9_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_9_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_9_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_9_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_9_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_9_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_9_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_9_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_9_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_9_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_9_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_9_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_9_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_10_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_10_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_10_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_10_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_10_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_10_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_10_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_10_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_10_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_10_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_10_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_10_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_10_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_10_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_10_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_10_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_10_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_10_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_10_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_10_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_10_is_br; // @[rob.scala 310:28]
  reg  rob_uop_10_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_10_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_10_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_10_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_10_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_10_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_10_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_10_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_10_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_10_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_10_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_10_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_10_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_10_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_10_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_10_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_10_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_10_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_10_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_10_ppred; // @[rob.scala 310:28]
  reg  rob_uop_10_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_10_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_10_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_10_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_10_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_10_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_10_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_10_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_10_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_10_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_10_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_10_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_10_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_10_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_10_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_10_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_10_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_10_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_10_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_10_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_10_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_10_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_10_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_10_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_10_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_10_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_10_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_10_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_10_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_10_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_10_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_10_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_10_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_10_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_10_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_10_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_10_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_10_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_11_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_11_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_11_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_11_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_11_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_11_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_11_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_11_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_11_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_11_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_11_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_11_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_11_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_11_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_11_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_11_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_11_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_11_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_11_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_11_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_11_is_br; // @[rob.scala 310:28]
  reg  rob_uop_11_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_11_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_11_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_11_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_11_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_11_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_11_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_11_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_11_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_11_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_11_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_11_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_11_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_11_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_11_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_11_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_11_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_11_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_11_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_11_ppred; // @[rob.scala 310:28]
  reg  rob_uop_11_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_11_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_11_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_11_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_11_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_11_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_11_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_11_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_11_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_11_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_11_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_11_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_11_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_11_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_11_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_11_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_11_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_11_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_11_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_11_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_11_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_11_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_11_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_11_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_11_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_11_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_11_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_11_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_11_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_11_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_11_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_11_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_11_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_11_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_11_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_11_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_11_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_11_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_12_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_12_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_12_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_12_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_12_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_12_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_12_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_12_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_12_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_12_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_12_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_12_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_12_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_12_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_12_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_12_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_12_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_12_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_12_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_12_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_12_is_br; // @[rob.scala 310:28]
  reg  rob_uop_12_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_12_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_12_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_12_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_12_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_12_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_12_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_12_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_12_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_12_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_12_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_12_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_12_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_12_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_12_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_12_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_12_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_12_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_12_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_12_ppred; // @[rob.scala 310:28]
  reg  rob_uop_12_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_12_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_12_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_12_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_12_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_12_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_12_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_12_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_12_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_12_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_12_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_12_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_12_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_12_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_12_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_12_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_12_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_12_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_12_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_12_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_12_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_12_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_12_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_12_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_12_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_12_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_12_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_12_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_12_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_12_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_12_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_12_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_12_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_12_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_12_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_12_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_12_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_12_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_13_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_13_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_13_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_13_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_13_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_13_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_13_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_13_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_13_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_13_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_13_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_13_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_13_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_13_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_13_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_13_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_13_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_13_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_13_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_13_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_13_is_br; // @[rob.scala 310:28]
  reg  rob_uop_13_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_13_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_13_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_13_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_13_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_13_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_13_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_13_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_13_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_13_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_13_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_13_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_13_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_13_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_13_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_13_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_13_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_13_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_13_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_13_ppred; // @[rob.scala 310:28]
  reg  rob_uop_13_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_13_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_13_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_13_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_13_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_13_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_13_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_13_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_13_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_13_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_13_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_13_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_13_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_13_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_13_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_13_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_13_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_13_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_13_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_13_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_13_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_13_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_13_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_13_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_13_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_13_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_13_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_13_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_13_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_13_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_13_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_13_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_13_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_13_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_13_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_13_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_13_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_13_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_14_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_14_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_14_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_14_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_14_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_14_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_14_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_14_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_14_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_14_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_14_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_14_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_14_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_14_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_14_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_14_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_14_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_14_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_14_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_14_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_14_is_br; // @[rob.scala 310:28]
  reg  rob_uop_14_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_14_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_14_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_14_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_14_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_14_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_14_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_14_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_14_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_14_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_14_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_14_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_14_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_14_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_14_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_14_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_14_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_14_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_14_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_14_ppred; // @[rob.scala 310:28]
  reg  rob_uop_14_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_14_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_14_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_14_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_14_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_14_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_14_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_14_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_14_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_14_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_14_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_14_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_14_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_14_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_14_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_14_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_14_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_14_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_14_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_14_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_14_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_14_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_14_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_14_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_14_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_14_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_14_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_14_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_14_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_14_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_14_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_14_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_14_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_14_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_14_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_14_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_14_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_14_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_15_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_15_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_15_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_15_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_15_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_15_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_15_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_15_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_15_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_15_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_15_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_15_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_15_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_15_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_15_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_15_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_15_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_15_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_15_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_15_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_15_is_br; // @[rob.scala 310:28]
  reg  rob_uop_15_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_15_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_15_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_15_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_15_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_15_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_15_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_15_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_15_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_15_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_15_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_15_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_15_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_15_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_15_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_15_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_15_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_15_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_15_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_15_ppred; // @[rob.scala 310:28]
  reg  rob_uop_15_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_15_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_15_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_15_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_15_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_15_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_15_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_15_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_15_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_15_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_15_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_15_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_15_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_15_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_15_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_15_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_15_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_15_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_15_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_15_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_15_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_15_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_15_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_15_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_15_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_15_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_15_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_15_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_15_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_15_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_15_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_15_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_15_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_15_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_15_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_15_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_15_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_15_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_16_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_16_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_16_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_16_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_16_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_16_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_16_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_16_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_16_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_16_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_16_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_16_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_16_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_16_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_16_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_16_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_16_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_16_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_16_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_16_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_16_is_br; // @[rob.scala 310:28]
  reg  rob_uop_16_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_16_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_16_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_16_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_16_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_16_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_16_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_16_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_16_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_16_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_16_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_16_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_16_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_16_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_16_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_16_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_16_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_16_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_16_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_16_ppred; // @[rob.scala 310:28]
  reg  rob_uop_16_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_16_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_16_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_16_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_16_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_16_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_16_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_16_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_16_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_16_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_16_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_16_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_16_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_16_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_16_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_16_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_16_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_16_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_16_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_16_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_16_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_16_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_16_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_16_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_16_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_16_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_16_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_16_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_16_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_16_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_16_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_16_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_16_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_16_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_16_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_16_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_16_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_16_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_17_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_17_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_17_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_17_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_17_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_17_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_17_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_17_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_17_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_17_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_17_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_17_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_17_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_17_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_17_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_17_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_17_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_17_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_17_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_17_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_17_is_br; // @[rob.scala 310:28]
  reg  rob_uop_17_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_17_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_17_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_17_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_17_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_17_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_17_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_17_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_17_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_17_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_17_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_17_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_17_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_17_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_17_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_17_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_17_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_17_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_17_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_17_ppred; // @[rob.scala 310:28]
  reg  rob_uop_17_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_17_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_17_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_17_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_17_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_17_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_17_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_17_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_17_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_17_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_17_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_17_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_17_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_17_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_17_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_17_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_17_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_17_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_17_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_17_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_17_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_17_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_17_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_17_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_17_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_17_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_17_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_17_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_17_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_17_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_17_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_17_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_17_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_17_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_17_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_17_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_17_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_17_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_18_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_18_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_18_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_18_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_18_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_18_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_18_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_18_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_18_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_18_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_18_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_18_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_18_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_18_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_18_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_18_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_18_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_18_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_18_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_18_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_18_is_br; // @[rob.scala 310:28]
  reg  rob_uop_18_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_18_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_18_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_18_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_18_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_18_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_18_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_18_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_18_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_18_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_18_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_18_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_18_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_18_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_18_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_18_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_18_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_18_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_18_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_18_ppred; // @[rob.scala 310:28]
  reg  rob_uop_18_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_18_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_18_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_18_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_18_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_18_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_18_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_18_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_18_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_18_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_18_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_18_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_18_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_18_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_18_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_18_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_18_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_18_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_18_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_18_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_18_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_18_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_18_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_18_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_18_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_18_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_18_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_18_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_18_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_18_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_18_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_18_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_18_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_18_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_18_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_18_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_18_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_18_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_19_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_19_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_19_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_19_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_19_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_19_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_19_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_19_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_19_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_19_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_19_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_19_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_19_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_19_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_19_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_19_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_19_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_19_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_19_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_19_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_19_is_br; // @[rob.scala 310:28]
  reg  rob_uop_19_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_19_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_19_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_19_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_19_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_19_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_19_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_19_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_19_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_19_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_19_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_19_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_19_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_19_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_19_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_19_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_19_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_19_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_19_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_19_ppred; // @[rob.scala 310:28]
  reg  rob_uop_19_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_19_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_19_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_19_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_19_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_19_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_19_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_19_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_19_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_19_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_19_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_19_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_19_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_19_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_19_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_19_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_19_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_19_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_19_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_19_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_19_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_19_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_19_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_19_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_19_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_19_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_19_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_19_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_19_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_19_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_19_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_19_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_19_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_19_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_19_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_19_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_19_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_19_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_20_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_20_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_20_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_20_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_20_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_20_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_20_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_20_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_20_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_20_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_20_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_20_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_20_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_20_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_20_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_20_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_20_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_20_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_20_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_20_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_20_is_br; // @[rob.scala 310:28]
  reg  rob_uop_20_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_20_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_20_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_20_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_20_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_20_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_20_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_20_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_20_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_20_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_20_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_20_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_20_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_20_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_20_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_20_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_20_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_20_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_20_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_20_ppred; // @[rob.scala 310:28]
  reg  rob_uop_20_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_20_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_20_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_20_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_20_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_20_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_20_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_20_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_20_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_20_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_20_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_20_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_20_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_20_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_20_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_20_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_20_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_20_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_20_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_20_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_20_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_20_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_20_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_20_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_20_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_20_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_20_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_20_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_20_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_20_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_20_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_20_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_20_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_20_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_20_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_20_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_20_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_20_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_21_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_21_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_21_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_21_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_21_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_21_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_21_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_21_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_21_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_21_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_21_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_21_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_21_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_21_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_21_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_21_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_21_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_21_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_21_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_21_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_21_is_br; // @[rob.scala 310:28]
  reg  rob_uop_21_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_21_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_21_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_21_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_21_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_21_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_21_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_21_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_21_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_21_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_21_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_21_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_21_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_21_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_21_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_21_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_21_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_21_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_21_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_21_ppred; // @[rob.scala 310:28]
  reg  rob_uop_21_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_21_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_21_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_21_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_21_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_21_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_21_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_21_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_21_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_21_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_21_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_21_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_21_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_21_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_21_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_21_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_21_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_21_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_21_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_21_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_21_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_21_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_21_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_21_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_21_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_21_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_21_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_21_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_21_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_21_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_21_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_21_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_21_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_21_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_21_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_21_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_21_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_21_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_22_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_22_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_22_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_22_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_22_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_22_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_22_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_22_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_22_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_22_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_22_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_22_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_22_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_22_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_22_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_22_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_22_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_22_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_22_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_22_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_22_is_br; // @[rob.scala 310:28]
  reg  rob_uop_22_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_22_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_22_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_22_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_22_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_22_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_22_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_22_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_22_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_22_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_22_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_22_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_22_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_22_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_22_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_22_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_22_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_22_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_22_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_22_ppred; // @[rob.scala 310:28]
  reg  rob_uop_22_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_22_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_22_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_22_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_22_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_22_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_22_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_22_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_22_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_22_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_22_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_22_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_22_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_22_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_22_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_22_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_22_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_22_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_22_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_22_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_22_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_22_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_22_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_22_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_22_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_22_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_22_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_22_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_22_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_22_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_22_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_22_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_22_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_22_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_22_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_22_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_22_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_22_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_23_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_23_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_23_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_23_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_23_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_23_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_23_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_23_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_23_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_23_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_23_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_23_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_23_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_23_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_23_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_23_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_23_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_23_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_23_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_23_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_23_is_br; // @[rob.scala 310:28]
  reg  rob_uop_23_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_23_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_23_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_23_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_23_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_23_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_23_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_23_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_23_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_23_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_23_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_23_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_23_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_23_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_23_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_23_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_23_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_23_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_23_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_23_ppred; // @[rob.scala 310:28]
  reg  rob_uop_23_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_23_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_23_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_23_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_23_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_23_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_23_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_23_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_23_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_23_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_23_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_23_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_23_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_23_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_23_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_23_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_23_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_23_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_23_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_23_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_23_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_23_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_23_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_23_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_23_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_23_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_23_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_23_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_23_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_23_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_23_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_23_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_23_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_23_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_23_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_23_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_23_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_23_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_24_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_24_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_24_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_24_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_24_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_24_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_24_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_24_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_24_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_24_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_24_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_24_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_24_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_24_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_24_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_24_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_24_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_24_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_24_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_24_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_24_is_br; // @[rob.scala 310:28]
  reg  rob_uop_24_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_24_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_24_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_24_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_24_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_24_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_24_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_24_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_24_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_24_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_24_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_24_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_24_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_24_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_24_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_24_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_24_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_24_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_24_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_24_ppred; // @[rob.scala 310:28]
  reg  rob_uop_24_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_24_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_24_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_24_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_24_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_24_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_24_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_24_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_24_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_24_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_24_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_24_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_24_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_24_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_24_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_24_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_24_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_24_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_24_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_24_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_24_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_24_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_24_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_24_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_24_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_24_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_24_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_24_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_24_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_24_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_24_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_24_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_24_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_24_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_24_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_24_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_24_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_24_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_25_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_25_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_25_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_25_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_25_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_25_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_25_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_25_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_25_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_25_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_25_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_25_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_25_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_25_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_25_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_25_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_25_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_25_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_25_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_25_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_25_is_br; // @[rob.scala 310:28]
  reg  rob_uop_25_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_25_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_25_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_25_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_25_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_25_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_25_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_25_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_25_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_25_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_25_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_25_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_25_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_25_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_25_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_25_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_25_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_25_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_25_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_25_ppred; // @[rob.scala 310:28]
  reg  rob_uop_25_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_25_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_25_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_25_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_25_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_25_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_25_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_25_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_25_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_25_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_25_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_25_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_25_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_25_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_25_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_25_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_25_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_25_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_25_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_25_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_25_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_25_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_25_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_25_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_25_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_25_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_25_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_25_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_25_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_25_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_25_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_25_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_25_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_25_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_25_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_25_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_25_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_25_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_26_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_26_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_26_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_26_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_26_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_26_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_26_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_26_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_26_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_26_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_26_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_26_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_26_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_26_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_26_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_26_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_26_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_26_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_26_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_26_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_26_is_br; // @[rob.scala 310:28]
  reg  rob_uop_26_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_26_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_26_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_26_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_26_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_26_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_26_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_26_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_26_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_26_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_26_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_26_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_26_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_26_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_26_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_26_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_26_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_26_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_26_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_26_ppred; // @[rob.scala 310:28]
  reg  rob_uop_26_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_26_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_26_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_26_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_26_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_26_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_26_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_26_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_26_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_26_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_26_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_26_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_26_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_26_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_26_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_26_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_26_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_26_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_26_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_26_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_26_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_26_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_26_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_26_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_26_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_26_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_26_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_26_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_26_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_26_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_26_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_26_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_26_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_26_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_26_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_26_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_26_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_26_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_27_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_27_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_27_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_27_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_27_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_27_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_27_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_27_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_27_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_27_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_27_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_27_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_27_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_27_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_27_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_27_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_27_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_27_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_27_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_27_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_27_is_br; // @[rob.scala 310:28]
  reg  rob_uop_27_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_27_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_27_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_27_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_27_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_27_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_27_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_27_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_27_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_27_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_27_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_27_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_27_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_27_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_27_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_27_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_27_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_27_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_27_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_27_ppred; // @[rob.scala 310:28]
  reg  rob_uop_27_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_27_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_27_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_27_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_27_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_27_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_27_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_27_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_27_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_27_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_27_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_27_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_27_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_27_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_27_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_27_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_27_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_27_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_27_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_27_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_27_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_27_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_27_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_27_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_27_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_27_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_27_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_27_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_27_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_27_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_27_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_27_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_27_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_27_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_27_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_27_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_27_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_27_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_28_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_28_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_28_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_28_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_28_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_28_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_28_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_28_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_28_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_28_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_28_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_28_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_28_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_28_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_28_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_28_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_28_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_28_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_28_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_28_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_28_is_br; // @[rob.scala 310:28]
  reg  rob_uop_28_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_28_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_28_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_28_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_28_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_28_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_28_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_28_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_28_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_28_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_28_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_28_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_28_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_28_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_28_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_28_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_28_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_28_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_28_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_28_ppred; // @[rob.scala 310:28]
  reg  rob_uop_28_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_28_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_28_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_28_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_28_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_28_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_28_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_28_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_28_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_28_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_28_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_28_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_28_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_28_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_28_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_28_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_28_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_28_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_28_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_28_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_28_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_28_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_28_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_28_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_28_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_28_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_28_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_28_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_28_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_28_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_28_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_28_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_28_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_28_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_28_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_28_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_28_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_28_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_29_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_29_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_29_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_29_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_29_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_29_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_29_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_29_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_29_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_29_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_29_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_29_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_29_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_29_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_29_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_29_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_29_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_29_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_29_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_29_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_29_is_br; // @[rob.scala 310:28]
  reg  rob_uop_29_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_29_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_29_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_29_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_29_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_29_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_29_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_29_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_29_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_29_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_29_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_29_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_29_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_29_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_29_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_29_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_29_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_29_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_29_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_29_ppred; // @[rob.scala 310:28]
  reg  rob_uop_29_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_29_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_29_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_29_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_29_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_29_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_29_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_29_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_29_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_29_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_29_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_29_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_29_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_29_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_29_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_29_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_29_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_29_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_29_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_29_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_29_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_29_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_29_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_29_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_29_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_29_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_29_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_29_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_29_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_29_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_29_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_29_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_29_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_29_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_29_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_29_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_29_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_29_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_30_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_30_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_30_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_30_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_30_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_30_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_30_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_30_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_30_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_30_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_30_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_30_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_30_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_30_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_30_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_30_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_30_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_30_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_30_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_30_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_30_is_br; // @[rob.scala 310:28]
  reg  rob_uop_30_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_30_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_30_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_30_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_30_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_30_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_30_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_30_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_30_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_30_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_30_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_30_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_30_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_30_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_30_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_30_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_30_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_30_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_30_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_30_ppred; // @[rob.scala 310:28]
  reg  rob_uop_30_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_30_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_30_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_30_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_30_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_30_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_30_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_30_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_30_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_30_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_30_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_30_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_30_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_30_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_30_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_30_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_30_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_30_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_30_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_30_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_30_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_30_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_30_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_30_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_30_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_30_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_30_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_30_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_30_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_30_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_30_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_30_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_30_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_30_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_30_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_30_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_30_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_30_debug_tsrc; // @[rob.scala 310:28]
  reg [6:0] rob_uop_31_uopc; // @[rob.scala 310:28]
  reg [31:0] rob_uop_31_inst; // @[rob.scala 310:28]
  reg [31:0] rob_uop_31_debug_inst; // @[rob.scala 310:28]
  reg  rob_uop_31_is_rvc; // @[rob.scala 310:28]
  reg [39:0] rob_uop_31_debug_pc; // @[rob.scala 310:28]
  reg [2:0] rob_uop_31_iq_type; // @[rob.scala 310:28]
  reg [9:0] rob_uop_31_fu_code; // @[rob.scala 310:28]
  reg [3:0] rob_uop_31_ctrl_br_type; // @[rob.scala 310:28]
  reg [1:0] rob_uop_31_ctrl_op1_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_31_ctrl_op2_sel; // @[rob.scala 310:28]
  reg [2:0] rob_uop_31_ctrl_imm_sel; // @[rob.scala 310:28]
  reg [3:0] rob_uop_31_ctrl_op_fcn; // @[rob.scala 310:28]
  reg  rob_uop_31_ctrl_fcn_dw; // @[rob.scala 310:28]
  reg [2:0] rob_uop_31_ctrl_csr_cmd; // @[rob.scala 310:28]
  reg  rob_uop_31_ctrl_is_load; // @[rob.scala 310:28]
  reg  rob_uop_31_ctrl_is_sta; // @[rob.scala 310:28]
  reg  rob_uop_31_ctrl_is_std; // @[rob.scala 310:28]
  reg [1:0] rob_uop_31_iw_state; // @[rob.scala 310:28]
  reg  rob_uop_31_iw_p1_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_31_iw_p2_poisoned; // @[rob.scala 310:28]
  reg  rob_uop_31_is_br; // @[rob.scala 310:28]
  reg  rob_uop_31_is_jalr; // @[rob.scala 310:28]
  reg  rob_uop_31_is_jal; // @[rob.scala 310:28]
  reg  rob_uop_31_is_sfb; // @[rob.scala 310:28]
  reg [7:0] rob_uop_31_br_mask; // @[rob.scala 310:28]
  reg [2:0] rob_uop_31_br_tag; // @[rob.scala 310:28]
  reg [3:0] rob_uop_31_ftq_idx; // @[rob.scala 310:28]
  reg  rob_uop_31_edge_inst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_31_pc_lob; // @[rob.scala 310:28]
  reg  rob_uop_31_taken; // @[rob.scala 310:28]
  reg [19:0] rob_uop_31_imm_packed; // @[rob.scala 310:28]
  reg [11:0] rob_uop_31_csr_addr; // @[rob.scala 310:28]
  reg [4:0] rob_uop_31_rob_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_31_ldq_idx; // @[rob.scala 310:28]
  reg [2:0] rob_uop_31_stq_idx; // @[rob.scala 310:28]
  reg [1:0] rob_uop_31_rxq_idx; // @[rob.scala 310:28]
  reg [5:0] rob_uop_31_pdst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_31_prs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_31_prs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_31_prs3; // @[rob.scala 310:28]
  reg [3:0] rob_uop_31_ppred; // @[rob.scala 310:28]
  reg  rob_uop_31_prs1_busy; // @[rob.scala 310:28]
  reg  rob_uop_31_prs2_busy; // @[rob.scala 310:28]
  reg  rob_uop_31_prs3_busy; // @[rob.scala 310:28]
  reg  rob_uop_31_ppred_busy; // @[rob.scala 310:28]
  reg [5:0] rob_uop_31_stale_pdst; // @[rob.scala 310:28]
  reg  rob_uop_31_exception; // @[rob.scala 310:28]
  reg [63:0] rob_uop_31_exc_cause; // @[rob.scala 310:28]
  reg  rob_uop_31_bypassable; // @[rob.scala 310:28]
  reg [4:0] rob_uop_31_mem_cmd; // @[rob.scala 310:28]
  reg [1:0] rob_uop_31_mem_size; // @[rob.scala 310:28]
  reg  rob_uop_31_mem_signed; // @[rob.scala 310:28]
  reg  rob_uop_31_is_fence; // @[rob.scala 310:28]
  reg  rob_uop_31_is_fencei; // @[rob.scala 310:28]
  reg  rob_uop_31_is_amo; // @[rob.scala 310:28]
  reg  rob_uop_31_uses_ldq; // @[rob.scala 310:28]
  reg  rob_uop_31_uses_stq; // @[rob.scala 310:28]
  reg  rob_uop_31_is_sys_pc2epc; // @[rob.scala 310:28]
  reg  rob_uop_31_is_unique; // @[rob.scala 310:28]
  reg  rob_uop_31_flush_on_commit; // @[rob.scala 310:28]
  reg  rob_uop_31_ldst_is_rs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_31_ldst; // @[rob.scala 310:28]
  reg [5:0] rob_uop_31_lrs1; // @[rob.scala 310:28]
  reg [5:0] rob_uop_31_lrs2; // @[rob.scala 310:28]
  reg [5:0] rob_uop_31_lrs3; // @[rob.scala 310:28]
  reg  rob_uop_31_ldst_val; // @[rob.scala 310:28]
  reg [1:0] rob_uop_31_dst_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_31_lrs1_rtype; // @[rob.scala 310:28]
  reg [1:0] rob_uop_31_lrs2_rtype; // @[rob.scala 310:28]
  reg  rob_uop_31_frs3_en; // @[rob.scala 310:28]
  reg  rob_uop_31_fp_val; // @[rob.scala 310:28]
  reg  rob_uop_31_fp_single; // @[rob.scala 310:28]
  reg  rob_uop_31_xcpt_pf_if; // @[rob.scala 310:28]
  reg  rob_uop_31_xcpt_ae_if; // @[rob.scala 310:28]
  reg  rob_uop_31_xcpt_ma_if; // @[rob.scala 310:28]
  reg  rob_uop_31_bp_debug_if; // @[rob.scala 310:28]
  reg  rob_uop_31_bp_xcpt_if; // @[rob.scala 310:28]
  reg [1:0] rob_uop_31_debug_fsrc; // @[rob.scala 310:28]
  reg [1:0] rob_uop_31_debug_tsrc; // @[rob.scala 310:28]
  reg  rob_predicated_0; // @[rob.scala 312:29]
  reg  rob_predicated_1; // @[rob.scala 312:29]
  reg  rob_predicated_2; // @[rob.scala 312:29]
  reg  rob_predicated_3; // @[rob.scala 312:29]
  reg  rob_predicated_4; // @[rob.scala 312:29]
  reg  rob_predicated_5; // @[rob.scala 312:29]
  reg  rob_predicated_6; // @[rob.scala 312:29]
  reg  rob_predicated_7; // @[rob.scala 312:29]
  reg  rob_predicated_8; // @[rob.scala 312:29]
  reg  rob_predicated_9; // @[rob.scala 312:29]
  reg  rob_predicated_10; // @[rob.scala 312:29]
  reg  rob_predicated_11; // @[rob.scala 312:29]
  reg  rob_predicated_12; // @[rob.scala 312:29]
  reg  rob_predicated_13; // @[rob.scala 312:29]
  reg  rob_predicated_14; // @[rob.scala 312:29]
  reg  rob_predicated_15; // @[rob.scala 312:29]
  reg  rob_predicated_16; // @[rob.scala 312:29]
  reg  rob_predicated_17; // @[rob.scala 312:29]
  reg  rob_predicated_18; // @[rob.scala 312:29]
  reg  rob_predicated_19; // @[rob.scala 312:29]
  reg  rob_predicated_20; // @[rob.scala 312:29]
  reg  rob_predicated_21; // @[rob.scala 312:29]
  reg  rob_predicated_22; // @[rob.scala 312:29]
  reg  rob_predicated_23; // @[rob.scala 312:29]
  reg  rob_predicated_24; // @[rob.scala 312:29]
  reg  rob_predicated_25; // @[rob.scala 312:29]
  reg  rob_predicated_26; // @[rob.scala 312:29]
  reg  rob_predicated_27; // @[rob.scala 312:29]
  reg  rob_predicated_28; // @[rob.scala 312:29]
  reg  rob_predicated_29; // @[rob.scala 312:29]
  reg  rob_predicated_30; // @[rob.scala 312:29]
  reg  rob_predicated_31; // @[rob.scala 312:29]
  wire  _GEN_6 = 5'h0 == rob_tail | rob_val_0; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_7 = 5'h1 == rob_tail | rob_val_1; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_8 = 5'h2 == rob_tail | rob_val_2; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_9 = 5'h3 == rob_tail | rob_val_3; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_10 = 5'h4 == rob_tail | rob_val_4; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_11 = 5'h5 == rob_tail | rob_val_5; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_12 = 5'h6 == rob_tail | rob_val_6; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_13 = 5'h7 == rob_tail | rob_val_7; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_14 = 5'h8 == rob_tail | rob_val_8; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_15 = 5'h9 == rob_tail | rob_val_9; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_16 = 5'ha == rob_tail | rob_val_10; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_17 = 5'hb == rob_tail | rob_val_11; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_18 = 5'hc == rob_tail | rob_val_12; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_19 = 5'hd == rob_tail | rob_val_13; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_20 = 5'he == rob_tail | rob_val_14; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_21 = 5'hf == rob_tail | rob_val_15; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_22 = 5'h10 == rob_tail | rob_val_16; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_23 = 5'h11 == rob_tail | rob_val_17; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_24 = 5'h12 == rob_tail | rob_val_18; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_25 = 5'h13 == rob_tail | rob_val_19; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_26 = 5'h14 == rob_tail | rob_val_20; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_27 = 5'h15 == rob_tail | rob_val_21; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_28 = 5'h16 == rob_tail | rob_val_22; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_29 = 5'h17 == rob_tail | rob_val_23; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_30 = 5'h18 == rob_tail | rob_val_24; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_31 = 5'h19 == rob_tail | rob_val_25; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_32 = 5'h1a == rob_tail | rob_val_26; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_33 = 5'h1b == rob_tail | rob_val_27; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_34 = 5'h1c == rob_tail | rob_val_28; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_35 = 5'h1d == rob_tail | rob_val_29; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_36 = 5'h1e == rob_tail | rob_val_30; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_37 = 5'h1f == rob_tail | rob_val_31; // @[rob.scala 324:{31,31} 307:32]
  wire  _GEN_38 = 5'h0 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_0; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_39 = 5'h1 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_1; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_40 = 5'h2 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_2; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_41 = 5'h3 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_3; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_42 = 5'h4 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_4; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_43 = 5'h5 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_5; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_44 = 5'h6 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_6; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_45 = 5'h7 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_7; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_46 = 5'h8 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_8; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_47 = 5'h9 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_9; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_48 = 5'ha == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_10; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_49 = 5'hb == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_11; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_50 = 5'hc == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_12; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_51 = 5'hd == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_13; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_52 = 5'he == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_14; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_53 = 5'hf == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_15; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_54 = 5'h10 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_16; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_55 = 5'h11 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_17; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_56 = 5'h12 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_18; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_57 = 5'h13 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_19; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_58 = 5'h14 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_20; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_59 = 5'h15 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_21; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_60 = 5'h16 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_22; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_61 = 5'h17 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_23; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_62 = 5'h18 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_24; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_63 = 5'h19 == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_25; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_64 = 5'h1a == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_26; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_65 = 5'h1b == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_27; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_66 = 5'h1c == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_28; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_67 = 5'h1d == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_29; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_68 = 5'h1e == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_30; // @[rob.scala 308:28 325:{31,31}]
  wire  _GEN_69 = 5'h1f == rob_tail ? ~(io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei) : rob_bsy_31; // @[rob.scala 308:28 325:{31,31}]
  wire  _T_14 = io_enq_uops_0_uses_ldq | io_enq_uops_0_uses_stq & ~io_enq_uops_0_is_fence | io_enq_uops_0_is_br |
    io_enq_uops_0_is_jalr; // @[micro-op.scala 152:71]
  wire  _GEN_70 = 5'h0 == rob_tail ? _T_14 : rob_unsafe_0; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_71 = 5'h1 == rob_tail ? _T_14 : rob_unsafe_1; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_72 = 5'h2 == rob_tail ? _T_14 : rob_unsafe_2; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_73 = 5'h3 == rob_tail ? _T_14 : rob_unsafe_3; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_74 = 5'h4 == rob_tail ? _T_14 : rob_unsafe_4; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_75 = 5'h5 == rob_tail ? _T_14 : rob_unsafe_5; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_76 = 5'h6 == rob_tail ? _T_14 : rob_unsafe_6; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_77 = 5'h7 == rob_tail ? _T_14 : rob_unsafe_7; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_78 = 5'h8 == rob_tail ? _T_14 : rob_unsafe_8; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_79 = 5'h9 == rob_tail ? _T_14 : rob_unsafe_9; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_80 = 5'ha == rob_tail ? _T_14 : rob_unsafe_10; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_81 = 5'hb == rob_tail ? _T_14 : rob_unsafe_11; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_82 = 5'hc == rob_tail ? _T_14 : rob_unsafe_12; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_83 = 5'hd == rob_tail ? _T_14 : rob_unsafe_13; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_84 = 5'he == rob_tail ? _T_14 : rob_unsafe_14; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_85 = 5'hf == rob_tail ? _T_14 : rob_unsafe_15; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_86 = 5'h10 == rob_tail ? _T_14 : rob_unsafe_16; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_87 = 5'h11 == rob_tail ? _T_14 : rob_unsafe_17; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_88 = 5'h12 == rob_tail ? _T_14 : rob_unsafe_18; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_89 = 5'h13 == rob_tail ? _T_14 : rob_unsafe_19; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_90 = 5'h14 == rob_tail ? _T_14 : rob_unsafe_20; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_91 = 5'h15 == rob_tail ? _T_14 : rob_unsafe_21; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_92 = 5'h16 == rob_tail ? _T_14 : rob_unsafe_22; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_93 = 5'h17 == rob_tail ? _T_14 : rob_unsafe_23; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_94 = 5'h18 == rob_tail ? _T_14 : rob_unsafe_24; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_95 = 5'h19 == rob_tail ? _T_14 : rob_unsafe_25; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_96 = 5'h1a == rob_tail ? _T_14 : rob_unsafe_26; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_97 = 5'h1b == rob_tail ? _T_14 : rob_unsafe_27; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_98 = 5'h1c == rob_tail ? _T_14 : rob_unsafe_28; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_99 = 5'h1d == rob_tail ? _T_14 : rob_unsafe_29; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_100 = 5'h1e == rob_tail ? _T_14 : rob_unsafe_30; // @[rob.scala 309:28 327:{31,31}]
  wire  _GEN_101 = 5'h1f == rob_tail ? _T_14 : rob_unsafe_31; // @[rob.scala 309:28 327:{31,31}]
  wire [1:0] _GEN_134 = 5'h0 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_0_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_135 = 5'h1 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_1_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_136 = 5'h2 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_2_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_137 = 5'h3 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_3_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_138 = 5'h4 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_4_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_139 = 5'h5 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_5_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_140 = 5'h6 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_6_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_141 = 5'h7 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_7_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_142 = 5'h8 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_8_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_143 = 5'h9 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_9_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_144 = 5'ha == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_10_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_145 = 5'hb == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_11_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_146 = 5'hc == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_12_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_147 = 5'hd == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_13_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_148 = 5'he == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_14_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_149 = 5'hf == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_15_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_150 = 5'h10 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_16_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_151 = 5'h11 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_17_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_152 = 5'h12 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_18_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_153 = 5'h13 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_19_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_154 = 5'h14 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_20_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_155 = 5'h15 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_21_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_156 = 5'h16 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_22_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_157 = 5'h17 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_23_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_158 = 5'h18 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_24_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_159 = 5'h19 == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_25_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_160 = 5'h1a == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_26_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_161 = 5'h1b == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_27_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_162 = 5'h1c == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_28_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_163 = 5'h1d == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_29_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_164 = 5'h1e == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_30_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire [1:0] _GEN_165 = 5'h1f == rob_tail ? io_enq_uops_0_debug_fsrc : rob_uop_31_debug_fsrc; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1670 = 5'h0 == rob_tail ? io_enq_uops_0_taken : rob_uop_0_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1671 = 5'h1 == rob_tail ? io_enq_uops_0_taken : rob_uop_1_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1672 = 5'h2 == rob_tail ? io_enq_uops_0_taken : rob_uop_2_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1673 = 5'h3 == rob_tail ? io_enq_uops_0_taken : rob_uop_3_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1674 = 5'h4 == rob_tail ? io_enq_uops_0_taken : rob_uop_4_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1675 = 5'h5 == rob_tail ? io_enq_uops_0_taken : rob_uop_5_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1676 = 5'h6 == rob_tail ? io_enq_uops_0_taken : rob_uop_6_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1677 = 5'h7 == rob_tail ? io_enq_uops_0_taken : rob_uop_7_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1678 = 5'h8 == rob_tail ? io_enq_uops_0_taken : rob_uop_8_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1679 = 5'h9 == rob_tail ? io_enq_uops_0_taken : rob_uop_9_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1680 = 5'ha == rob_tail ? io_enq_uops_0_taken : rob_uop_10_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1681 = 5'hb == rob_tail ? io_enq_uops_0_taken : rob_uop_11_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1682 = 5'hc == rob_tail ? io_enq_uops_0_taken : rob_uop_12_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1683 = 5'hd == rob_tail ? io_enq_uops_0_taken : rob_uop_13_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1684 = 5'he == rob_tail ? io_enq_uops_0_taken : rob_uop_14_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1685 = 5'hf == rob_tail ? io_enq_uops_0_taken : rob_uop_15_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1686 = 5'h10 == rob_tail ? io_enq_uops_0_taken : rob_uop_16_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1687 = 5'h11 == rob_tail ? io_enq_uops_0_taken : rob_uop_17_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1688 = 5'h12 == rob_tail ? io_enq_uops_0_taken : rob_uop_18_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1689 = 5'h13 == rob_tail ? io_enq_uops_0_taken : rob_uop_19_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1690 = 5'h14 == rob_tail ? io_enq_uops_0_taken : rob_uop_20_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1691 = 5'h15 == rob_tail ? io_enq_uops_0_taken : rob_uop_21_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1692 = 5'h16 == rob_tail ? io_enq_uops_0_taken : rob_uop_22_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1693 = 5'h17 == rob_tail ? io_enq_uops_0_taken : rob_uop_23_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1694 = 5'h18 == rob_tail ? io_enq_uops_0_taken : rob_uop_24_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1695 = 5'h19 == rob_tail ? io_enq_uops_0_taken : rob_uop_25_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1696 = 5'h1a == rob_tail ? io_enq_uops_0_taken : rob_uop_26_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1697 = 5'h1b == rob_tail ? io_enq_uops_0_taken : rob_uop_27_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1698 = 5'h1c == rob_tail ? io_enq_uops_0_taken : rob_uop_28_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1699 = 5'h1d == rob_tail ? io_enq_uops_0_taken : rob_uop_29_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1700 = 5'h1e == rob_tail ? io_enq_uops_0_taken : rob_uop_30_taken; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_1701 = 5'h1f == rob_tail ? io_enq_uops_0_taken : rob_uop_31_taken; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1830 = 5'h0 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_0_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1831 = 5'h1 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_1_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1832 = 5'h2 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_2_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1833 = 5'h3 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_3_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1834 = 5'h4 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_4_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1835 = 5'h5 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_5_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1836 = 5'h6 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_6_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1837 = 5'h7 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_7_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1838 = 5'h8 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_8_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1839 = 5'h9 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_9_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1840 = 5'ha == rob_tail ? io_enq_uops_0_br_mask : rob_uop_10_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1841 = 5'hb == rob_tail ? io_enq_uops_0_br_mask : rob_uop_11_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1842 = 5'hc == rob_tail ? io_enq_uops_0_br_mask : rob_uop_12_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1843 = 5'hd == rob_tail ? io_enq_uops_0_br_mask : rob_uop_13_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1844 = 5'he == rob_tail ? io_enq_uops_0_br_mask : rob_uop_14_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1845 = 5'hf == rob_tail ? io_enq_uops_0_br_mask : rob_uop_15_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1846 = 5'h10 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_16_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1847 = 5'h11 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_17_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1848 = 5'h12 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_18_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1849 = 5'h13 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_19_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1850 = 5'h14 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_20_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1851 = 5'h15 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_21_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1852 = 5'h16 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_22_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1853 = 5'h17 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_23_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1854 = 5'h18 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_24_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1855 = 5'h19 == rob_tail ? io_enq_uops_0_br_mask : rob_uop_25_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1856 = 5'h1a == rob_tail ? io_enq_uops_0_br_mask : rob_uop_26_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1857 = 5'h1b == rob_tail ? io_enq_uops_0_br_mask : rob_uop_27_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1858 = 5'h1c == rob_tail ? io_enq_uops_0_br_mask : rob_uop_28_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1859 = 5'h1d == rob_tail ? io_enq_uops_0_br_mask : rob_uop_29_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1860 = 5'h1e == rob_tail ? io_enq_uops_0_br_mask : rob_uop_30_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [7:0] _GEN_1861 = 5'h1f == rob_tail ? io_enq_uops_0_br_mask : rob_uop_31_br_mask; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2534 = 5'h0 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_0_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2535 = 5'h1 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_1_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2536 = 5'h2 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_2_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2537 = 5'h3 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_3_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2538 = 5'h4 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_4_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2539 = 5'h5 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_5_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2540 = 5'h6 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_6_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2541 = 5'h7 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_7_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2542 = 5'h8 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_8_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2543 = 5'h9 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_9_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2544 = 5'ha == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_10_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2545 = 5'hb == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_11_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2546 = 5'hc == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_12_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2547 = 5'hd == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_13_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2548 = 5'he == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_14_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2549 = 5'hf == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_15_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2550 = 5'h10 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_16_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2551 = 5'h11 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_17_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2552 = 5'h12 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_18_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2553 = 5'h13 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_19_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2554 = 5'h14 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_20_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2555 = 5'h15 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_21_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2556 = 5'h16 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_22_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2557 = 5'h17 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_23_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2558 = 5'h18 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_24_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2559 = 5'h19 == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_25_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2560 = 5'h1a == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_26_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2561 = 5'h1b == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_27_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2562 = 5'h1c == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_28_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2563 = 5'h1d == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_29_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2564 = 5'h1e == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_30_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire [31:0] _GEN_2565 = 5'h1f == rob_tail ? io_enq_uops_0_debug_inst : rob_uop_31_debug_inst; // @[rob.scala 310:28 328:{31,31}]
  wire  _GEN_2630 = 5'h0 == rob_tail ? io_enq_uops_0_exception : rob_exception_0; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2631 = 5'h1 == rob_tail ? io_enq_uops_0_exception : rob_exception_1; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2632 = 5'h2 == rob_tail ? io_enq_uops_0_exception : rob_exception_2; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2633 = 5'h3 == rob_tail ? io_enq_uops_0_exception : rob_exception_3; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2634 = 5'h4 == rob_tail ? io_enq_uops_0_exception : rob_exception_4; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2635 = 5'h5 == rob_tail ? io_enq_uops_0_exception : rob_exception_5; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2636 = 5'h6 == rob_tail ? io_enq_uops_0_exception : rob_exception_6; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2637 = 5'h7 == rob_tail ? io_enq_uops_0_exception : rob_exception_7; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2638 = 5'h8 == rob_tail ? io_enq_uops_0_exception : rob_exception_8; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2639 = 5'h9 == rob_tail ? io_enq_uops_0_exception : rob_exception_9; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2640 = 5'ha == rob_tail ? io_enq_uops_0_exception : rob_exception_10; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2641 = 5'hb == rob_tail ? io_enq_uops_0_exception : rob_exception_11; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2642 = 5'hc == rob_tail ? io_enq_uops_0_exception : rob_exception_12; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2643 = 5'hd == rob_tail ? io_enq_uops_0_exception : rob_exception_13; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2644 = 5'he == rob_tail ? io_enq_uops_0_exception : rob_exception_14; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2645 = 5'hf == rob_tail ? io_enq_uops_0_exception : rob_exception_15; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2646 = 5'h10 == rob_tail ? io_enq_uops_0_exception : rob_exception_16; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2647 = 5'h11 == rob_tail ? io_enq_uops_0_exception : rob_exception_17; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2648 = 5'h12 == rob_tail ? io_enq_uops_0_exception : rob_exception_18; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2649 = 5'h13 == rob_tail ? io_enq_uops_0_exception : rob_exception_19; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2650 = 5'h14 == rob_tail ? io_enq_uops_0_exception : rob_exception_20; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2651 = 5'h15 == rob_tail ? io_enq_uops_0_exception : rob_exception_21; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2652 = 5'h16 == rob_tail ? io_enq_uops_0_exception : rob_exception_22; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2653 = 5'h17 == rob_tail ? io_enq_uops_0_exception : rob_exception_23; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2654 = 5'h18 == rob_tail ? io_enq_uops_0_exception : rob_exception_24; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2655 = 5'h19 == rob_tail ? io_enq_uops_0_exception : rob_exception_25; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2656 = 5'h1a == rob_tail ? io_enq_uops_0_exception : rob_exception_26; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2657 = 5'h1b == rob_tail ? io_enq_uops_0_exception : rob_exception_27; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2658 = 5'h1c == rob_tail ? io_enq_uops_0_exception : rob_exception_28; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2659 = 5'h1d == rob_tail ? io_enq_uops_0_exception : rob_exception_29; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2660 = 5'h1e == rob_tail ? io_enq_uops_0_exception : rob_exception_30; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2661 = 5'h1f == rob_tail ? io_enq_uops_0_exception : rob_exception_31; // @[rob.scala 311:28 329:{31,31}]
  wire  _GEN_2662 = 5'h0 == rob_tail ? 1'h0 : rob_predicated_0; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2663 = 5'h1 == rob_tail ? 1'h0 : rob_predicated_1; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2664 = 5'h2 == rob_tail ? 1'h0 : rob_predicated_2; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2665 = 5'h3 == rob_tail ? 1'h0 : rob_predicated_3; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2666 = 5'h4 == rob_tail ? 1'h0 : rob_predicated_4; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2667 = 5'h5 == rob_tail ? 1'h0 : rob_predicated_5; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2668 = 5'h6 == rob_tail ? 1'h0 : rob_predicated_6; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2669 = 5'h7 == rob_tail ? 1'h0 : rob_predicated_7; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2670 = 5'h8 == rob_tail ? 1'h0 : rob_predicated_8; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2671 = 5'h9 == rob_tail ? 1'h0 : rob_predicated_9; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2672 = 5'ha == rob_tail ? 1'h0 : rob_predicated_10; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2673 = 5'hb == rob_tail ? 1'h0 : rob_predicated_11; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2674 = 5'hc == rob_tail ? 1'h0 : rob_predicated_12; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2675 = 5'hd == rob_tail ? 1'h0 : rob_predicated_13; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2676 = 5'he == rob_tail ? 1'h0 : rob_predicated_14; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2677 = 5'hf == rob_tail ? 1'h0 : rob_predicated_15; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2678 = 5'h10 == rob_tail ? 1'h0 : rob_predicated_16; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2679 = 5'h11 == rob_tail ? 1'h0 : rob_predicated_17; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2680 = 5'h12 == rob_tail ? 1'h0 : rob_predicated_18; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2681 = 5'h13 == rob_tail ? 1'h0 : rob_predicated_19; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2682 = 5'h14 == rob_tail ? 1'h0 : rob_predicated_20; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2683 = 5'h15 == rob_tail ? 1'h0 : rob_predicated_21; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2684 = 5'h16 == rob_tail ? 1'h0 : rob_predicated_22; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2685 = 5'h17 == rob_tail ? 1'h0 : rob_predicated_23; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2686 = 5'h18 == rob_tail ? 1'h0 : rob_predicated_24; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2687 = 5'h19 == rob_tail ? 1'h0 : rob_predicated_25; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2688 = 5'h1a == rob_tail ? 1'h0 : rob_predicated_26; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2689 = 5'h1b == rob_tail ? 1'h0 : rob_predicated_27; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2690 = 5'h1c == rob_tail ? 1'h0 : rob_predicated_28; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2691 = 5'h1d == rob_tail ? 1'h0 : rob_predicated_29; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2692 = 5'h1e == rob_tail ? 1'h0 : rob_predicated_30; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2693 = 5'h1f == rob_tail ? 1'h0 : rob_predicated_31; // @[rob.scala 312:29 330:{34,34}]
  wire  _GEN_2695 = 5'h1 == rob_tail ? rob_val_1 : rob_val_0; // @[rob.scala 333:{33,33}]
  wire  _GEN_2696 = 5'h2 == rob_tail ? rob_val_2 : _GEN_2695; // @[rob.scala 333:{33,33}]
  wire  _GEN_2697 = 5'h3 == rob_tail ? rob_val_3 : _GEN_2696; // @[rob.scala 333:{33,33}]
  wire  _GEN_2698 = 5'h4 == rob_tail ? rob_val_4 : _GEN_2697; // @[rob.scala 333:{33,33}]
  wire  _GEN_2699 = 5'h5 == rob_tail ? rob_val_5 : _GEN_2698; // @[rob.scala 333:{33,33}]
  wire  _GEN_2700 = 5'h6 == rob_tail ? rob_val_6 : _GEN_2699; // @[rob.scala 333:{33,33}]
  wire  _GEN_2701 = 5'h7 == rob_tail ? rob_val_7 : _GEN_2700; // @[rob.scala 333:{33,33}]
  wire  _GEN_2702 = 5'h8 == rob_tail ? rob_val_8 : _GEN_2701; // @[rob.scala 333:{33,33}]
  wire  _GEN_2703 = 5'h9 == rob_tail ? rob_val_9 : _GEN_2702; // @[rob.scala 333:{33,33}]
  wire  _GEN_2704 = 5'ha == rob_tail ? rob_val_10 : _GEN_2703; // @[rob.scala 333:{33,33}]
  wire  _GEN_2705 = 5'hb == rob_tail ? rob_val_11 : _GEN_2704; // @[rob.scala 333:{33,33}]
  wire  _GEN_2706 = 5'hc == rob_tail ? rob_val_12 : _GEN_2705; // @[rob.scala 333:{33,33}]
  wire  _GEN_2707 = 5'hd == rob_tail ? rob_val_13 : _GEN_2706; // @[rob.scala 333:{33,33}]
  wire  _GEN_2708 = 5'he == rob_tail ? rob_val_14 : _GEN_2707; // @[rob.scala 333:{33,33}]
  wire  _GEN_2709 = 5'hf == rob_tail ? rob_val_15 : _GEN_2708; // @[rob.scala 333:{33,33}]
  wire  _GEN_2710 = 5'h10 == rob_tail ? rob_val_16 : _GEN_2709; // @[rob.scala 333:{33,33}]
  wire  _GEN_2711 = 5'h11 == rob_tail ? rob_val_17 : _GEN_2710; // @[rob.scala 333:{33,33}]
  wire  _GEN_2712 = 5'h12 == rob_tail ? rob_val_18 : _GEN_2711; // @[rob.scala 333:{33,33}]
  wire  _GEN_2713 = 5'h13 == rob_tail ? rob_val_19 : _GEN_2712; // @[rob.scala 333:{33,33}]
  wire  _GEN_2714 = 5'h14 == rob_tail ? rob_val_20 : _GEN_2713; // @[rob.scala 333:{33,33}]
  wire  _GEN_2715 = 5'h15 == rob_tail ? rob_val_21 : _GEN_2714; // @[rob.scala 333:{33,33}]
  wire  _GEN_2716 = 5'h16 == rob_tail ? rob_val_22 : _GEN_2715; // @[rob.scala 333:{33,33}]
  wire  _GEN_2717 = 5'h17 == rob_tail ? rob_val_23 : _GEN_2716; // @[rob.scala 333:{33,33}]
  wire  _GEN_2718 = 5'h18 == rob_tail ? rob_val_24 : _GEN_2717; // @[rob.scala 333:{33,33}]
  wire  _GEN_2719 = 5'h19 == rob_tail ? rob_val_25 : _GEN_2718; // @[rob.scala 333:{33,33}]
  wire  _GEN_2720 = 5'h1a == rob_tail ? rob_val_26 : _GEN_2719; // @[rob.scala 333:{33,33}]
  wire  _GEN_2721 = 5'h1b == rob_tail ? rob_val_27 : _GEN_2720; // @[rob.scala 333:{33,33}]
  wire  _GEN_2722 = 5'h1c == rob_tail ? rob_val_28 : _GEN_2721; // @[rob.scala 333:{33,33}]
  wire  _GEN_2723 = 5'h1d == rob_tail ? rob_val_29 : _GEN_2722; // @[rob.scala 333:{33,33}]
  wire  _GEN_2724 = 5'h1e == rob_tail ? rob_val_30 : _GEN_2723; // @[rob.scala 333:{33,33}]
  wire  rob_tail_vals_0 = 5'h1f == rob_tail ? rob_val_31 : _GEN_2724; // @[rob.scala 333:{33,33}]
  wire  _T_16 = ~rob_tail_vals_0; // @[rob.scala 333:33]
  wire [31:0] _GEN_2726 = 5'h0 == rob_tail ? 32'h4033 : rob_uop_0_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2727 = 5'h1 == rob_tail ? 32'h4033 : rob_uop_1_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2728 = 5'h2 == rob_tail ? 32'h4033 : rob_uop_2_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2729 = 5'h3 == rob_tail ? 32'h4033 : rob_uop_3_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2730 = 5'h4 == rob_tail ? 32'h4033 : rob_uop_4_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2731 = 5'h5 == rob_tail ? 32'h4033 : rob_uop_5_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2732 = 5'h6 == rob_tail ? 32'h4033 : rob_uop_6_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2733 = 5'h7 == rob_tail ? 32'h4033 : rob_uop_7_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2734 = 5'h8 == rob_tail ? 32'h4033 : rob_uop_8_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2735 = 5'h9 == rob_tail ? 32'h4033 : rob_uop_9_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2736 = 5'ha == rob_tail ? 32'h4033 : rob_uop_10_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2737 = 5'hb == rob_tail ? 32'h4033 : rob_uop_11_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2738 = 5'hc == rob_tail ? 32'h4033 : rob_uop_12_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2739 = 5'hd == rob_tail ? 32'h4033 : rob_uop_13_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2740 = 5'he == rob_tail ? 32'h4033 : rob_uop_14_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2741 = 5'hf == rob_tail ? 32'h4033 : rob_uop_15_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2742 = 5'h10 == rob_tail ? 32'h4033 : rob_uop_16_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2743 = 5'h11 == rob_tail ? 32'h4033 : rob_uop_17_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2744 = 5'h12 == rob_tail ? 32'h4033 : rob_uop_18_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2745 = 5'h13 == rob_tail ? 32'h4033 : rob_uop_19_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2746 = 5'h14 == rob_tail ? 32'h4033 : rob_uop_20_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2747 = 5'h15 == rob_tail ? 32'h4033 : rob_uop_21_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2748 = 5'h16 == rob_tail ? 32'h4033 : rob_uop_22_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2749 = 5'h17 == rob_tail ? 32'h4033 : rob_uop_23_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2750 = 5'h18 == rob_tail ? 32'h4033 : rob_uop_24_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2751 = 5'h19 == rob_tail ? 32'h4033 : rob_uop_25_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2752 = 5'h1a == rob_tail ? 32'h4033 : rob_uop_26_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2753 = 5'h1b == rob_tail ? 32'h4033 : rob_uop_27_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2754 = 5'h1c == rob_tail ? 32'h4033 : rob_uop_28_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2755 = 5'h1d == rob_tail ? 32'h4033 : rob_uop_29_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2756 = 5'h1e == rob_tail ? 32'h4033 : rob_uop_30_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2757 = 5'h1f == rob_tail ? 32'h4033 : rob_uop_31_debug_inst; // @[rob.scala 310:28 336:{36,36}]
  wire [31:0] _GEN_2758 = io_enq_valids_0 & _T_16 ? _GEN_2726 : rob_uop_0_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2759 = io_enq_valids_0 & _T_16 ? _GEN_2727 : rob_uop_1_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2760 = io_enq_valids_0 & _T_16 ? _GEN_2728 : rob_uop_2_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2761 = io_enq_valids_0 & _T_16 ? _GEN_2729 : rob_uop_3_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2762 = io_enq_valids_0 & _T_16 ? _GEN_2730 : rob_uop_4_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2763 = io_enq_valids_0 & _T_16 ? _GEN_2731 : rob_uop_5_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2764 = io_enq_valids_0 & _T_16 ? _GEN_2732 : rob_uop_6_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2765 = io_enq_valids_0 & _T_16 ? _GEN_2733 : rob_uop_7_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2766 = io_enq_valids_0 & _T_16 ? _GEN_2734 : rob_uop_8_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2767 = io_enq_valids_0 & _T_16 ? _GEN_2735 : rob_uop_9_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2768 = io_enq_valids_0 & _T_16 ? _GEN_2736 : rob_uop_10_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2769 = io_enq_valids_0 & _T_16 ? _GEN_2737 : rob_uop_11_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2770 = io_enq_valids_0 & _T_16 ? _GEN_2738 : rob_uop_12_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2771 = io_enq_valids_0 & _T_16 ? _GEN_2739 : rob_uop_13_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2772 = io_enq_valids_0 & _T_16 ? _GEN_2740 : rob_uop_14_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2773 = io_enq_valids_0 & _T_16 ? _GEN_2741 : rob_uop_15_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2774 = io_enq_valids_0 & _T_16 ? _GEN_2742 : rob_uop_16_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2775 = io_enq_valids_0 & _T_16 ? _GEN_2743 : rob_uop_17_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2776 = io_enq_valids_0 & _T_16 ? _GEN_2744 : rob_uop_18_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2777 = io_enq_valids_0 & _T_16 ? _GEN_2745 : rob_uop_19_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2778 = io_enq_valids_0 & _T_16 ? _GEN_2746 : rob_uop_20_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2779 = io_enq_valids_0 & _T_16 ? _GEN_2747 : rob_uop_21_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2780 = io_enq_valids_0 & _T_16 ? _GEN_2748 : rob_uop_22_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2781 = io_enq_valids_0 & _T_16 ? _GEN_2749 : rob_uop_23_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2782 = io_enq_valids_0 & _T_16 ? _GEN_2750 : rob_uop_24_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2783 = io_enq_valids_0 & _T_16 ? _GEN_2751 : rob_uop_25_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2784 = io_enq_valids_0 & _T_16 ? _GEN_2752 : rob_uop_26_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2785 = io_enq_valids_0 & _T_16 ? _GEN_2753 : rob_uop_27_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2786 = io_enq_valids_0 & _T_16 ? _GEN_2754 : rob_uop_28_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2787 = io_enq_valids_0 & _T_16 ? _GEN_2755 : rob_uop_29_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2788 = io_enq_valids_0 & _T_16 ? _GEN_2756 : rob_uop_30_debug_inst; // @[rob.scala 310:28 335:67]
  wire [31:0] _GEN_2789 = io_enq_valids_0 & _T_16 ? _GEN_2757 : rob_uop_31_debug_inst; // @[rob.scala 310:28 335:67]
  wire  _GEN_2790 = io_enq_valids_0 ? _GEN_6 : rob_val_0; // @[rob.scala 323:29 307:32]
  wire  _GEN_2791 = io_enq_valids_0 ? _GEN_7 : rob_val_1; // @[rob.scala 323:29 307:32]
  wire  _GEN_2792 = io_enq_valids_0 ? _GEN_8 : rob_val_2; // @[rob.scala 323:29 307:32]
  wire  _GEN_2793 = io_enq_valids_0 ? _GEN_9 : rob_val_3; // @[rob.scala 323:29 307:32]
  wire  _GEN_2794 = io_enq_valids_0 ? _GEN_10 : rob_val_4; // @[rob.scala 323:29 307:32]
  wire  _GEN_2795 = io_enq_valids_0 ? _GEN_11 : rob_val_5; // @[rob.scala 323:29 307:32]
  wire  _GEN_2796 = io_enq_valids_0 ? _GEN_12 : rob_val_6; // @[rob.scala 323:29 307:32]
  wire  _GEN_2797 = io_enq_valids_0 ? _GEN_13 : rob_val_7; // @[rob.scala 323:29 307:32]
  wire  _GEN_2798 = io_enq_valids_0 ? _GEN_14 : rob_val_8; // @[rob.scala 323:29 307:32]
  wire  _GEN_2799 = io_enq_valids_0 ? _GEN_15 : rob_val_9; // @[rob.scala 323:29 307:32]
  wire  _GEN_2800 = io_enq_valids_0 ? _GEN_16 : rob_val_10; // @[rob.scala 323:29 307:32]
  wire  _GEN_2801 = io_enq_valids_0 ? _GEN_17 : rob_val_11; // @[rob.scala 323:29 307:32]
  wire  _GEN_2802 = io_enq_valids_0 ? _GEN_18 : rob_val_12; // @[rob.scala 323:29 307:32]
  wire  _GEN_2803 = io_enq_valids_0 ? _GEN_19 : rob_val_13; // @[rob.scala 323:29 307:32]
  wire  _GEN_2804 = io_enq_valids_0 ? _GEN_20 : rob_val_14; // @[rob.scala 323:29 307:32]
  wire  _GEN_2805 = io_enq_valids_0 ? _GEN_21 : rob_val_15; // @[rob.scala 323:29 307:32]
  wire  _GEN_2806 = io_enq_valids_0 ? _GEN_22 : rob_val_16; // @[rob.scala 323:29 307:32]
  wire  _GEN_2807 = io_enq_valids_0 ? _GEN_23 : rob_val_17; // @[rob.scala 323:29 307:32]
  wire  _GEN_2808 = io_enq_valids_0 ? _GEN_24 : rob_val_18; // @[rob.scala 323:29 307:32]
  wire  _GEN_2809 = io_enq_valids_0 ? _GEN_25 : rob_val_19; // @[rob.scala 323:29 307:32]
  wire  _GEN_2810 = io_enq_valids_0 ? _GEN_26 : rob_val_20; // @[rob.scala 323:29 307:32]
  wire  _GEN_2811 = io_enq_valids_0 ? _GEN_27 : rob_val_21; // @[rob.scala 323:29 307:32]
  wire  _GEN_2812 = io_enq_valids_0 ? _GEN_28 : rob_val_22; // @[rob.scala 323:29 307:32]
  wire  _GEN_2813 = io_enq_valids_0 ? _GEN_29 : rob_val_23; // @[rob.scala 323:29 307:32]
  wire  _GEN_2814 = io_enq_valids_0 ? _GEN_30 : rob_val_24; // @[rob.scala 323:29 307:32]
  wire  _GEN_2815 = io_enq_valids_0 ? _GEN_31 : rob_val_25; // @[rob.scala 323:29 307:32]
  wire  _GEN_2816 = io_enq_valids_0 ? _GEN_32 : rob_val_26; // @[rob.scala 323:29 307:32]
  wire  _GEN_2817 = io_enq_valids_0 ? _GEN_33 : rob_val_27; // @[rob.scala 323:29 307:32]
  wire  _GEN_2818 = io_enq_valids_0 ? _GEN_34 : rob_val_28; // @[rob.scala 323:29 307:32]
  wire  _GEN_2819 = io_enq_valids_0 ? _GEN_35 : rob_val_29; // @[rob.scala 323:29 307:32]
  wire  _GEN_2820 = io_enq_valids_0 ? _GEN_36 : rob_val_30; // @[rob.scala 323:29 307:32]
  wire  _GEN_2821 = io_enq_valids_0 ? _GEN_37 : rob_val_31; // @[rob.scala 323:29 307:32]
  wire  _GEN_2822 = io_enq_valids_0 ? _GEN_38 : rob_bsy_0; // @[rob.scala 308:28 323:29]
  wire  _GEN_2823 = io_enq_valids_0 ? _GEN_39 : rob_bsy_1; // @[rob.scala 308:28 323:29]
  wire  _GEN_2824 = io_enq_valids_0 ? _GEN_40 : rob_bsy_2; // @[rob.scala 308:28 323:29]
  wire  _GEN_2825 = io_enq_valids_0 ? _GEN_41 : rob_bsy_3; // @[rob.scala 308:28 323:29]
  wire  _GEN_2826 = io_enq_valids_0 ? _GEN_42 : rob_bsy_4; // @[rob.scala 308:28 323:29]
  wire  _GEN_2827 = io_enq_valids_0 ? _GEN_43 : rob_bsy_5; // @[rob.scala 308:28 323:29]
  wire  _GEN_2828 = io_enq_valids_0 ? _GEN_44 : rob_bsy_6; // @[rob.scala 308:28 323:29]
  wire  _GEN_2829 = io_enq_valids_0 ? _GEN_45 : rob_bsy_7; // @[rob.scala 308:28 323:29]
  wire  _GEN_2830 = io_enq_valids_0 ? _GEN_46 : rob_bsy_8; // @[rob.scala 308:28 323:29]
  wire  _GEN_2831 = io_enq_valids_0 ? _GEN_47 : rob_bsy_9; // @[rob.scala 308:28 323:29]
  wire  _GEN_2832 = io_enq_valids_0 ? _GEN_48 : rob_bsy_10; // @[rob.scala 308:28 323:29]
  wire  _GEN_2833 = io_enq_valids_0 ? _GEN_49 : rob_bsy_11; // @[rob.scala 308:28 323:29]
  wire  _GEN_2834 = io_enq_valids_0 ? _GEN_50 : rob_bsy_12; // @[rob.scala 308:28 323:29]
  wire  _GEN_2835 = io_enq_valids_0 ? _GEN_51 : rob_bsy_13; // @[rob.scala 308:28 323:29]
  wire  _GEN_2836 = io_enq_valids_0 ? _GEN_52 : rob_bsy_14; // @[rob.scala 308:28 323:29]
  wire  _GEN_2837 = io_enq_valids_0 ? _GEN_53 : rob_bsy_15; // @[rob.scala 308:28 323:29]
  wire  _GEN_2838 = io_enq_valids_0 ? _GEN_54 : rob_bsy_16; // @[rob.scala 308:28 323:29]
  wire  _GEN_2839 = io_enq_valids_0 ? _GEN_55 : rob_bsy_17; // @[rob.scala 308:28 323:29]
  wire  _GEN_2840 = io_enq_valids_0 ? _GEN_56 : rob_bsy_18; // @[rob.scala 308:28 323:29]
  wire  _GEN_2841 = io_enq_valids_0 ? _GEN_57 : rob_bsy_19; // @[rob.scala 308:28 323:29]
  wire  _GEN_2842 = io_enq_valids_0 ? _GEN_58 : rob_bsy_20; // @[rob.scala 308:28 323:29]
  wire  _GEN_2843 = io_enq_valids_0 ? _GEN_59 : rob_bsy_21; // @[rob.scala 308:28 323:29]
  wire  _GEN_2844 = io_enq_valids_0 ? _GEN_60 : rob_bsy_22; // @[rob.scala 308:28 323:29]
  wire  _GEN_2845 = io_enq_valids_0 ? _GEN_61 : rob_bsy_23; // @[rob.scala 308:28 323:29]
  wire  _GEN_2846 = io_enq_valids_0 ? _GEN_62 : rob_bsy_24; // @[rob.scala 308:28 323:29]
  wire  _GEN_2847 = io_enq_valids_0 ? _GEN_63 : rob_bsy_25; // @[rob.scala 308:28 323:29]
  wire  _GEN_2848 = io_enq_valids_0 ? _GEN_64 : rob_bsy_26; // @[rob.scala 308:28 323:29]
  wire  _GEN_2849 = io_enq_valids_0 ? _GEN_65 : rob_bsy_27; // @[rob.scala 308:28 323:29]
  wire  _GEN_2850 = io_enq_valids_0 ? _GEN_66 : rob_bsy_28; // @[rob.scala 308:28 323:29]
  wire  _GEN_2851 = io_enq_valids_0 ? _GEN_67 : rob_bsy_29; // @[rob.scala 308:28 323:29]
  wire  _GEN_2852 = io_enq_valids_0 ? _GEN_68 : rob_bsy_30; // @[rob.scala 308:28 323:29]
  wire  _GEN_2853 = io_enq_valids_0 ? _GEN_69 : rob_bsy_31; // @[rob.scala 308:28 323:29]
  wire  _GEN_2854 = io_enq_valids_0 ? _GEN_70 : rob_unsafe_0; // @[rob.scala 309:28 323:29]
  wire  _GEN_2855 = io_enq_valids_0 ? _GEN_71 : rob_unsafe_1; // @[rob.scala 309:28 323:29]
  wire  _GEN_2856 = io_enq_valids_0 ? _GEN_72 : rob_unsafe_2; // @[rob.scala 309:28 323:29]
  wire  _GEN_2857 = io_enq_valids_0 ? _GEN_73 : rob_unsafe_3; // @[rob.scala 309:28 323:29]
  wire  _GEN_2858 = io_enq_valids_0 ? _GEN_74 : rob_unsafe_4; // @[rob.scala 309:28 323:29]
  wire  _GEN_2859 = io_enq_valids_0 ? _GEN_75 : rob_unsafe_5; // @[rob.scala 309:28 323:29]
  wire  _GEN_2860 = io_enq_valids_0 ? _GEN_76 : rob_unsafe_6; // @[rob.scala 309:28 323:29]
  wire  _GEN_2861 = io_enq_valids_0 ? _GEN_77 : rob_unsafe_7; // @[rob.scala 309:28 323:29]
  wire  _GEN_2862 = io_enq_valids_0 ? _GEN_78 : rob_unsafe_8; // @[rob.scala 309:28 323:29]
  wire  _GEN_2863 = io_enq_valids_0 ? _GEN_79 : rob_unsafe_9; // @[rob.scala 309:28 323:29]
  wire  _GEN_2864 = io_enq_valids_0 ? _GEN_80 : rob_unsafe_10; // @[rob.scala 309:28 323:29]
  wire  _GEN_2865 = io_enq_valids_0 ? _GEN_81 : rob_unsafe_11; // @[rob.scala 309:28 323:29]
  wire  _GEN_2866 = io_enq_valids_0 ? _GEN_82 : rob_unsafe_12; // @[rob.scala 309:28 323:29]
  wire  _GEN_2867 = io_enq_valids_0 ? _GEN_83 : rob_unsafe_13; // @[rob.scala 309:28 323:29]
  wire  _GEN_2868 = io_enq_valids_0 ? _GEN_84 : rob_unsafe_14; // @[rob.scala 309:28 323:29]
  wire  _GEN_2869 = io_enq_valids_0 ? _GEN_85 : rob_unsafe_15; // @[rob.scala 309:28 323:29]
  wire  _GEN_2870 = io_enq_valids_0 ? _GEN_86 : rob_unsafe_16; // @[rob.scala 309:28 323:29]
  wire  _GEN_2871 = io_enq_valids_0 ? _GEN_87 : rob_unsafe_17; // @[rob.scala 309:28 323:29]
  wire  _GEN_2872 = io_enq_valids_0 ? _GEN_88 : rob_unsafe_18; // @[rob.scala 309:28 323:29]
  wire  _GEN_2873 = io_enq_valids_0 ? _GEN_89 : rob_unsafe_19; // @[rob.scala 309:28 323:29]
  wire  _GEN_2874 = io_enq_valids_0 ? _GEN_90 : rob_unsafe_20; // @[rob.scala 309:28 323:29]
  wire  _GEN_2875 = io_enq_valids_0 ? _GEN_91 : rob_unsafe_21; // @[rob.scala 309:28 323:29]
  wire  _GEN_2876 = io_enq_valids_0 ? _GEN_92 : rob_unsafe_22; // @[rob.scala 309:28 323:29]
  wire  _GEN_2877 = io_enq_valids_0 ? _GEN_93 : rob_unsafe_23; // @[rob.scala 309:28 323:29]
  wire  _GEN_2878 = io_enq_valids_0 ? _GEN_94 : rob_unsafe_24; // @[rob.scala 309:28 323:29]
  wire  _GEN_2879 = io_enq_valids_0 ? _GEN_95 : rob_unsafe_25; // @[rob.scala 309:28 323:29]
  wire  _GEN_2880 = io_enq_valids_0 ? _GEN_96 : rob_unsafe_26; // @[rob.scala 309:28 323:29]
  wire  _GEN_2881 = io_enq_valids_0 ? _GEN_97 : rob_unsafe_27; // @[rob.scala 309:28 323:29]
  wire  _GEN_2882 = io_enq_valids_0 ? _GEN_98 : rob_unsafe_28; // @[rob.scala 309:28 323:29]
  wire  _GEN_2883 = io_enq_valids_0 ? _GEN_99 : rob_unsafe_29; // @[rob.scala 309:28 323:29]
  wire  _GEN_2884 = io_enq_valids_0 ? _GEN_100 : rob_unsafe_30; // @[rob.scala 309:28 323:29]
  wire  _GEN_2885 = io_enq_valids_0 ? _GEN_101 : rob_unsafe_31; // @[rob.scala 309:28 323:29]
  wire [1:0] _GEN_2918 = io_enq_valids_0 ? _GEN_134 : rob_uop_0_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2919 = io_enq_valids_0 ? _GEN_135 : rob_uop_1_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2920 = io_enq_valids_0 ? _GEN_136 : rob_uop_2_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2921 = io_enq_valids_0 ? _GEN_137 : rob_uop_3_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2922 = io_enq_valids_0 ? _GEN_138 : rob_uop_4_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2923 = io_enq_valids_0 ? _GEN_139 : rob_uop_5_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2924 = io_enq_valids_0 ? _GEN_140 : rob_uop_6_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2925 = io_enq_valids_0 ? _GEN_141 : rob_uop_7_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2926 = io_enq_valids_0 ? _GEN_142 : rob_uop_8_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2927 = io_enq_valids_0 ? _GEN_143 : rob_uop_9_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2928 = io_enq_valids_0 ? _GEN_144 : rob_uop_10_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2929 = io_enq_valids_0 ? _GEN_145 : rob_uop_11_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2930 = io_enq_valids_0 ? _GEN_146 : rob_uop_12_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2931 = io_enq_valids_0 ? _GEN_147 : rob_uop_13_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2932 = io_enq_valids_0 ? _GEN_148 : rob_uop_14_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2933 = io_enq_valids_0 ? _GEN_149 : rob_uop_15_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2934 = io_enq_valids_0 ? _GEN_150 : rob_uop_16_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2935 = io_enq_valids_0 ? _GEN_151 : rob_uop_17_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2936 = io_enq_valids_0 ? _GEN_152 : rob_uop_18_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2937 = io_enq_valids_0 ? _GEN_153 : rob_uop_19_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2938 = io_enq_valids_0 ? _GEN_154 : rob_uop_20_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2939 = io_enq_valids_0 ? _GEN_155 : rob_uop_21_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2940 = io_enq_valids_0 ? _GEN_156 : rob_uop_22_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2941 = io_enq_valids_0 ? _GEN_157 : rob_uop_23_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2942 = io_enq_valids_0 ? _GEN_158 : rob_uop_24_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2943 = io_enq_valids_0 ? _GEN_159 : rob_uop_25_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2944 = io_enq_valids_0 ? _GEN_160 : rob_uop_26_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2945 = io_enq_valids_0 ? _GEN_161 : rob_uop_27_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2946 = io_enq_valids_0 ? _GEN_162 : rob_uop_28_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2947 = io_enq_valids_0 ? _GEN_163 : rob_uop_29_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2948 = io_enq_valids_0 ? _GEN_164 : rob_uop_30_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire [1:0] _GEN_2949 = io_enq_valids_0 ? _GEN_165 : rob_uop_31_debug_fsrc; // @[rob.scala 310:28 323:29]
  wire  _GEN_4454 = io_enq_valids_0 ? _GEN_1670 : rob_uop_0_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4455 = io_enq_valids_0 ? _GEN_1671 : rob_uop_1_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4456 = io_enq_valids_0 ? _GEN_1672 : rob_uop_2_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4457 = io_enq_valids_0 ? _GEN_1673 : rob_uop_3_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4458 = io_enq_valids_0 ? _GEN_1674 : rob_uop_4_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4459 = io_enq_valids_0 ? _GEN_1675 : rob_uop_5_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4460 = io_enq_valids_0 ? _GEN_1676 : rob_uop_6_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4461 = io_enq_valids_0 ? _GEN_1677 : rob_uop_7_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4462 = io_enq_valids_0 ? _GEN_1678 : rob_uop_8_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4463 = io_enq_valids_0 ? _GEN_1679 : rob_uop_9_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4464 = io_enq_valids_0 ? _GEN_1680 : rob_uop_10_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4465 = io_enq_valids_0 ? _GEN_1681 : rob_uop_11_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4466 = io_enq_valids_0 ? _GEN_1682 : rob_uop_12_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4467 = io_enq_valids_0 ? _GEN_1683 : rob_uop_13_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4468 = io_enq_valids_0 ? _GEN_1684 : rob_uop_14_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4469 = io_enq_valids_0 ? _GEN_1685 : rob_uop_15_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4470 = io_enq_valids_0 ? _GEN_1686 : rob_uop_16_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4471 = io_enq_valids_0 ? _GEN_1687 : rob_uop_17_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4472 = io_enq_valids_0 ? _GEN_1688 : rob_uop_18_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4473 = io_enq_valids_0 ? _GEN_1689 : rob_uop_19_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4474 = io_enq_valids_0 ? _GEN_1690 : rob_uop_20_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4475 = io_enq_valids_0 ? _GEN_1691 : rob_uop_21_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4476 = io_enq_valids_0 ? _GEN_1692 : rob_uop_22_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4477 = io_enq_valids_0 ? _GEN_1693 : rob_uop_23_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4478 = io_enq_valids_0 ? _GEN_1694 : rob_uop_24_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4479 = io_enq_valids_0 ? _GEN_1695 : rob_uop_25_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4480 = io_enq_valids_0 ? _GEN_1696 : rob_uop_26_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4481 = io_enq_valids_0 ? _GEN_1697 : rob_uop_27_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4482 = io_enq_valids_0 ? _GEN_1698 : rob_uop_28_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4483 = io_enq_valids_0 ? _GEN_1699 : rob_uop_29_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4484 = io_enq_valids_0 ? _GEN_1700 : rob_uop_30_taken; // @[rob.scala 310:28 323:29]
  wire  _GEN_4485 = io_enq_valids_0 ? _GEN_1701 : rob_uop_31_taken; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4614 = io_enq_valids_0 ? _GEN_1830 : rob_uop_0_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4615 = io_enq_valids_0 ? _GEN_1831 : rob_uop_1_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4616 = io_enq_valids_0 ? _GEN_1832 : rob_uop_2_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4617 = io_enq_valids_0 ? _GEN_1833 : rob_uop_3_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4618 = io_enq_valids_0 ? _GEN_1834 : rob_uop_4_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4619 = io_enq_valids_0 ? _GEN_1835 : rob_uop_5_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4620 = io_enq_valids_0 ? _GEN_1836 : rob_uop_6_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4621 = io_enq_valids_0 ? _GEN_1837 : rob_uop_7_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4622 = io_enq_valids_0 ? _GEN_1838 : rob_uop_8_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4623 = io_enq_valids_0 ? _GEN_1839 : rob_uop_9_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4624 = io_enq_valids_0 ? _GEN_1840 : rob_uop_10_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4625 = io_enq_valids_0 ? _GEN_1841 : rob_uop_11_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4626 = io_enq_valids_0 ? _GEN_1842 : rob_uop_12_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4627 = io_enq_valids_0 ? _GEN_1843 : rob_uop_13_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4628 = io_enq_valids_0 ? _GEN_1844 : rob_uop_14_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4629 = io_enq_valids_0 ? _GEN_1845 : rob_uop_15_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4630 = io_enq_valids_0 ? _GEN_1846 : rob_uop_16_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4631 = io_enq_valids_0 ? _GEN_1847 : rob_uop_17_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4632 = io_enq_valids_0 ? _GEN_1848 : rob_uop_18_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4633 = io_enq_valids_0 ? _GEN_1849 : rob_uop_19_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4634 = io_enq_valids_0 ? _GEN_1850 : rob_uop_20_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4635 = io_enq_valids_0 ? _GEN_1851 : rob_uop_21_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4636 = io_enq_valids_0 ? _GEN_1852 : rob_uop_22_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4637 = io_enq_valids_0 ? _GEN_1853 : rob_uop_23_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4638 = io_enq_valids_0 ? _GEN_1854 : rob_uop_24_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4639 = io_enq_valids_0 ? _GEN_1855 : rob_uop_25_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4640 = io_enq_valids_0 ? _GEN_1856 : rob_uop_26_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4641 = io_enq_valids_0 ? _GEN_1857 : rob_uop_27_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4642 = io_enq_valids_0 ? _GEN_1858 : rob_uop_28_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4643 = io_enq_valids_0 ? _GEN_1859 : rob_uop_29_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4644 = io_enq_valids_0 ? _GEN_1860 : rob_uop_30_br_mask; // @[rob.scala 310:28 323:29]
  wire [7:0] _GEN_4645 = io_enq_valids_0 ? _GEN_1861 : rob_uop_31_br_mask; // @[rob.scala 310:28 323:29]
  wire [31:0] _GEN_5318 = io_enq_valids_0 ? _GEN_2534 : _GEN_2758; // @[rob.scala 323:29]
  wire [31:0] _GEN_5319 = io_enq_valids_0 ? _GEN_2535 : _GEN_2759; // @[rob.scala 323:29]
  wire [31:0] _GEN_5320 = io_enq_valids_0 ? _GEN_2536 : _GEN_2760; // @[rob.scala 323:29]
  wire [31:0] _GEN_5321 = io_enq_valids_0 ? _GEN_2537 : _GEN_2761; // @[rob.scala 323:29]
  wire [31:0] _GEN_5322 = io_enq_valids_0 ? _GEN_2538 : _GEN_2762; // @[rob.scala 323:29]
  wire [31:0] _GEN_5323 = io_enq_valids_0 ? _GEN_2539 : _GEN_2763; // @[rob.scala 323:29]
  wire [31:0] _GEN_5324 = io_enq_valids_0 ? _GEN_2540 : _GEN_2764; // @[rob.scala 323:29]
  wire [31:0] _GEN_5325 = io_enq_valids_0 ? _GEN_2541 : _GEN_2765; // @[rob.scala 323:29]
  wire [31:0] _GEN_5326 = io_enq_valids_0 ? _GEN_2542 : _GEN_2766; // @[rob.scala 323:29]
  wire [31:0] _GEN_5327 = io_enq_valids_0 ? _GEN_2543 : _GEN_2767; // @[rob.scala 323:29]
  wire [31:0] _GEN_5328 = io_enq_valids_0 ? _GEN_2544 : _GEN_2768; // @[rob.scala 323:29]
  wire [31:0] _GEN_5329 = io_enq_valids_0 ? _GEN_2545 : _GEN_2769; // @[rob.scala 323:29]
  wire [31:0] _GEN_5330 = io_enq_valids_0 ? _GEN_2546 : _GEN_2770; // @[rob.scala 323:29]
  wire [31:0] _GEN_5331 = io_enq_valids_0 ? _GEN_2547 : _GEN_2771; // @[rob.scala 323:29]
  wire [31:0] _GEN_5332 = io_enq_valids_0 ? _GEN_2548 : _GEN_2772; // @[rob.scala 323:29]
  wire [31:0] _GEN_5333 = io_enq_valids_0 ? _GEN_2549 : _GEN_2773; // @[rob.scala 323:29]
  wire [31:0] _GEN_5334 = io_enq_valids_0 ? _GEN_2550 : _GEN_2774; // @[rob.scala 323:29]
  wire [31:0] _GEN_5335 = io_enq_valids_0 ? _GEN_2551 : _GEN_2775; // @[rob.scala 323:29]
  wire [31:0] _GEN_5336 = io_enq_valids_0 ? _GEN_2552 : _GEN_2776; // @[rob.scala 323:29]
  wire [31:0] _GEN_5337 = io_enq_valids_0 ? _GEN_2553 : _GEN_2777; // @[rob.scala 323:29]
  wire [31:0] _GEN_5338 = io_enq_valids_0 ? _GEN_2554 : _GEN_2778; // @[rob.scala 323:29]
  wire [31:0] _GEN_5339 = io_enq_valids_0 ? _GEN_2555 : _GEN_2779; // @[rob.scala 323:29]
  wire [31:0] _GEN_5340 = io_enq_valids_0 ? _GEN_2556 : _GEN_2780; // @[rob.scala 323:29]
  wire [31:0] _GEN_5341 = io_enq_valids_0 ? _GEN_2557 : _GEN_2781; // @[rob.scala 323:29]
  wire [31:0] _GEN_5342 = io_enq_valids_0 ? _GEN_2558 : _GEN_2782; // @[rob.scala 323:29]
  wire [31:0] _GEN_5343 = io_enq_valids_0 ? _GEN_2559 : _GEN_2783; // @[rob.scala 323:29]
  wire [31:0] _GEN_5344 = io_enq_valids_0 ? _GEN_2560 : _GEN_2784; // @[rob.scala 323:29]
  wire [31:0] _GEN_5345 = io_enq_valids_0 ? _GEN_2561 : _GEN_2785; // @[rob.scala 323:29]
  wire [31:0] _GEN_5346 = io_enq_valids_0 ? _GEN_2562 : _GEN_2786; // @[rob.scala 323:29]
  wire [31:0] _GEN_5347 = io_enq_valids_0 ? _GEN_2563 : _GEN_2787; // @[rob.scala 323:29]
  wire [31:0] _GEN_5348 = io_enq_valids_0 ? _GEN_2564 : _GEN_2788; // @[rob.scala 323:29]
  wire [31:0] _GEN_5349 = io_enq_valids_0 ? _GEN_2565 : _GEN_2789; // @[rob.scala 323:29]
  wire  _GEN_5414 = io_enq_valids_0 ? _GEN_2630 : rob_exception_0; // @[rob.scala 311:28 323:29]
  wire  _GEN_5415 = io_enq_valids_0 ? _GEN_2631 : rob_exception_1; // @[rob.scala 311:28 323:29]
  wire  _GEN_5416 = io_enq_valids_0 ? _GEN_2632 : rob_exception_2; // @[rob.scala 311:28 323:29]
  wire  _GEN_5417 = io_enq_valids_0 ? _GEN_2633 : rob_exception_3; // @[rob.scala 311:28 323:29]
  wire  _GEN_5418 = io_enq_valids_0 ? _GEN_2634 : rob_exception_4; // @[rob.scala 311:28 323:29]
  wire  _GEN_5419 = io_enq_valids_0 ? _GEN_2635 : rob_exception_5; // @[rob.scala 311:28 323:29]
  wire  _GEN_5420 = io_enq_valids_0 ? _GEN_2636 : rob_exception_6; // @[rob.scala 311:28 323:29]
  wire  _GEN_5421 = io_enq_valids_0 ? _GEN_2637 : rob_exception_7; // @[rob.scala 311:28 323:29]
  wire  _GEN_5422 = io_enq_valids_0 ? _GEN_2638 : rob_exception_8; // @[rob.scala 311:28 323:29]
  wire  _GEN_5423 = io_enq_valids_0 ? _GEN_2639 : rob_exception_9; // @[rob.scala 311:28 323:29]
  wire  _GEN_5424 = io_enq_valids_0 ? _GEN_2640 : rob_exception_10; // @[rob.scala 311:28 323:29]
  wire  _GEN_5425 = io_enq_valids_0 ? _GEN_2641 : rob_exception_11; // @[rob.scala 311:28 323:29]
  wire  _GEN_5426 = io_enq_valids_0 ? _GEN_2642 : rob_exception_12; // @[rob.scala 311:28 323:29]
  wire  _GEN_5427 = io_enq_valids_0 ? _GEN_2643 : rob_exception_13; // @[rob.scala 311:28 323:29]
  wire  _GEN_5428 = io_enq_valids_0 ? _GEN_2644 : rob_exception_14; // @[rob.scala 311:28 323:29]
  wire  _GEN_5429 = io_enq_valids_0 ? _GEN_2645 : rob_exception_15; // @[rob.scala 311:28 323:29]
  wire  _GEN_5430 = io_enq_valids_0 ? _GEN_2646 : rob_exception_16; // @[rob.scala 311:28 323:29]
  wire  _GEN_5431 = io_enq_valids_0 ? _GEN_2647 : rob_exception_17; // @[rob.scala 311:28 323:29]
  wire  _GEN_5432 = io_enq_valids_0 ? _GEN_2648 : rob_exception_18; // @[rob.scala 311:28 323:29]
  wire  _GEN_5433 = io_enq_valids_0 ? _GEN_2649 : rob_exception_19; // @[rob.scala 311:28 323:29]
  wire  _GEN_5434 = io_enq_valids_0 ? _GEN_2650 : rob_exception_20; // @[rob.scala 311:28 323:29]
  wire  _GEN_5435 = io_enq_valids_0 ? _GEN_2651 : rob_exception_21; // @[rob.scala 311:28 323:29]
  wire  _GEN_5436 = io_enq_valids_0 ? _GEN_2652 : rob_exception_22; // @[rob.scala 311:28 323:29]
  wire  _GEN_5437 = io_enq_valids_0 ? _GEN_2653 : rob_exception_23; // @[rob.scala 311:28 323:29]
  wire  _GEN_5438 = io_enq_valids_0 ? _GEN_2654 : rob_exception_24; // @[rob.scala 311:28 323:29]
  wire  _GEN_5439 = io_enq_valids_0 ? _GEN_2655 : rob_exception_25; // @[rob.scala 311:28 323:29]
  wire  _GEN_5440 = io_enq_valids_0 ? _GEN_2656 : rob_exception_26; // @[rob.scala 311:28 323:29]
  wire  _GEN_5441 = io_enq_valids_0 ? _GEN_2657 : rob_exception_27; // @[rob.scala 311:28 323:29]
  wire  _GEN_5442 = io_enq_valids_0 ? _GEN_2658 : rob_exception_28; // @[rob.scala 311:28 323:29]
  wire  _GEN_5443 = io_enq_valids_0 ? _GEN_2659 : rob_exception_29; // @[rob.scala 311:28 323:29]
  wire  _GEN_5444 = io_enq_valids_0 ? _GEN_2660 : rob_exception_30; // @[rob.scala 311:28 323:29]
  wire  _GEN_5445 = io_enq_valids_0 ? _GEN_2661 : rob_exception_31; // @[rob.scala 311:28 323:29]
  wire  _GEN_5446 = io_enq_valids_0 ? _GEN_2662 : rob_predicated_0; // @[rob.scala 312:29 323:29]
  wire  _GEN_5447 = io_enq_valids_0 ? _GEN_2663 : rob_predicated_1; // @[rob.scala 312:29 323:29]
  wire  _GEN_5448 = io_enq_valids_0 ? _GEN_2664 : rob_predicated_2; // @[rob.scala 312:29 323:29]
  wire  _GEN_5449 = io_enq_valids_0 ? _GEN_2665 : rob_predicated_3; // @[rob.scala 312:29 323:29]
  wire  _GEN_5450 = io_enq_valids_0 ? _GEN_2666 : rob_predicated_4; // @[rob.scala 312:29 323:29]
  wire  _GEN_5451 = io_enq_valids_0 ? _GEN_2667 : rob_predicated_5; // @[rob.scala 312:29 323:29]
  wire  _GEN_5452 = io_enq_valids_0 ? _GEN_2668 : rob_predicated_6; // @[rob.scala 312:29 323:29]
  wire  _GEN_5453 = io_enq_valids_0 ? _GEN_2669 : rob_predicated_7; // @[rob.scala 312:29 323:29]
  wire  _GEN_5454 = io_enq_valids_0 ? _GEN_2670 : rob_predicated_8; // @[rob.scala 312:29 323:29]
  wire  _GEN_5455 = io_enq_valids_0 ? _GEN_2671 : rob_predicated_9; // @[rob.scala 312:29 323:29]
  wire  _GEN_5456 = io_enq_valids_0 ? _GEN_2672 : rob_predicated_10; // @[rob.scala 312:29 323:29]
  wire  _GEN_5457 = io_enq_valids_0 ? _GEN_2673 : rob_predicated_11; // @[rob.scala 312:29 323:29]
  wire  _GEN_5458 = io_enq_valids_0 ? _GEN_2674 : rob_predicated_12; // @[rob.scala 312:29 323:29]
  wire  _GEN_5459 = io_enq_valids_0 ? _GEN_2675 : rob_predicated_13; // @[rob.scala 312:29 323:29]
  wire  _GEN_5460 = io_enq_valids_0 ? _GEN_2676 : rob_predicated_14; // @[rob.scala 312:29 323:29]
  wire  _GEN_5461 = io_enq_valids_0 ? _GEN_2677 : rob_predicated_15; // @[rob.scala 312:29 323:29]
  wire  _GEN_5462 = io_enq_valids_0 ? _GEN_2678 : rob_predicated_16; // @[rob.scala 312:29 323:29]
  wire  _GEN_5463 = io_enq_valids_0 ? _GEN_2679 : rob_predicated_17; // @[rob.scala 312:29 323:29]
  wire  _GEN_5464 = io_enq_valids_0 ? _GEN_2680 : rob_predicated_18; // @[rob.scala 312:29 323:29]
  wire  _GEN_5465 = io_enq_valids_0 ? _GEN_2681 : rob_predicated_19; // @[rob.scala 312:29 323:29]
  wire  _GEN_5466 = io_enq_valids_0 ? _GEN_2682 : rob_predicated_20; // @[rob.scala 312:29 323:29]
  wire  _GEN_5467 = io_enq_valids_0 ? _GEN_2683 : rob_predicated_21; // @[rob.scala 312:29 323:29]
  wire  _GEN_5468 = io_enq_valids_0 ? _GEN_2684 : rob_predicated_22; // @[rob.scala 312:29 323:29]
  wire  _GEN_5469 = io_enq_valids_0 ? _GEN_2685 : rob_predicated_23; // @[rob.scala 312:29 323:29]
  wire  _GEN_5470 = io_enq_valids_0 ? _GEN_2686 : rob_predicated_24; // @[rob.scala 312:29 323:29]
  wire  _GEN_5471 = io_enq_valids_0 ? _GEN_2687 : rob_predicated_25; // @[rob.scala 312:29 323:29]
  wire  _GEN_5472 = io_enq_valids_0 ? _GEN_2688 : rob_predicated_26; // @[rob.scala 312:29 323:29]
  wire  _GEN_5473 = io_enq_valids_0 ? _GEN_2689 : rob_predicated_27; // @[rob.scala 312:29 323:29]
  wire  _GEN_5474 = io_enq_valids_0 ? _GEN_2690 : rob_predicated_28; // @[rob.scala 312:29 323:29]
  wire  _GEN_5475 = io_enq_valids_0 ? _GEN_2691 : rob_predicated_29; // @[rob.scala 312:29 323:29]
  wire  _GEN_5476 = io_enq_valids_0 ? _GEN_2692 : rob_predicated_30; // @[rob.scala 312:29 323:29]
  wire  _GEN_5477 = io_enq_valids_0 ? _GEN_2693 : rob_predicated_31; // @[rob.scala 312:29 323:29]
  wire  _GEN_5483 = 5'h0 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2822; // @[rob.scala 347:{31,31}]
  wire  _GEN_5484 = 5'h1 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2823; // @[rob.scala 347:{31,31}]
  wire  _GEN_5485 = 5'h2 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2824; // @[rob.scala 347:{31,31}]
  wire  _GEN_5486 = 5'h3 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2825; // @[rob.scala 347:{31,31}]
  wire  _GEN_5487 = 5'h4 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2826; // @[rob.scala 347:{31,31}]
  wire  _GEN_5488 = 5'h5 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2827; // @[rob.scala 347:{31,31}]
  wire  _GEN_5489 = 5'h6 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2828; // @[rob.scala 347:{31,31}]
  wire  _GEN_5490 = 5'h7 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2829; // @[rob.scala 347:{31,31}]
  wire  _GEN_5491 = 5'h8 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2830; // @[rob.scala 347:{31,31}]
  wire  _GEN_5492 = 5'h9 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2831; // @[rob.scala 347:{31,31}]
  wire  _GEN_5493 = 5'ha == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2832; // @[rob.scala 347:{31,31}]
  wire  _GEN_5494 = 5'hb == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2833; // @[rob.scala 347:{31,31}]
  wire  _GEN_5495 = 5'hc == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2834; // @[rob.scala 347:{31,31}]
  wire  _GEN_5496 = 5'hd == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2835; // @[rob.scala 347:{31,31}]
  wire  _GEN_5497 = 5'he == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2836; // @[rob.scala 347:{31,31}]
  wire  _GEN_5498 = 5'hf == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2837; // @[rob.scala 347:{31,31}]
  wire  _GEN_5499 = 5'h10 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2838; // @[rob.scala 347:{31,31}]
  wire  _GEN_5500 = 5'h11 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2839; // @[rob.scala 347:{31,31}]
  wire  _GEN_5501 = 5'h12 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2840; // @[rob.scala 347:{31,31}]
  wire  _GEN_5502 = 5'h13 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2841; // @[rob.scala 347:{31,31}]
  wire  _GEN_5503 = 5'h14 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2842; // @[rob.scala 347:{31,31}]
  wire  _GEN_5504 = 5'h15 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2843; // @[rob.scala 347:{31,31}]
  wire  _GEN_5505 = 5'h16 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2844; // @[rob.scala 347:{31,31}]
  wire  _GEN_5506 = 5'h17 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2845; // @[rob.scala 347:{31,31}]
  wire  _GEN_5507 = 5'h18 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2846; // @[rob.scala 347:{31,31}]
  wire  _GEN_5508 = 5'h19 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2847; // @[rob.scala 347:{31,31}]
  wire  _GEN_5509 = 5'h1a == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2848; // @[rob.scala 347:{31,31}]
  wire  _GEN_5510 = 5'h1b == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2849; // @[rob.scala 347:{31,31}]
  wire  _GEN_5511 = 5'h1c == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2850; // @[rob.scala 347:{31,31}]
  wire  _GEN_5512 = 5'h1d == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2851; // @[rob.scala 347:{31,31}]
  wire  _GEN_5513 = 5'h1e == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2852; // @[rob.scala 347:{31,31}]
  wire  _GEN_5514 = 5'h1f == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2853; // @[rob.scala 347:{31,31}]
  wire  _GEN_5515 = 5'h0 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2854; // @[rob.scala 348:{31,31}]
  wire  _GEN_5516 = 5'h1 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2855; // @[rob.scala 348:{31,31}]
  wire  _GEN_5517 = 5'h2 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2856; // @[rob.scala 348:{31,31}]
  wire  _GEN_5518 = 5'h3 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2857; // @[rob.scala 348:{31,31}]
  wire  _GEN_5519 = 5'h4 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2858; // @[rob.scala 348:{31,31}]
  wire  _GEN_5520 = 5'h5 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2859; // @[rob.scala 348:{31,31}]
  wire  _GEN_5521 = 5'h6 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2860; // @[rob.scala 348:{31,31}]
  wire  _GEN_5522 = 5'h7 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2861; // @[rob.scala 348:{31,31}]
  wire  _GEN_5523 = 5'h8 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2862; // @[rob.scala 348:{31,31}]
  wire  _GEN_5524 = 5'h9 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2863; // @[rob.scala 348:{31,31}]
  wire  _GEN_5525 = 5'ha == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2864; // @[rob.scala 348:{31,31}]
  wire  _GEN_5526 = 5'hb == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2865; // @[rob.scala 348:{31,31}]
  wire  _GEN_5527 = 5'hc == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2866; // @[rob.scala 348:{31,31}]
  wire  _GEN_5528 = 5'hd == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2867; // @[rob.scala 348:{31,31}]
  wire  _GEN_5529 = 5'he == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2868; // @[rob.scala 348:{31,31}]
  wire  _GEN_5530 = 5'hf == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2869; // @[rob.scala 348:{31,31}]
  wire  _GEN_5531 = 5'h10 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2870; // @[rob.scala 348:{31,31}]
  wire  _GEN_5532 = 5'h11 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2871; // @[rob.scala 348:{31,31}]
  wire  _GEN_5533 = 5'h12 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2872; // @[rob.scala 348:{31,31}]
  wire  _GEN_5534 = 5'h13 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2873; // @[rob.scala 348:{31,31}]
  wire  _GEN_5535 = 5'h14 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2874; // @[rob.scala 348:{31,31}]
  wire  _GEN_5536 = 5'h15 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2875; // @[rob.scala 348:{31,31}]
  wire  _GEN_5537 = 5'h16 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2876; // @[rob.scala 348:{31,31}]
  wire  _GEN_5538 = 5'h17 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2877; // @[rob.scala 348:{31,31}]
  wire  _GEN_5539 = 5'h18 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2878; // @[rob.scala 348:{31,31}]
  wire  _GEN_5540 = 5'h19 == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2879; // @[rob.scala 348:{31,31}]
  wire  _GEN_5541 = 5'h1a == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2880; // @[rob.scala 348:{31,31}]
  wire  _GEN_5542 = 5'h1b == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2881; // @[rob.scala 348:{31,31}]
  wire  _GEN_5543 = 5'h1c == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2882; // @[rob.scala 348:{31,31}]
  wire  _GEN_5544 = 5'h1d == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2883; // @[rob.scala 348:{31,31}]
  wire  _GEN_5545 = 5'h1e == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2884; // @[rob.scala 348:{31,31}]
  wire  _GEN_5546 = 5'h1f == io_wb_resps_0_bits_uop_rob_idx ? 1'h0 : _GEN_2885; // @[rob.scala 348:{31,31}]
  wire  _GEN_5547 = 5'h0 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5446; // @[rob.scala 349:{34,34}]
  wire  _GEN_5548 = 5'h1 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5447; // @[rob.scala 349:{34,34}]
  wire  _GEN_5549 = 5'h2 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5448; // @[rob.scala 349:{34,34}]
  wire  _GEN_5550 = 5'h3 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5449; // @[rob.scala 349:{34,34}]
  wire  _GEN_5551 = 5'h4 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5450; // @[rob.scala 349:{34,34}]
  wire  _GEN_5552 = 5'h5 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5451; // @[rob.scala 349:{34,34}]
  wire  _GEN_5553 = 5'h6 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5452; // @[rob.scala 349:{34,34}]
  wire  _GEN_5554 = 5'h7 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5453; // @[rob.scala 349:{34,34}]
  wire  _GEN_5555 = 5'h8 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5454; // @[rob.scala 349:{34,34}]
  wire  _GEN_5556 = 5'h9 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5455; // @[rob.scala 349:{34,34}]
  wire  _GEN_5557 = 5'ha == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5456; // @[rob.scala 349:{34,34}]
  wire  _GEN_5558 = 5'hb == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5457; // @[rob.scala 349:{34,34}]
  wire  _GEN_5559 = 5'hc == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5458; // @[rob.scala 349:{34,34}]
  wire  _GEN_5560 = 5'hd == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5459; // @[rob.scala 349:{34,34}]
  wire  _GEN_5561 = 5'he == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5460; // @[rob.scala 349:{34,34}]
  wire  _GEN_5562 = 5'hf == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5461; // @[rob.scala 349:{34,34}]
  wire  _GEN_5563 = 5'h10 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5462; // @[rob.scala 349:{34,34}]
  wire  _GEN_5564 = 5'h11 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5463; // @[rob.scala 349:{34,34}]
  wire  _GEN_5565 = 5'h12 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5464; // @[rob.scala 349:{34,34}]
  wire  _GEN_5566 = 5'h13 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5465; // @[rob.scala 349:{34,34}]
  wire  _GEN_5567 = 5'h14 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5466; // @[rob.scala 349:{34,34}]
  wire  _GEN_5568 = 5'h15 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5467; // @[rob.scala 349:{34,34}]
  wire  _GEN_5569 = 5'h16 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5468; // @[rob.scala 349:{34,34}]
  wire  _GEN_5570 = 5'h17 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5469; // @[rob.scala 349:{34,34}]
  wire  _GEN_5571 = 5'h18 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5470; // @[rob.scala 349:{34,34}]
  wire  _GEN_5572 = 5'h19 == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5471; // @[rob.scala 349:{34,34}]
  wire  _GEN_5573 = 5'h1a == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5472; // @[rob.scala 349:{34,34}]
  wire  _GEN_5574 = 5'h1b == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5473; // @[rob.scala 349:{34,34}]
  wire  _GEN_5575 = 5'h1c == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5474; // @[rob.scala 349:{34,34}]
  wire  _GEN_5576 = 5'h1d == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5475; // @[rob.scala 349:{34,34}]
  wire  _GEN_5577 = 5'h1e == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5476; // @[rob.scala 349:{34,34}]
  wire  _GEN_5578 = 5'h1f == io_wb_resps_0_bits_uop_rob_idx ? io_wb_resps_0_bits_predicated : _GEN_5477; // @[rob.scala 349:{34,34}]
  wire  _GEN_5579 = io_wb_resps_0_valid ? _GEN_5483 : _GEN_2822; // @[rob.scala 346:69]
  wire  _GEN_5580 = io_wb_resps_0_valid ? _GEN_5484 : _GEN_2823; // @[rob.scala 346:69]
  wire  _GEN_5581 = io_wb_resps_0_valid ? _GEN_5485 : _GEN_2824; // @[rob.scala 346:69]
  wire  _GEN_5582 = io_wb_resps_0_valid ? _GEN_5486 : _GEN_2825; // @[rob.scala 346:69]
  wire  _GEN_5583 = io_wb_resps_0_valid ? _GEN_5487 : _GEN_2826; // @[rob.scala 346:69]
  wire  _GEN_5584 = io_wb_resps_0_valid ? _GEN_5488 : _GEN_2827; // @[rob.scala 346:69]
  wire  _GEN_5585 = io_wb_resps_0_valid ? _GEN_5489 : _GEN_2828; // @[rob.scala 346:69]
  wire  _GEN_5586 = io_wb_resps_0_valid ? _GEN_5490 : _GEN_2829; // @[rob.scala 346:69]
  wire  _GEN_5587 = io_wb_resps_0_valid ? _GEN_5491 : _GEN_2830; // @[rob.scala 346:69]
  wire  _GEN_5588 = io_wb_resps_0_valid ? _GEN_5492 : _GEN_2831; // @[rob.scala 346:69]
  wire  _GEN_5589 = io_wb_resps_0_valid ? _GEN_5493 : _GEN_2832; // @[rob.scala 346:69]
  wire  _GEN_5590 = io_wb_resps_0_valid ? _GEN_5494 : _GEN_2833; // @[rob.scala 346:69]
  wire  _GEN_5591 = io_wb_resps_0_valid ? _GEN_5495 : _GEN_2834; // @[rob.scala 346:69]
  wire  _GEN_5592 = io_wb_resps_0_valid ? _GEN_5496 : _GEN_2835; // @[rob.scala 346:69]
  wire  _GEN_5593 = io_wb_resps_0_valid ? _GEN_5497 : _GEN_2836; // @[rob.scala 346:69]
  wire  _GEN_5594 = io_wb_resps_0_valid ? _GEN_5498 : _GEN_2837; // @[rob.scala 346:69]
  wire  _GEN_5595 = io_wb_resps_0_valid ? _GEN_5499 : _GEN_2838; // @[rob.scala 346:69]
  wire  _GEN_5596 = io_wb_resps_0_valid ? _GEN_5500 : _GEN_2839; // @[rob.scala 346:69]
  wire  _GEN_5597 = io_wb_resps_0_valid ? _GEN_5501 : _GEN_2840; // @[rob.scala 346:69]
  wire  _GEN_5598 = io_wb_resps_0_valid ? _GEN_5502 : _GEN_2841; // @[rob.scala 346:69]
  wire  _GEN_5599 = io_wb_resps_0_valid ? _GEN_5503 : _GEN_2842; // @[rob.scala 346:69]
  wire  _GEN_5600 = io_wb_resps_0_valid ? _GEN_5504 : _GEN_2843; // @[rob.scala 346:69]
  wire  _GEN_5601 = io_wb_resps_0_valid ? _GEN_5505 : _GEN_2844; // @[rob.scala 346:69]
  wire  _GEN_5602 = io_wb_resps_0_valid ? _GEN_5506 : _GEN_2845; // @[rob.scala 346:69]
  wire  _GEN_5603 = io_wb_resps_0_valid ? _GEN_5507 : _GEN_2846; // @[rob.scala 346:69]
  wire  _GEN_5604 = io_wb_resps_0_valid ? _GEN_5508 : _GEN_2847; // @[rob.scala 346:69]
  wire  _GEN_5605 = io_wb_resps_0_valid ? _GEN_5509 : _GEN_2848; // @[rob.scala 346:69]
  wire  _GEN_5606 = io_wb_resps_0_valid ? _GEN_5510 : _GEN_2849; // @[rob.scala 346:69]
  wire  _GEN_5607 = io_wb_resps_0_valid ? _GEN_5511 : _GEN_2850; // @[rob.scala 346:69]
  wire  _GEN_5608 = io_wb_resps_0_valid ? _GEN_5512 : _GEN_2851; // @[rob.scala 346:69]
  wire  _GEN_5609 = io_wb_resps_0_valid ? _GEN_5513 : _GEN_2852; // @[rob.scala 346:69]
  wire  _GEN_5610 = io_wb_resps_0_valid ? _GEN_5514 : _GEN_2853; // @[rob.scala 346:69]
  wire  _GEN_5611 = io_wb_resps_0_valid ? _GEN_5515 : _GEN_2854; // @[rob.scala 346:69]
  wire  _GEN_5612 = io_wb_resps_0_valid ? _GEN_5516 : _GEN_2855; // @[rob.scala 346:69]
  wire  _GEN_5613 = io_wb_resps_0_valid ? _GEN_5517 : _GEN_2856; // @[rob.scala 346:69]
  wire  _GEN_5614 = io_wb_resps_0_valid ? _GEN_5518 : _GEN_2857; // @[rob.scala 346:69]
  wire  _GEN_5615 = io_wb_resps_0_valid ? _GEN_5519 : _GEN_2858; // @[rob.scala 346:69]
  wire  _GEN_5616 = io_wb_resps_0_valid ? _GEN_5520 : _GEN_2859; // @[rob.scala 346:69]
  wire  _GEN_5617 = io_wb_resps_0_valid ? _GEN_5521 : _GEN_2860; // @[rob.scala 346:69]
  wire  _GEN_5618 = io_wb_resps_0_valid ? _GEN_5522 : _GEN_2861; // @[rob.scala 346:69]
  wire  _GEN_5619 = io_wb_resps_0_valid ? _GEN_5523 : _GEN_2862; // @[rob.scala 346:69]
  wire  _GEN_5620 = io_wb_resps_0_valid ? _GEN_5524 : _GEN_2863; // @[rob.scala 346:69]
  wire  _GEN_5621 = io_wb_resps_0_valid ? _GEN_5525 : _GEN_2864; // @[rob.scala 346:69]
  wire  _GEN_5622 = io_wb_resps_0_valid ? _GEN_5526 : _GEN_2865; // @[rob.scala 346:69]
  wire  _GEN_5623 = io_wb_resps_0_valid ? _GEN_5527 : _GEN_2866; // @[rob.scala 346:69]
  wire  _GEN_5624 = io_wb_resps_0_valid ? _GEN_5528 : _GEN_2867; // @[rob.scala 346:69]
  wire  _GEN_5625 = io_wb_resps_0_valid ? _GEN_5529 : _GEN_2868; // @[rob.scala 346:69]
  wire  _GEN_5626 = io_wb_resps_0_valid ? _GEN_5530 : _GEN_2869; // @[rob.scala 346:69]
  wire  _GEN_5627 = io_wb_resps_0_valid ? _GEN_5531 : _GEN_2870; // @[rob.scala 346:69]
  wire  _GEN_5628 = io_wb_resps_0_valid ? _GEN_5532 : _GEN_2871; // @[rob.scala 346:69]
  wire  _GEN_5629 = io_wb_resps_0_valid ? _GEN_5533 : _GEN_2872; // @[rob.scala 346:69]
  wire  _GEN_5630 = io_wb_resps_0_valid ? _GEN_5534 : _GEN_2873; // @[rob.scala 346:69]
  wire  _GEN_5631 = io_wb_resps_0_valid ? _GEN_5535 : _GEN_2874; // @[rob.scala 346:69]
  wire  _GEN_5632 = io_wb_resps_0_valid ? _GEN_5536 : _GEN_2875; // @[rob.scala 346:69]
  wire  _GEN_5633 = io_wb_resps_0_valid ? _GEN_5537 : _GEN_2876; // @[rob.scala 346:69]
  wire  _GEN_5634 = io_wb_resps_0_valid ? _GEN_5538 : _GEN_2877; // @[rob.scala 346:69]
  wire  _GEN_5635 = io_wb_resps_0_valid ? _GEN_5539 : _GEN_2878; // @[rob.scala 346:69]
  wire  _GEN_5636 = io_wb_resps_0_valid ? _GEN_5540 : _GEN_2879; // @[rob.scala 346:69]
  wire  _GEN_5637 = io_wb_resps_0_valid ? _GEN_5541 : _GEN_2880; // @[rob.scala 346:69]
  wire  _GEN_5638 = io_wb_resps_0_valid ? _GEN_5542 : _GEN_2881; // @[rob.scala 346:69]
  wire  _GEN_5639 = io_wb_resps_0_valid ? _GEN_5543 : _GEN_2882; // @[rob.scala 346:69]
  wire  _GEN_5640 = io_wb_resps_0_valid ? _GEN_5544 : _GEN_2883; // @[rob.scala 346:69]
  wire  _GEN_5641 = io_wb_resps_0_valid ? _GEN_5545 : _GEN_2884; // @[rob.scala 346:69]
  wire  _GEN_5642 = io_wb_resps_0_valid ? _GEN_5546 : _GEN_2885; // @[rob.scala 346:69]
  wire  _GEN_5643 = io_wb_resps_0_valid ? _GEN_5547 : _GEN_5446; // @[rob.scala 346:69]
  wire  _GEN_5644 = io_wb_resps_0_valid ? _GEN_5548 : _GEN_5447; // @[rob.scala 346:69]
  wire  _GEN_5645 = io_wb_resps_0_valid ? _GEN_5549 : _GEN_5448; // @[rob.scala 346:69]
  wire  _GEN_5646 = io_wb_resps_0_valid ? _GEN_5550 : _GEN_5449; // @[rob.scala 346:69]
  wire  _GEN_5647 = io_wb_resps_0_valid ? _GEN_5551 : _GEN_5450; // @[rob.scala 346:69]
  wire  _GEN_5648 = io_wb_resps_0_valid ? _GEN_5552 : _GEN_5451; // @[rob.scala 346:69]
  wire  _GEN_5649 = io_wb_resps_0_valid ? _GEN_5553 : _GEN_5452; // @[rob.scala 346:69]
  wire  _GEN_5650 = io_wb_resps_0_valid ? _GEN_5554 : _GEN_5453; // @[rob.scala 346:69]
  wire  _GEN_5651 = io_wb_resps_0_valid ? _GEN_5555 : _GEN_5454; // @[rob.scala 346:69]
  wire  _GEN_5652 = io_wb_resps_0_valid ? _GEN_5556 : _GEN_5455; // @[rob.scala 346:69]
  wire  _GEN_5653 = io_wb_resps_0_valid ? _GEN_5557 : _GEN_5456; // @[rob.scala 346:69]
  wire  _GEN_5654 = io_wb_resps_0_valid ? _GEN_5558 : _GEN_5457; // @[rob.scala 346:69]
  wire  _GEN_5655 = io_wb_resps_0_valid ? _GEN_5559 : _GEN_5458; // @[rob.scala 346:69]
  wire  _GEN_5656 = io_wb_resps_0_valid ? _GEN_5560 : _GEN_5459; // @[rob.scala 346:69]
  wire  _GEN_5657 = io_wb_resps_0_valid ? _GEN_5561 : _GEN_5460; // @[rob.scala 346:69]
  wire  _GEN_5658 = io_wb_resps_0_valid ? _GEN_5562 : _GEN_5461; // @[rob.scala 346:69]
  wire  _GEN_5659 = io_wb_resps_0_valid ? _GEN_5563 : _GEN_5462; // @[rob.scala 346:69]
  wire  _GEN_5660 = io_wb_resps_0_valid ? _GEN_5564 : _GEN_5463; // @[rob.scala 346:69]
  wire  _GEN_5661 = io_wb_resps_0_valid ? _GEN_5565 : _GEN_5464; // @[rob.scala 346:69]
  wire  _GEN_5662 = io_wb_resps_0_valid ? _GEN_5566 : _GEN_5465; // @[rob.scala 346:69]
  wire  _GEN_5663 = io_wb_resps_0_valid ? _GEN_5567 : _GEN_5466; // @[rob.scala 346:69]
  wire  _GEN_5664 = io_wb_resps_0_valid ? _GEN_5568 : _GEN_5467; // @[rob.scala 346:69]
  wire  _GEN_5665 = io_wb_resps_0_valid ? _GEN_5569 : _GEN_5468; // @[rob.scala 346:69]
  wire  _GEN_5666 = io_wb_resps_0_valid ? _GEN_5570 : _GEN_5469; // @[rob.scala 346:69]
  wire  _GEN_5667 = io_wb_resps_0_valid ? _GEN_5571 : _GEN_5470; // @[rob.scala 346:69]
  wire  _GEN_5668 = io_wb_resps_0_valid ? _GEN_5572 : _GEN_5471; // @[rob.scala 346:69]
  wire  _GEN_5669 = io_wb_resps_0_valid ? _GEN_5573 : _GEN_5472; // @[rob.scala 346:69]
  wire  _GEN_5670 = io_wb_resps_0_valid ? _GEN_5574 : _GEN_5473; // @[rob.scala 346:69]
  wire  _GEN_5671 = io_wb_resps_0_valid ? _GEN_5575 : _GEN_5474; // @[rob.scala 346:69]
  wire  _GEN_5672 = io_wb_resps_0_valid ? _GEN_5576 : _GEN_5475; // @[rob.scala 346:69]
  wire  _GEN_5673 = io_wb_resps_0_valid ? _GEN_5577 : _GEN_5476; // @[rob.scala 346:69]
  wire  _GEN_5674 = io_wb_resps_0_valid ? _GEN_5578 : _GEN_5477; // @[rob.scala 346:69]
  wire  _GEN_5675 = 5'h0 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5579; // @[rob.scala 347:{31,31}]
  wire  _GEN_5676 = 5'h1 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5580; // @[rob.scala 347:{31,31}]
  wire  _GEN_5677 = 5'h2 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5581; // @[rob.scala 347:{31,31}]
  wire  _GEN_5678 = 5'h3 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5582; // @[rob.scala 347:{31,31}]
  wire  _GEN_5679 = 5'h4 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5583; // @[rob.scala 347:{31,31}]
  wire  _GEN_5680 = 5'h5 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5584; // @[rob.scala 347:{31,31}]
  wire  _GEN_5681 = 5'h6 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5585; // @[rob.scala 347:{31,31}]
  wire  _GEN_5682 = 5'h7 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5586; // @[rob.scala 347:{31,31}]
  wire  _GEN_5683 = 5'h8 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5587; // @[rob.scala 347:{31,31}]
  wire  _GEN_5684 = 5'h9 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5588; // @[rob.scala 347:{31,31}]
  wire  _GEN_5685 = 5'ha == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5589; // @[rob.scala 347:{31,31}]
  wire  _GEN_5686 = 5'hb == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5590; // @[rob.scala 347:{31,31}]
  wire  _GEN_5687 = 5'hc == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5591; // @[rob.scala 347:{31,31}]
  wire  _GEN_5688 = 5'hd == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5592; // @[rob.scala 347:{31,31}]
  wire  _GEN_5689 = 5'he == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5593; // @[rob.scala 347:{31,31}]
  wire  _GEN_5690 = 5'hf == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5594; // @[rob.scala 347:{31,31}]
  wire  _GEN_5691 = 5'h10 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5595; // @[rob.scala 347:{31,31}]
  wire  _GEN_5692 = 5'h11 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5596; // @[rob.scala 347:{31,31}]
  wire  _GEN_5693 = 5'h12 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5597; // @[rob.scala 347:{31,31}]
  wire  _GEN_5694 = 5'h13 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5598; // @[rob.scala 347:{31,31}]
  wire  _GEN_5695 = 5'h14 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5599; // @[rob.scala 347:{31,31}]
  wire  _GEN_5696 = 5'h15 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5600; // @[rob.scala 347:{31,31}]
  wire  _GEN_5697 = 5'h16 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5601; // @[rob.scala 347:{31,31}]
  wire  _GEN_5698 = 5'h17 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5602; // @[rob.scala 347:{31,31}]
  wire  _GEN_5699 = 5'h18 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5603; // @[rob.scala 347:{31,31}]
  wire  _GEN_5700 = 5'h19 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5604; // @[rob.scala 347:{31,31}]
  wire  _GEN_5701 = 5'h1a == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5605; // @[rob.scala 347:{31,31}]
  wire  _GEN_5702 = 5'h1b == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5606; // @[rob.scala 347:{31,31}]
  wire  _GEN_5703 = 5'h1c == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5607; // @[rob.scala 347:{31,31}]
  wire  _GEN_5704 = 5'h1d == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5608; // @[rob.scala 347:{31,31}]
  wire  _GEN_5705 = 5'h1e == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5609; // @[rob.scala 347:{31,31}]
  wire  _GEN_5706 = 5'h1f == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5610; // @[rob.scala 347:{31,31}]
  wire  _GEN_5707 = 5'h0 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5611; // @[rob.scala 348:{31,31}]
  wire  _GEN_5708 = 5'h1 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5612; // @[rob.scala 348:{31,31}]
  wire  _GEN_5709 = 5'h2 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5613; // @[rob.scala 348:{31,31}]
  wire  _GEN_5710 = 5'h3 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5614; // @[rob.scala 348:{31,31}]
  wire  _GEN_5711 = 5'h4 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5615; // @[rob.scala 348:{31,31}]
  wire  _GEN_5712 = 5'h5 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5616; // @[rob.scala 348:{31,31}]
  wire  _GEN_5713 = 5'h6 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5617; // @[rob.scala 348:{31,31}]
  wire  _GEN_5714 = 5'h7 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5618; // @[rob.scala 348:{31,31}]
  wire  _GEN_5715 = 5'h8 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5619; // @[rob.scala 348:{31,31}]
  wire  _GEN_5716 = 5'h9 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5620; // @[rob.scala 348:{31,31}]
  wire  _GEN_5717 = 5'ha == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5621; // @[rob.scala 348:{31,31}]
  wire  _GEN_5718 = 5'hb == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5622; // @[rob.scala 348:{31,31}]
  wire  _GEN_5719 = 5'hc == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5623; // @[rob.scala 348:{31,31}]
  wire  _GEN_5720 = 5'hd == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5624; // @[rob.scala 348:{31,31}]
  wire  _GEN_5721 = 5'he == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5625; // @[rob.scala 348:{31,31}]
  wire  _GEN_5722 = 5'hf == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5626; // @[rob.scala 348:{31,31}]
  wire  _GEN_5723 = 5'h10 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5627; // @[rob.scala 348:{31,31}]
  wire  _GEN_5724 = 5'h11 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5628; // @[rob.scala 348:{31,31}]
  wire  _GEN_5725 = 5'h12 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5629; // @[rob.scala 348:{31,31}]
  wire  _GEN_5726 = 5'h13 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5630; // @[rob.scala 348:{31,31}]
  wire  _GEN_5727 = 5'h14 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5631; // @[rob.scala 348:{31,31}]
  wire  _GEN_5728 = 5'h15 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5632; // @[rob.scala 348:{31,31}]
  wire  _GEN_5729 = 5'h16 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5633; // @[rob.scala 348:{31,31}]
  wire  _GEN_5730 = 5'h17 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5634; // @[rob.scala 348:{31,31}]
  wire  _GEN_5731 = 5'h18 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5635; // @[rob.scala 348:{31,31}]
  wire  _GEN_5732 = 5'h19 == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5636; // @[rob.scala 348:{31,31}]
  wire  _GEN_5733 = 5'h1a == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5637; // @[rob.scala 348:{31,31}]
  wire  _GEN_5734 = 5'h1b == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5638; // @[rob.scala 348:{31,31}]
  wire  _GEN_5735 = 5'h1c == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5639; // @[rob.scala 348:{31,31}]
  wire  _GEN_5736 = 5'h1d == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5640; // @[rob.scala 348:{31,31}]
  wire  _GEN_5737 = 5'h1e == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5641; // @[rob.scala 348:{31,31}]
  wire  _GEN_5738 = 5'h1f == io_wb_resps_1_bits_uop_rob_idx ? 1'h0 : _GEN_5642; // @[rob.scala 348:{31,31}]
  wire  _GEN_5739 = 5'h0 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5643; // @[rob.scala 349:{34,34}]
  wire  _GEN_5740 = 5'h1 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5644; // @[rob.scala 349:{34,34}]
  wire  _GEN_5741 = 5'h2 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5645; // @[rob.scala 349:{34,34}]
  wire  _GEN_5742 = 5'h3 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5646; // @[rob.scala 349:{34,34}]
  wire  _GEN_5743 = 5'h4 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5647; // @[rob.scala 349:{34,34}]
  wire  _GEN_5744 = 5'h5 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5648; // @[rob.scala 349:{34,34}]
  wire  _GEN_5745 = 5'h6 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5649; // @[rob.scala 349:{34,34}]
  wire  _GEN_5746 = 5'h7 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5650; // @[rob.scala 349:{34,34}]
  wire  _GEN_5747 = 5'h8 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5651; // @[rob.scala 349:{34,34}]
  wire  _GEN_5748 = 5'h9 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5652; // @[rob.scala 349:{34,34}]
  wire  _GEN_5749 = 5'ha == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5653; // @[rob.scala 349:{34,34}]
  wire  _GEN_5750 = 5'hb == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5654; // @[rob.scala 349:{34,34}]
  wire  _GEN_5751 = 5'hc == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5655; // @[rob.scala 349:{34,34}]
  wire  _GEN_5752 = 5'hd == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5656; // @[rob.scala 349:{34,34}]
  wire  _GEN_5753 = 5'he == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5657; // @[rob.scala 349:{34,34}]
  wire  _GEN_5754 = 5'hf == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5658; // @[rob.scala 349:{34,34}]
  wire  _GEN_5755 = 5'h10 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5659; // @[rob.scala 349:{34,34}]
  wire  _GEN_5756 = 5'h11 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5660; // @[rob.scala 349:{34,34}]
  wire  _GEN_5757 = 5'h12 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5661; // @[rob.scala 349:{34,34}]
  wire  _GEN_5758 = 5'h13 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5662; // @[rob.scala 349:{34,34}]
  wire  _GEN_5759 = 5'h14 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5663; // @[rob.scala 349:{34,34}]
  wire  _GEN_5760 = 5'h15 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5664; // @[rob.scala 349:{34,34}]
  wire  _GEN_5761 = 5'h16 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5665; // @[rob.scala 349:{34,34}]
  wire  _GEN_5762 = 5'h17 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5666; // @[rob.scala 349:{34,34}]
  wire  _GEN_5763 = 5'h18 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5667; // @[rob.scala 349:{34,34}]
  wire  _GEN_5764 = 5'h19 == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5668; // @[rob.scala 349:{34,34}]
  wire  _GEN_5765 = 5'h1a == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5669; // @[rob.scala 349:{34,34}]
  wire  _GEN_5766 = 5'h1b == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5670; // @[rob.scala 349:{34,34}]
  wire  _GEN_5767 = 5'h1c == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5671; // @[rob.scala 349:{34,34}]
  wire  _GEN_5768 = 5'h1d == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5672; // @[rob.scala 349:{34,34}]
  wire  _GEN_5769 = 5'h1e == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5673; // @[rob.scala 349:{34,34}]
  wire  _GEN_5770 = 5'h1f == io_wb_resps_1_bits_uop_rob_idx ? io_wb_resps_1_bits_predicated : _GEN_5674; // @[rob.scala 349:{34,34}]
  wire  _GEN_5771 = io_wb_resps_1_valid ? _GEN_5675 : _GEN_5579; // @[rob.scala 346:69]
  wire  _GEN_5772 = io_wb_resps_1_valid ? _GEN_5676 : _GEN_5580; // @[rob.scala 346:69]
  wire  _GEN_5773 = io_wb_resps_1_valid ? _GEN_5677 : _GEN_5581; // @[rob.scala 346:69]
  wire  _GEN_5774 = io_wb_resps_1_valid ? _GEN_5678 : _GEN_5582; // @[rob.scala 346:69]
  wire  _GEN_5775 = io_wb_resps_1_valid ? _GEN_5679 : _GEN_5583; // @[rob.scala 346:69]
  wire  _GEN_5776 = io_wb_resps_1_valid ? _GEN_5680 : _GEN_5584; // @[rob.scala 346:69]
  wire  _GEN_5777 = io_wb_resps_1_valid ? _GEN_5681 : _GEN_5585; // @[rob.scala 346:69]
  wire  _GEN_5778 = io_wb_resps_1_valid ? _GEN_5682 : _GEN_5586; // @[rob.scala 346:69]
  wire  _GEN_5779 = io_wb_resps_1_valid ? _GEN_5683 : _GEN_5587; // @[rob.scala 346:69]
  wire  _GEN_5780 = io_wb_resps_1_valid ? _GEN_5684 : _GEN_5588; // @[rob.scala 346:69]
  wire  _GEN_5781 = io_wb_resps_1_valid ? _GEN_5685 : _GEN_5589; // @[rob.scala 346:69]
  wire  _GEN_5782 = io_wb_resps_1_valid ? _GEN_5686 : _GEN_5590; // @[rob.scala 346:69]
  wire  _GEN_5783 = io_wb_resps_1_valid ? _GEN_5687 : _GEN_5591; // @[rob.scala 346:69]
  wire  _GEN_5784 = io_wb_resps_1_valid ? _GEN_5688 : _GEN_5592; // @[rob.scala 346:69]
  wire  _GEN_5785 = io_wb_resps_1_valid ? _GEN_5689 : _GEN_5593; // @[rob.scala 346:69]
  wire  _GEN_5786 = io_wb_resps_1_valid ? _GEN_5690 : _GEN_5594; // @[rob.scala 346:69]
  wire  _GEN_5787 = io_wb_resps_1_valid ? _GEN_5691 : _GEN_5595; // @[rob.scala 346:69]
  wire  _GEN_5788 = io_wb_resps_1_valid ? _GEN_5692 : _GEN_5596; // @[rob.scala 346:69]
  wire  _GEN_5789 = io_wb_resps_1_valid ? _GEN_5693 : _GEN_5597; // @[rob.scala 346:69]
  wire  _GEN_5790 = io_wb_resps_1_valid ? _GEN_5694 : _GEN_5598; // @[rob.scala 346:69]
  wire  _GEN_5791 = io_wb_resps_1_valid ? _GEN_5695 : _GEN_5599; // @[rob.scala 346:69]
  wire  _GEN_5792 = io_wb_resps_1_valid ? _GEN_5696 : _GEN_5600; // @[rob.scala 346:69]
  wire  _GEN_5793 = io_wb_resps_1_valid ? _GEN_5697 : _GEN_5601; // @[rob.scala 346:69]
  wire  _GEN_5794 = io_wb_resps_1_valid ? _GEN_5698 : _GEN_5602; // @[rob.scala 346:69]
  wire  _GEN_5795 = io_wb_resps_1_valid ? _GEN_5699 : _GEN_5603; // @[rob.scala 346:69]
  wire  _GEN_5796 = io_wb_resps_1_valid ? _GEN_5700 : _GEN_5604; // @[rob.scala 346:69]
  wire  _GEN_5797 = io_wb_resps_1_valid ? _GEN_5701 : _GEN_5605; // @[rob.scala 346:69]
  wire  _GEN_5798 = io_wb_resps_1_valid ? _GEN_5702 : _GEN_5606; // @[rob.scala 346:69]
  wire  _GEN_5799 = io_wb_resps_1_valid ? _GEN_5703 : _GEN_5607; // @[rob.scala 346:69]
  wire  _GEN_5800 = io_wb_resps_1_valid ? _GEN_5704 : _GEN_5608; // @[rob.scala 346:69]
  wire  _GEN_5801 = io_wb_resps_1_valid ? _GEN_5705 : _GEN_5609; // @[rob.scala 346:69]
  wire  _GEN_5802 = io_wb_resps_1_valid ? _GEN_5706 : _GEN_5610; // @[rob.scala 346:69]
  wire  _GEN_5803 = io_wb_resps_1_valid ? _GEN_5707 : _GEN_5611; // @[rob.scala 346:69]
  wire  _GEN_5804 = io_wb_resps_1_valid ? _GEN_5708 : _GEN_5612; // @[rob.scala 346:69]
  wire  _GEN_5805 = io_wb_resps_1_valid ? _GEN_5709 : _GEN_5613; // @[rob.scala 346:69]
  wire  _GEN_5806 = io_wb_resps_1_valid ? _GEN_5710 : _GEN_5614; // @[rob.scala 346:69]
  wire  _GEN_5807 = io_wb_resps_1_valid ? _GEN_5711 : _GEN_5615; // @[rob.scala 346:69]
  wire  _GEN_5808 = io_wb_resps_1_valid ? _GEN_5712 : _GEN_5616; // @[rob.scala 346:69]
  wire  _GEN_5809 = io_wb_resps_1_valid ? _GEN_5713 : _GEN_5617; // @[rob.scala 346:69]
  wire  _GEN_5810 = io_wb_resps_1_valid ? _GEN_5714 : _GEN_5618; // @[rob.scala 346:69]
  wire  _GEN_5811 = io_wb_resps_1_valid ? _GEN_5715 : _GEN_5619; // @[rob.scala 346:69]
  wire  _GEN_5812 = io_wb_resps_1_valid ? _GEN_5716 : _GEN_5620; // @[rob.scala 346:69]
  wire  _GEN_5813 = io_wb_resps_1_valid ? _GEN_5717 : _GEN_5621; // @[rob.scala 346:69]
  wire  _GEN_5814 = io_wb_resps_1_valid ? _GEN_5718 : _GEN_5622; // @[rob.scala 346:69]
  wire  _GEN_5815 = io_wb_resps_1_valid ? _GEN_5719 : _GEN_5623; // @[rob.scala 346:69]
  wire  _GEN_5816 = io_wb_resps_1_valid ? _GEN_5720 : _GEN_5624; // @[rob.scala 346:69]
  wire  _GEN_5817 = io_wb_resps_1_valid ? _GEN_5721 : _GEN_5625; // @[rob.scala 346:69]
  wire  _GEN_5818 = io_wb_resps_1_valid ? _GEN_5722 : _GEN_5626; // @[rob.scala 346:69]
  wire  _GEN_5819 = io_wb_resps_1_valid ? _GEN_5723 : _GEN_5627; // @[rob.scala 346:69]
  wire  _GEN_5820 = io_wb_resps_1_valid ? _GEN_5724 : _GEN_5628; // @[rob.scala 346:69]
  wire  _GEN_5821 = io_wb_resps_1_valid ? _GEN_5725 : _GEN_5629; // @[rob.scala 346:69]
  wire  _GEN_5822 = io_wb_resps_1_valid ? _GEN_5726 : _GEN_5630; // @[rob.scala 346:69]
  wire  _GEN_5823 = io_wb_resps_1_valid ? _GEN_5727 : _GEN_5631; // @[rob.scala 346:69]
  wire  _GEN_5824 = io_wb_resps_1_valid ? _GEN_5728 : _GEN_5632; // @[rob.scala 346:69]
  wire  _GEN_5825 = io_wb_resps_1_valid ? _GEN_5729 : _GEN_5633; // @[rob.scala 346:69]
  wire  _GEN_5826 = io_wb_resps_1_valid ? _GEN_5730 : _GEN_5634; // @[rob.scala 346:69]
  wire  _GEN_5827 = io_wb_resps_1_valid ? _GEN_5731 : _GEN_5635; // @[rob.scala 346:69]
  wire  _GEN_5828 = io_wb_resps_1_valid ? _GEN_5732 : _GEN_5636; // @[rob.scala 346:69]
  wire  _GEN_5829 = io_wb_resps_1_valid ? _GEN_5733 : _GEN_5637; // @[rob.scala 346:69]
  wire  _GEN_5830 = io_wb_resps_1_valid ? _GEN_5734 : _GEN_5638; // @[rob.scala 346:69]
  wire  _GEN_5831 = io_wb_resps_1_valid ? _GEN_5735 : _GEN_5639; // @[rob.scala 346:69]
  wire  _GEN_5832 = io_wb_resps_1_valid ? _GEN_5736 : _GEN_5640; // @[rob.scala 346:69]
  wire  _GEN_5833 = io_wb_resps_1_valid ? _GEN_5737 : _GEN_5641; // @[rob.scala 346:69]
  wire  _GEN_5834 = io_wb_resps_1_valid ? _GEN_5738 : _GEN_5642; // @[rob.scala 346:69]
  wire  _GEN_5835 = io_wb_resps_1_valid ? _GEN_5739 : _GEN_5643; // @[rob.scala 346:69]
  wire  _GEN_5836 = io_wb_resps_1_valid ? _GEN_5740 : _GEN_5644; // @[rob.scala 346:69]
  wire  _GEN_5837 = io_wb_resps_1_valid ? _GEN_5741 : _GEN_5645; // @[rob.scala 346:69]
  wire  _GEN_5838 = io_wb_resps_1_valid ? _GEN_5742 : _GEN_5646; // @[rob.scala 346:69]
  wire  _GEN_5839 = io_wb_resps_1_valid ? _GEN_5743 : _GEN_5647; // @[rob.scala 346:69]
  wire  _GEN_5840 = io_wb_resps_1_valid ? _GEN_5744 : _GEN_5648; // @[rob.scala 346:69]
  wire  _GEN_5841 = io_wb_resps_1_valid ? _GEN_5745 : _GEN_5649; // @[rob.scala 346:69]
  wire  _GEN_5842 = io_wb_resps_1_valid ? _GEN_5746 : _GEN_5650; // @[rob.scala 346:69]
  wire  _GEN_5843 = io_wb_resps_1_valid ? _GEN_5747 : _GEN_5651; // @[rob.scala 346:69]
  wire  _GEN_5844 = io_wb_resps_1_valid ? _GEN_5748 : _GEN_5652; // @[rob.scala 346:69]
  wire  _GEN_5845 = io_wb_resps_1_valid ? _GEN_5749 : _GEN_5653; // @[rob.scala 346:69]
  wire  _GEN_5846 = io_wb_resps_1_valid ? _GEN_5750 : _GEN_5654; // @[rob.scala 346:69]
  wire  _GEN_5847 = io_wb_resps_1_valid ? _GEN_5751 : _GEN_5655; // @[rob.scala 346:69]
  wire  _GEN_5848 = io_wb_resps_1_valid ? _GEN_5752 : _GEN_5656; // @[rob.scala 346:69]
  wire  _GEN_5849 = io_wb_resps_1_valid ? _GEN_5753 : _GEN_5657; // @[rob.scala 346:69]
  wire  _GEN_5850 = io_wb_resps_1_valid ? _GEN_5754 : _GEN_5658; // @[rob.scala 346:69]
  wire  _GEN_5851 = io_wb_resps_1_valid ? _GEN_5755 : _GEN_5659; // @[rob.scala 346:69]
  wire  _GEN_5852 = io_wb_resps_1_valid ? _GEN_5756 : _GEN_5660; // @[rob.scala 346:69]
  wire  _GEN_5853 = io_wb_resps_1_valid ? _GEN_5757 : _GEN_5661; // @[rob.scala 346:69]
  wire  _GEN_5854 = io_wb_resps_1_valid ? _GEN_5758 : _GEN_5662; // @[rob.scala 346:69]
  wire  _GEN_5855 = io_wb_resps_1_valid ? _GEN_5759 : _GEN_5663; // @[rob.scala 346:69]
  wire  _GEN_5856 = io_wb_resps_1_valid ? _GEN_5760 : _GEN_5664; // @[rob.scala 346:69]
  wire  _GEN_5857 = io_wb_resps_1_valid ? _GEN_5761 : _GEN_5665; // @[rob.scala 346:69]
  wire  _GEN_5858 = io_wb_resps_1_valid ? _GEN_5762 : _GEN_5666; // @[rob.scala 346:69]
  wire  _GEN_5859 = io_wb_resps_1_valid ? _GEN_5763 : _GEN_5667; // @[rob.scala 346:69]
  wire  _GEN_5860 = io_wb_resps_1_valid ? _GEN_5764 : _GEN_5668; // @[rob.scala 346:69]
  wire  _GEN_5861 = io_wb_resps_1_valid ? _GEN_5765 : _GEN_5669; // @[rob.scala 346:69]
  wire  _GEN_5862 = io_wb_resps_1_valid ? _GEN_5766 : _GEN_5670; // @[rob.scala 346:69]
  wire  _GEN_5863 = io_wb_resps_1_valid ? _GEN_5767 : _GEN_5671; // @[rob.scala 346:69]
  wire  _GEN_5864 = io_wb_resps_1_valid ? _GEN_5768 : _GEN_5672; // @[rob.scala 346:69]
  wire  _GEN_5865 = io_wb_resps_1_valid ? _GEN_5769 : _GEN_5673; // @[rob.scala 346:69]
  wire  _GEN_5866 = io_wb_resps_1_valid ? _GEN_5770 : _GEN_5674; // @[rob.scala 346:69]
  wire  _GEN_5867 = 5'h0 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5771; // @[rob.scala 347:{31,31}]
  wire  _GEN_5868 = 5'h1 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5772; // @[rob.scala 347:{31,31}]
  wire  _GEN_5869 = 5'h2 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5773; // @[rob.scala 347:{31,31}]
  wire  _GEN_5870 = 5'h3 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5774; // @[rob.scala 347:{31,31}]
  wire  _GEN_5871 = 5'h4 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5775; // @[rob.scala 347:{31,31}]
  wire  _GEN_5872 = 5'h5 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5776; // @[rob.scala 347:{31,31}]
  wire  _GEN_5873 = 5'h6 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5777; // @[rob.scala 347:{31,31}]
  wire  _GEN_5874 = 5'h7 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5778; // @[rob.scala 347:{31,31}]
  wire  _GEN_5875 = 5'h8 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5779; // @[rob.scala 347:{31,31}]
  wire  _GEN_5876 = 5'h9 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5780; // @[rob.scala 347:{31,31}]
  wire  _GEN_5877 = 5'ha == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5781; // @[rob.scala 347:{31,31}]
  wire  _GEN_5878 = 5'hb == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5782; // @[rob.scala 347:{31,31}]
  wire  _GEN_5879 = 5'hc == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5783; // @[rob.scala 347:{31,31}]
  wire  _GEN_5880 = 5'hd == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5784; // @[rob.scala 347:{31,31}]
  wire  _GEN_5881 = 5'he == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5785; // @[rob.scala 347:{31,31}]
  wire  _GEN_5882 = 5'hf == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5786; // @[rob.scala 347:{31,31}]
  wire  _GEN_5883 = 5'h10 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5787; // @[rob.scala 347:{31,31}]
  wire  _GEN_5884 = 5'h11 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5788; // @[rob.scala 347:{31,31}]
  wire  _GEN_5885 = 5'h12 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5789; // @[rob.scala 347:{31,31}]
  wire  _GEN_5886 = 5'h13 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5790; // @[rob.scala 347:{31,31}]
  wire  _GEN_5887 = 5'h14 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5791; // @[rob.scala 347:{31,31}]
  wire  _GEN_5888 = 5'h15 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5792; // @[rob.scala 347:{31,31}]
  wire  _GEN_5889 = 5'h16 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5793; // @[rob.scala 347:{31,31}]
  wire  _GEN_5890 = 5'h17 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5794; // @[rob.scala 347:{31,31}]
  wire  _GEN_5891 = 5'h18 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5795; // @[rob.scala 347:{31,31}]
  wire  _GEN_5892 = 5'h19 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5796; // @[rob.scala 347:{31,31}]
  wire  _GEN_5893 = 5'h1a == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5797; // @[rob.scala 347:{31,31}]
  wire  _GEN_5894 = 5'h1b == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5798; // @[rob.scala 347:{31,31}]
  wire  _GEN_5895 = 5'h1c == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5799; // @[rob.scala 347:{31,31}]
  wire  _GEN_5896 = 5'h1d == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5800; // @[rob.scala 347:{31,31}]
  wire  _GEN_5897 = 5'h1e == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5801; // @[rob.scala 347:{31,31}]
  wire  _GEN_5898 = 5'h1f == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5802; // @[rob.scala 347:{31,31}]
  wire  _GEN_5899 = 5'h0 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5803; // @[rob.scala 348:{31,31}]
  wire  _GEN_5900 = 5'h1 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5804; // @[rob.scala 348:{31,31}]
  wire  _GEN_5901 = 5'h2 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5805; // @[rob.scala 348:{31,31}]
  wire  _GEN_5902 = 5'h3 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5806; // @[rob.scala 348:{31,31}]
  wire  _GEN_5903 = 5'h4 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5807; // @[rob.scala 348:{31,31}]
  wire  _GEN_5904 = 5'h5 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5808; // @[rob.scala 348:{31,31}]
  wire  _GEN_5905 = 5'h6 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5809; // @[rob.scala 348:{31,31}]
  wire  _GEN_5906 = 5'h7 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5810; // @[rob.scala 348:{31,31}]
  wire  _GEN_5907 = 5'h8 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5811; // @[rob.scala 348:{31,31}]
  wire  _GEN_5908 = 5'h9 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5812; // @[rob.scala 348:{31,31}]
  wire  _GEN_5909 = 5'ha == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5813; // @[rob.scala 348:{31,31}]
  wire  _GEN_5910 = 5'hb == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5814; // @[rob.scala 348:{31,31}]
  wire  _GEN_5911 = 5'hc == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5815; // @[rob.scala 348:{31,31}]
  wire  _GEN_5912 = 5'hd == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5816; // @[rob.scala 348:{31,31}]
  wire  _GEN_5913 = 5'he == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5817; // @[rob.scala 348:{31,31}]
  wire  _GEN_5914 = 5'hf == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5818; // @[rob.scala 348:{31,31}]
  wire  _GEN_5915 = 5'h10 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5819; // @[rob.scala 348:{31,31}]
  wire  _GEN_5916 = 5'h11 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5820; // @[rob.scala 348:{31,31}]
  wire  _GEN_5917 = 5'h12 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5821; // @[rob.scala 348:{31,31}]
  wire  _GEN_5918 = 5'h13 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5822; // @[rob.scala 348:{31,31}]
  wire  _GEN_5919 = 5'h14 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5823; // @[rob.scala 348:{31,31}]
  wire  _GEN_5920 = 5'h15 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5824; // @[rob.scala 348:{31,31}]
  wire  _GEN_5921 = 5'h16 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5825; // @[rob.scala 348:{31,31}]
  wire  _GEN_5922 = 5'h17 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5826; // @[rob.scala 348:{31,31}]
  wire  _GEN_5923 = 5'h18 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5827; // @[rob.scala 348:{31,31}]
  wire  _GEN_5924 = 5'h19 == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5828; // @[rob.scala 348:{31,31}]
  wire  _GEN_5925 = 5'h1a == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5829; // @[rob.scala 348:{31,31}]
  wire  _GEN_5926 = 5'h1b == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5830; // @[rob.scala 348:{31,31}]
  wire  _GEN_5927 = 5'h1c == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5831; // @[rob.scala 348:{31,31}]
  wire  _GEN_5928 = 5'h1d == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5832; // @[rob.scala 348:{31,31}]
  wire  _GEN_5929 = 5'h1e == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5833; // @[rob.scala 348:{31,31}]
  wire  _GEN_5930 = 5'h1f == io_wb_resps_2_bits_uop_rob_idx ? 1'h0 : _GEN_5834; // @[rob.scala 348:{31,31}]
  wire  _GEN_5931 = 5'h0 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5835; // @[rob.scala 349:{34,34}]
  wire  _GEN_5932 = 5'h1 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5836; // @[rob.scala 349:{34,34}]
  wire  _GEN_5933 = 5'h2 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5837; // @[rob.scala 349:{34,34}]
  wire  _GEN_5934 = 5'h3 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5838; // @[rob.scala 349:{34,34}]
  wire  _GEN_5935 = 5'h4 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5839; // @[rob.scala 349:{34,34}]
  wire  _GEN_5936 = 5'h5 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5840; // @[rob.scala 349:{34,34}]
  wire  _GEN_5937 = 5'h6 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5841; // @[rob.scala 349:{34,34}]
  wire  _GEN_5938 = 5'h7 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5842; // @[rob.scala 349:{34,34}]
  wire  _GEN_5939 = 5'h8 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5843; // @[rob.scala 349:{34,34}]
  wire  _GEN_5940 = 5'h9 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5844; // @[rob.scala 349:{34,34}]
  wire  _GEN_5941 = 5'ha == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5845; // @[rob.scala 349:{34,34}]
  wire  _GEN_5942 = 5'hb == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5846; // @[rob.scala 349:{34,34}]
  wire  _GEN_5943 = 5'hc == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5847; // @[rob.scala 349:{34,34}]
  wire  _GEN_5944 = 5'hd == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5848; // @[rob.scala 349:{34,34}]
  wire  _GEN_5945 = 5'he == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5849; // @[rob.scala 349:{34,34}]
  wire  _GEN_5946 = 5'hf == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5850; // @[rob.scala 349:{34,34}]
  wire  _GEN_5947 = 5'h10 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5851; // @[rob.scala 349:{34,34}]
  wire  _GEN_5948 = 5'h11 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5852; // @[rob.scala 349:{34,34}]
  wire  _GEN_5949 = 5'h12 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5853; // @[rob.scala 349:{34,34}]
  wire  _GEN_5950 = 5'h13 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5854; // @[rob.scala 349:{34,34}]
  wire  _GEN_5951 = 5'h14 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5855; // @[rob.scala 349:{34,34}]
  wire  _GEN_5952 = 5'h15 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5856; // @[rob.scala 349:{34,34}]
  wire  _GEN_5953 = 5'h16 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5857; // @[rob.scala 349:{34,34}]
  wire  _GEN_5954 = 5'h17 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5858; // @[rob.scala 349:{34,34}]
  wire  _GEN_5955 = 5'h18 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5859; // @[rob.scala 349:{34,34}]
  wire  _GEN_5956 = 5'h19 == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5860; // @[rob.scala 349:{34,34}]
  wire  _GEN_5957 = 5'h1a == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5861; // @[rob.scala 349:{34,34}]
  wire  _GEN_5958 = 5'h1b == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5862; // @[rob.scala 349:{34,34}]
  wire  _GEN_5959 = 5'h1c == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5863; // @[rob.scala 349:{34,34}]
  wire  _GEN_5960 = 5'h1d == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5864; // @[rob.scala 349:{34,34}]
  wire  _GEN_5961 = 5'h1e == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5865; // @[rob.scala 349:{34,34}]
  wire  _GEN_5962 = 5'h1f == io_wb_resps_2_bits_uop_rob_idx ? io_wb_resps_2_bits_predicated : _GEN_5866; // @[rob.scala 349:{34,34}]
  wire  _GEN_5963 = io_wb_resps_2_valid ? _GEN_5867 : _GEN_5771; // @[rob.scala 346:69]
  wire  _GEN_5964 = io_wb_resps_2_valid ? _GEN_5868 : _GEN_5772; // @[rob.scala 346:69]
  wire  _GEN_5965 = io_wb_resps_2_valid ? _GEN_5869 : _GEN_5773; // @[rob.scala 346:69]
  wire  _GEN_5966 = io_wb_resps_2_valid ? _GEN_5870 : _GEN_5774; // @[rob.scala 346:69]
  wire  _GEN_5967 = io_wb_resps_2_valid ? _GEN_5871 : _GEN_5775; // @[rob.scala 346:69]
  wire  _GEN_5968 = io_wb_resps_2_valid ? _GEN_5872 : _GEN_5776; // @[rob.scala 346:69]
  wire  _GEN_5969 = io_wb_resps_2_valid ? _GEN_5873 : _GEN_5777; // @[rob.scala 346:69]
  wire  _GEN_5970 = io_wb_resps_2_valid ? _GEN_5874 : _GEN_5778; // @[rob.scala 346:69]
  wire  _GEN_5971 = io_wb_resps_2_valid ? _GEN_5875 : _GEN_5779; // @[rob.scala 346:69]
  wire  _GEN_5972 = io_wb_resps_2_valid ? _GEN_5876 : _GEN_5780; // @[rob.scala 346:69]
  wire  _GEN_5973 = io_wb_resps_2_valid ? _GEN_5877 : _GEN_5781; // @[rob.scala 346:69]
  wire  _GEN_5974 = io_wb_resps_2_valid ? _GEN_5878 : _GEN_5782; // @[rob.scala 346:69]
  wire  _GEN_5975 = io_wb_resps_2_valid ? _GEN_5879 : _GEN_5783; // @[rob.scala 346:69]
  wire  _GEN_5976 = io_wb_resps_2_valid ? _GEN_5880 : _GEN_5784; // @[rob.scala 346:69]
  wire  _GEN_5977 = io_wb_resps_2_valid ? _GEN_5881 : _GEN_5785; // @[rob.scala 346:69]
  wire  _GEN_5978 = io_wb_resps_2_valid ? _GEN_5882 : _GEN_5786; // @[rob.scala 346:69]
  wire  _GEN_5979 = io_wb_resps_2_valid ? _GEN_5883 : _GEN_5787; // @[rob.scala 346:69]
  wire  _GEN_5980 = io_wb_resps_2_valid ? _GEN_5884 : _GEN_5788; // @[rob.scala 346:69]
  wire  _GEN_5981 = io_wb_resps_2_valid ? _GEN_5885 : _GEN_5789; // @[rob.scala 346:69]
  wire  _GEN_5982 = io_wb_resps_2_valid ? _GEN_5886 : _GEN_5790; // @[rob.scala 346:69]
  wire  _GEN_5983 = io_wb_resps_2_valid ? _GEN_5887 : _GEN_5791; // @[rob.scala 346:69]
  wire  _GEN_5984 = io_wb_resps_2_valid ? _GEN_5888 : _GEN_5792; // @[rob.scala 346:69]
  wire  _GEN_5985 = io_wb_resps_2_valid ? _GEN_5889 : _GEN_5793; // @[rob.scala 346:69]
  wire  _GEN_5986 = io_wb_resps_2_valid ? _GEN_5890 : _GEN_5794; // @[rob.scala 346:69]
  wire  _GEN_5987 = io_wb_resps_2_valid ? _GEN_5891 : _GEN_5795; // @[rob.scala 346:69]
  wire  _GEN_5988 = io_wb_resps_2_valid ? _GEN_5892 : _GEN_5796; // @[rob.scala 346:69]
  wire  _GEN_5989 = io_wb_resps_2_valid ? _GEN_5893 : _GEN_5797; // @[rob.scala 346:69]
  wire  _GEN_5990 = io_wb_resps_2_valid ? _GEN_5894 : _GEN_5798; // @[rob.scala 346:69]
  wire  _GEN_5991 = io_wb_resps_2_valid ? _GEN_5895 : _GEN_5799; // @[rob.scala 346:69]
  wire  _GEN_5992 = io_wb_resps_2_valid ? _GEN_5896 : _GEN_5800; // @[rob.scala 346:69]
  wire  _GEN_5993 = io_wb_resps_2_valid ? _GEN_5897 : _GEN_5801; // @[rob.scala 346:69]
  wire  _GEN_5994 = io_wb_resps_2_valid ? _GEN_5898 : _GEN_5802; // @[rob.scala 346:69]
  wire  _GEN_5995 = io_wb_resps_2_valid ? _GEN_5899 : _GEN_5803; // @[rob.scala 346:69]
  wire  _GEN_5996 = io_wb_resps_2_valid ? _GEN_5900 : _GEN_5804; // @[rob.scala 346:69]
  wire  _GEN_5997 = io_wb_resps_2_valid ? _GEN_5901 : _GEN_5805; // @[rob.scala 346:69]
  wire  _GEN_5998 = io_wb_resps_2_valid ? _GEN_5902 : _GEN_5806; // @[rob.scala 346:69]
  wire  _GEN_5999 = io_wb_resps_2_valid ? _GEN_5903 : _GEN_5807; // @[rob.scala 346:69]
  wire  _GEN_6000 = io_wb_resps_2_valid ? _GEN_5904 : _GEN_5808; // @[rob.scala 346:69]
  wire  _GEN_6001 = io_wb_resps_2_valid ? _GEN_5905 : _GEN_5809; // @[rob.scala 346:69]
  wire  _GEN_6002 = io_wb_resps_2_valid ? _GEN_5906 : _GEN_5810; // @[rob.scala 346:69]
  wire  _GEN_6003 = io_wb_resps_2_valid ? _GEN_5907 : _GEN_5811; // @[rob.scala 346:69]
  wire  _GEN_6004 = io_wb_resps_2_valid ? _GEN_5908 : _GEN_5812; // @[rob.scala 346:69]
  wire  _GEN_6005 = io_wb_resps_2_valid ? _GEN_5909 : _GEN_5813; // @[rob.scala 346:69]
  wire  _GEN_6006 = io_wb_resps_2_valid ? _GEN_5910 : _GEN_5814; // @[rob.scala 346:69]
  wire  _GEN_6007 = io_wb_resps_2_valid ? _GEN_5911 : _GEN_5815; // @[rob.scala 346:69]
  wire  _GEN_6008 = io_wb_resps_2_valid ? _GEN_5912 : _GEN_5816; // @[rob.scala 346:69]
  wire  _GEN_6009 = io_wb_resps_2_valid ? _GEN_5913 : _GEN_5817; // @[rob.scala 346:69]
  wire  _GEN_6010 = io_wb_resps_2_valid ? _GEN_5914 : _GEN_5818; // @[rob.scala 346:69]
  wire  _GEN_6011 = io_wb_resps_2_valid ? _GEN_5915 : _GEN_5819; // @[rob.scala 346:69]
  wire  _GEN_6012 = io_wb_resps_2_valid ? _GEN_5916 : _GEN_5820; // @[rob.scala 346:69]
  wire  _GEN_6013 = io_wb_resps_2_valid ? _GEN_5917 : _GEN_5821; // @[rob.scala 346:69]
  wire  _GEN_6014 = io_wb_resps_2_valid ? _GEN_5918 : _GEN_5822; // @[rob.scala 346:69]
  wire  _GEN_6015 = io_wb_resps_2_valid ? _GEN_5919 : _GEN_5823; // @[rob.scala 346:69]
  wire  _GEN_6016 = io_wb_resps_2_valid ? _GEN_5920 : _GEN_5824; // @[rob.scala 346:69]
  wire  _GEN_6017 = io_wb_resps_2_valid ? _GEN_5921 : _GEN_5825; // @[rob.scala 346:69]
  wire  _GEN_6018 = io_wb_resps_2_valid ? _GEN_5922 : _GEN_5826; // @[rob.scala 346:69]
  wire  _GEN_6019 = io_wb_resps_2_valid ? _GEN_5923 : _GEN_5827; // @[rob.scala 346:69]
  wire  _GEN_6020 = io_wb_resps_2_valid ? _GEN_5924 : _GEN_5828; // @[rob.scala 346:69]
  wire  _GEN_6021 = io_wb_resps_2_valid ? _GEN_5925 : _GEN_5829; // @[rob.scala 346:69]
  wire  _GEN_6022 = io_wb_resps_2_valid ? _GEN_5926 : _GEN_5830; // @[rob.scala 346:69]
  wire  _GEN_6023 = io_wb_resps_2_valid ? _GEN_5927 : _GEN_5831; // @[rob.scala 346:69]
  wire  _GEN_6024 = io_wb_resps_2_valid ? _GEN_5928 : _GEN_5832; // @[rob.scala 346:69]
  wire  _GEN_6025 = io_wb_resps_2_valid ? _GEN_5929 : _GEN_5833; // @[rob.scala 346:69]
  wire  _GEN_6026 = io_wb_resps_2_valid ? _GEN_5930 : _GEN_5834; // @[rob.scala 346:69]
  wire  _GEN_6027 = io_wb_resps_2_valid ? _GEN_5931 : _GEN_5835; // @[rob.scala 346:69]
  wire  _GEN_6028 = io_wb_resps_2_valid ? _GEN_5932 : _GEN_5836; // @[rob.scala 346:69]
  wire  _GEN_6029 = io_wb_resps_2_valid ? _GEN_5933 : _GEN_5837; // @[rob.scala 346:69]
  wire  _GEN_6030 = io_wb_resps_2_valid ? _GEN_5934 : _GEN_5838; // @[rob.scala 346:69]
  wire  _GEN_6031 = io_wb_resps_2_valid ? _GEN_5935 : _GEN_5839; // @[rob.scala 346:69]
  wire  _GEN_6032 = io_wb_resps_2_valid ? _GEN_5936 : _GEN_5840; // @[rob.scala 346:69]
  wire  _GEN_6033 = io_wb_resps_2_valid ? _GEN_5937 : _GEN_5841; // @[rob.scala 346:69]
  wire  _GEN_6034 = io_wb_resps_2_valid ? _GEN_5938 : _GEN_5842; // @[rob.scala 346:69]
  wire  _GEN_6035 = io_wb_resps_2_valid ? _GEN_5939 : _GEN_5843; // @[rob.scala 346:69]
  wire  _GEN_6036 = io_wb_resps_2_valid ? _GEN_5940 : _GEN_5844; // @[rob.scala 346:69]
  wire  _GEN_6037 = io_wb_resps_2_valid ? _GEN_5941 : _GEN_5845; // @[rob.scala 346:69]
  wire  _GEN_6038 = io_wb_resps_2_valid ? _GEN_5942 : _GEN_5846; // @[rob.scala 346:69]
  wire  _GEN_6039 = io_wb_resps_2_valid ? _GEN_5943 : _GEN_5847; // @[rob.scala 346:69]
  wire  _GEN_6040 = io_wb_resps_2_valid ? _GEN_5944 : _GEN_5848; // @[rob.scala 346:69]
  wire  _GEN_6041 = io_wb_resps_2_valid ? _GEN_5945 : _GEN_5849; // @[rob.scala 346:69]
  wire  _GEN_6042 = io_wb_resps_2_valid ? _GEN_5946 : _GEN_5850; // @[rob.scala 346:69]
  wire  _GEN_6043 = io_wb_resps_2_valid ? _GEN_5947 : _GEN_5851; // @[rob.scala 346:69]
  wire  _GEN_6044 = io_wb_resps_2_valid ? _GEN_5948 : _GEN_5852; // @[rob.scala 346:69]
  wire  _GEN_6045 = io_wb_resps_2_valid ? _GEN_5949 : _GEN_5853; // @[rob.scala 346:69]
  wire  _GEN_6046 = io_wb_resps_2_valid ? _GEN_5950 : _GEN_5854; // @[rob.scala 346:69]
  wire  _GEN_6047 = io_wb_resps_2_valid ? _GEN_5951 : _GEN_5855; // @[rob.scala 346:69]
  wire  _GEN_6048 = io_wb_resps_2_valid ? _GEN_5952 : _GEN_5856; // @[rob.scala 346:69]
  wire  _GEN_6049 = io_wb_resps_2_valid ? _GEN_5953 : _GEN_5857; // @[rob.scala 346:69]
  wire  _GEN_6050 = io_wb_resps_2_valid ? _GEN_5954 : _GEN_5858; // @[rob.scala 346:69]
  wire  _GEN_6051 = io_wb_resps_2_valid ? _GEN_5955 : _GEN_5859; // @[rob.scala 346:69]
  wire  _GEN_6052 = io_wb_resps_2_valid ? _GEN_5956 : _GEN_5860; // @[rob.scala 346:69]
  wire  _GEN_6053 = io_wb_resps_2_valid ? _GEN_5957 : _GEN_5861; // @[rob.scala 346:69]
  wire  _GEN_6054 = io_wb_resps_2_valid ? _GEN_5958 : _GEN_5862; // @[rob.scala 346:69]
  wire  _GEN_6055 = io_wb_resps_2_valid ? _GEN_5959 : _GEN_5863; // @[rob.scala 346:69]
  wire  _GEN_6056 = io_wb_resps_2_valid ? _GEN_5960 : _GEN_5864; // @[rob.scala 346:69]
  wire  _GEN_6057 = io_wb_resps_2_valid ? _GEN_5961 : _GEN_5865; // @[rob.scala 346:69]
  wire  _GEN_6058 = io_wb_resps_2_valid ? _GEN_5962 : _GEN_5866; // @[rob.scala 346:69]
  wire  _GEN_6059 = 5'h0 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5963; // @[rob.scala 347:{31,31}]
  wire  _GEN_6060 = 5'h1 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5964; // @[rob.scala 347:{31,31}]
  wire  _GEN_6061 = 5'h2 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5965; // @[rob.scala 347:{31,31}]
  wire  _GEN_6062 = 5'h3 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5966; // @[rob.scala 347:{31,31}]
  wire  _GEN_6063 = 5'h4 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5967; // @[rob.scala 347:{31,31}]
  wire  _GEN_6064 = 5'h5 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5968; // @[rob.scala 347:{31,31}]
  wire  _GEN_6065 = 5'h6 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5969; // @[rob.scala 347:{31,31}]
  wire  _GEN_6066 = 5'h7 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5970; // @[rob.scala 347:{31,31}]
  wire  _GEN_6067 = 5'h8 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5971; // @[rob.scala 347:{31,31}]
  wire  _GEN_6068 = 5'h9 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5972; // @[rob.scala 347:{31,31}]
  wire  _GEN_6069 = 5'ha == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5973; // @[rob.scala 347:{31,31}]
  wire  _GEN_6070 = 5'hb == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5974; // @[rob.scala 347:{31,31}]
  wire  _GEN_6071 = 5'hc == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5975; // @[rob.scala 347:{31,31}]
  wire  _GEN_6072 = 5'hd == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5976; // @[rob.scala 347:{31,31}]
  wire  _GEN_6073 = 5'he == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5977; // @[rob.scala 347:{31,31}]
  wire  _GEN_6074 = 5'hf == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5978; // @[rob.scala 347:{31,31}]
  wire  _GEN_6075 = 5'h10 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5979; // @[rob.scala 347:{31,31}]
  wire  _GEN_6076 = 5'h11 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5980; // @[rob.scala 347:{31,31}]
  wire  _GEN_6077 = 5'h12 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5981; // @[rob.scala 347:{31,31}]
  wire  _GEN_6078 = 5'h13 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5982; // @[rob.scala 347:{31,31}]
  wire  _GEN_6079 = 5'h14 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5983; // @[rob.scala 347:{31,31}]
  wire  _GEN_6080 = 5'h15 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5984; // @[rob.scala 347:{31,31}]
  wire  _GEN_6081 = 5'h16 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5985; // @[rob.scala 347:{31,31}]
  wire  _GEN_6082 = 5'h17 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5986; // @[rob.scala 347:{31,31}]
  wire  _GEN_6083 = 5'h18 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5987; // @[rob.scala 347:{31,31}]
  wire  _GEN_6084 = 5'h19 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5988; // @[rob.scala 347:{31,31}]
  wire  _GEN_6085 = 5'h1a == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5989; // @[rob.scala 347:{31,31}]
  wire  _GEN_6086 = 5'h1b == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5990; // @[rob.scala 347:{31,31}]
  wire  _GEN_6087 = 5'h1c == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5991; // @[rob.scala 347:{31,31}]
  wire  _GEN_6088 = 5'h1d == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5992; // @[rob.scala 347:{31,31}]
  wire  _GEN_6089 = 5'h1e == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5993; // @[rob.scala 347:{31,31}]
  wire  _GEN_6090 = 5'h1f == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5994; // @[rob.scala 347:{31,31}]
  wire  _GEN_6091 = 5'h0 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5995; // @[rob.scala 348:{31,31}]
  wire  _GEN_6092 = 5'h1 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5996; // @[rob.scala 348:{31,31}]
  wire  _GEN_6093 = 5'h2 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5997; // @[rob.scala 348:{31,31}]
  wire  _GEN_6094 = 5'h3 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5998; // @[rob.scala 348:{31,31}]
  wire  _GEN_6095 = 5'h4 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_5999; // @[rob.scala 348:{31,31}]
  wire  _GEN_6096 = 5'h5 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6000; // @[rob.scala 348:{31,31}]
  wire  _GEN_6097 = 5'h6 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6001; // @[rob.scala 348:{31,31}]
  wire  _GEN_6098 = 5'h7 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6002; // @[rob.scala 348:{31,31}]
  wire  _GEN_6099 = 5'h8 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6003; // @[rob.scala 348:{31,31}]
  wire  _GEN_6100 = 5'h9 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6004; // @[rob.scala 348:{31,31}]
  wire  _GEN_6101 = 5'ha == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6005; // @[rob.scala 348:{31,31}]
  wire  _GEN_6102 = 5'hb == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6006; // @[rob.scala 348:{31,31}]
  wire  _GEN_6103 = 5'hc == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6007; // @[rob.scala 348:{31,31}]
  wire  _GEN_6104 = 5'hd == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6008; // @[rob.scala 348:{31,31}]
  wire  _GEN_6105 = 5'he == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6009; // @[rob.scala 348:{31,31}]
  wire  _GEN_6106 = 5'hf == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6010; // @[rob.scala 348:{31,31}]
  wire  _GEN_6107 = 5'h10 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6011; // @[rob.scala 348:{31,31}]
  wire  _GEN_6108 = 5'h11 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6012; // @[rob.scala 348:{31,31}]
  wire  _GEN_6109 = 5'h12 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6013; // @[rob.scala 348:{31,31}]
  wire  _GEN_6110 = 5'h13 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6014; // @[rob.scala 348:{31,31}]
  wire  _GEN_6111 = 5'h14 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6015; // @[rob.scala 348:{31,31}]
  wire  _GEN_6112 = 5'h15 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6016; // @[rob.scala 348:{31,31}]
  wire  _GEN_6113 = 5'h16 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6017; // @[rob.scala 348:{31,31}]
  wire  _GEN_6114 = 5'h17 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6018; // @[rob.scala 348:{31,31}]
  wire  _GEN_6115 = 5'h18 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6019; // @[rob.scala 348:{31,31}]
  wire  _GEN_6116 = 5'h19 == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6020; // @[rob.scala 348:{31,31}]
  wire  _GEN_6117 = 5'h1a == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6021; // @[rob.scala 348:{31,31}]
  wire  _GEN_6118 = 5'h1b == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6022; // @[rob.scala 348:{31,31}]
  wire  _GEN_6119 = 5'h1c == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6023; // @[rob.scala 348:{31,31}]
  wire  _GEN_6120 = 5'h1d == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6024; // @[rob.scala 348:{31,31}]
  wire  _GEN_6121 = 5'h1e == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6025; // @[rob.scala 348:{31,31}]
  wire  _GEN_6122 = 5'h1f == io_wb_resps_3_bits_uop_rob_idx ? 1'h0 : _GEN_6026; // @[rob.scala 348:{31,31}]
  wire  _GEN_6155 = io_wb_resps_3_valid ? _GEN_6059 : _GEN_5963; // @[rob.scala 346:69]
  wire  _GEN_6156 = io_wb_resps_3_valid ? _GEN_6060 : _GEN_5964; // @[rob.scala 346:69]
  wire  _GEN_6157 = io_wb_resps_3_valid ? _GEN_6061 : _GEN_5965; // @[rob.scala 346:69]
  wire  _GEN_6158 = io_wb_resps_3_valid ? _GEN_6062 : _GEN_5966; // @[rob.scala 346:69]
  wire  _GEN_6159 = io_wb_resps_3_valid ? _GEN_6063 : _GEN_5967; // @[rob.scala 346:69]
  wire  _GEN_6160 = io_wb_resps_3_valid ? _GEN_6064 : _GEN_5968; // @[rob.scala 346:69]
  wire  _GEN_6161 = io_wb_resps_3_valid ? _GEN_6065 : _GEN_5969; // @[rob.scala 346:69]
  wire  _GEN_6162 = io_wb_resps_3_valid ? _GEN_6066 : _GEN_5970; // @[rob.scala 346:69]
  wire  _GEN_6163 = io_wb_resps_3_valid ? _GEN_6067 : _GEN_5971; // @[rob.scala 346:69]
  wire  _GEN_6164 = io_wb_resps_3_valid ? _GEN_6068 : _GEN_5972; // @[rob.scala 346:69]
  wire  _GEN_6165 = io_wb_resps_3_valid ? _GEN_6069 : _GEN_5973; // @[rob.scala 346:69]
  wire  _GEN_6166 = io_wb_resps_3_valid ? _GEN_6070 : _GEN_5974; // @[rob.scala 346:69]
  wire  _GEN_6167 = io_wb_resps_3_valid ? _GEN_6071 : _GEN_5975; // @[rob.scala 346:69]
  wire  _GEN_6168 = io_wb_resps_3_valid ? _GEN_6072 : _GEN_5976; // @[rob.scala 346:69]
  wire  _GEN_6169 = io_wb_resps_3_valid ? _GEN_6073 : _GEN_5977; // @[rob.scala 346:69]
  wire  _GEN_6170 = io_wb_resps_3_valid ? _GEN_6074 : _GEN_5978; // @[rob.scala 346:69]
  wire  _GEN_6171 = io_wb_resps_3_valid ? _GEN_6075 : _GEN_5979; // @[rob.scala 346:69]
  wire  _GEN_6172 = io_wb_resps_3_valid ? _GEN_6076 : _GEN_5980; // @[rob.scala 346:69]
  wire  _GEN_6173 = io_wb_resps_3_valid ? _GEN_6077 : _GEN_5981; // @[rob.scala 346:69]
  wire  _GEN_6174 = io_wb_resps_3_valid ? _GEN_6078 : _GEN_5982; // @[rob.scala 346:69]
  wire  _GEN_6175 = io_wb_resps_3_valid ? _GEN_6079 : _GEN_5983; // @[rob.scala 346:69]
  wire  _GEN_6176 = io_wb_resps_3_valid ? _GEN_6080 : _GEN_5984; // @[rob.scala 346:69]
  wire  _GEN_6177 = io_wb_resps_3_valid ? _GEN_6081 : _GEN_5985; // @[rob.scala 346:69]
  wire  _GEN_6178 = io_wb_resps_3_valid ? _GEN_6082 : _GEN_5986; // @[rob.scala 346:69]
  wire  _GEN_6179 = io_wb_resps_3_valid ? _GEN_6083 : _GEN_5987; // @[rob.scala 346:69]
  wire  _GEN_6180 = io_wb_resps_3_valid ? _GEN_6084 : _GEN_5988; // @[rob.scala 346:69]
  wire  _GEN_6181 = io_wb_resps_3_valid ? _GEN_6085 : _GEN_5989; // @[rob.scala 346:69]
  wire  _GEN_6182 = io_wb_resps_3_valid ? _GEN_6086 : _GEN_5990; // @[rob.scala 346:69]
  wire  _GEN_6183 = io_wb_resps_3_valid ? _GEN_6087 : _GEN_5991; // @[rob.scala 346:69]
  wire  _GEN_6184 = io_wb_resps_3_valid ? _GEN_6088 : _GEN_5992; // @[rob.scala 346:69]
  wire  _GEN_6185 = io_wb_resps_3_valid ? _GEN_6089 : _GEN_5993; // @[rob.scala 346:69]
  wire  _GEN_6186 = io_wb_resps_3_valid ? _GEN_6090 : _GEN_5994; // @[rob.scala 346:69]
  wire  _GEN_6187 = io_wb_resps_3_valid ? _GEN_6091 : _GEN_5995; // @[rob.scala 346:69]
  wire  _GEN_6188 = io_wb_resps_3_valid ? _GEN_6092 : _GEN_5996; // @[rob.scala 346:69]
  wire  _GEN_6189 = io_wb_resps_3_valid ? _GEN_6093 : _GEN_5997; // @[rob.scala 346:69]
  wire  _GEN_6190 = io_wb_resps_3_valid ? _GEN_6094 : _GEN_5998; // @[rob.scala 346:69]
  wire  _GEN_6191 = io_wb_resps_3_valid ? _GEN_6095 : _GEN_5999; // @[rob.scala 346:69]
  wire  _GEN_6192 = io_wb_resps_3_valid ? _GEN_6096 : _GEN_6000; // @[rob.scala 346:69]
  wire  _GEN_6193 = io_wb_resps_3_valid ? _GEN_6097 : _GEN_6001; // @[rob.scala 346:69]
  wire  _GEN_6194 = io_wb_resps_3_valid ? _GEN_6098 : _GEN_6002; // @[rob.scala 346:69]
  wire  _GEN_6195 = io_wb_resps_3_valid ? _GEN_6099 : _GEN_6003; // @[rob.scala 346:69]
  wire  _GEN_6196 = io_wb_resps_3_valid ? _GEN_6100 : _GEN_6004; // @[rob.scala 346:69]
  wire  _GEN_6197 = io_wb_resps_3_valid ? _GEN_6101 : _GEN_6005; // @[rob.scala 346:69]
  wire  _GEN_6198 = io_wb_resps_3_valid ? _GEN_6102 : _GEN_6006; // @[rob.scala 346:69]
  wire  _GEN_6199 = io_wb_resps_3_valid ? _GEN_6103 : _GEN_6007; // @[rob.scala 346:69]
  wire  _GEN_6200 = io_wb_resps_3_valid ? _GEN_6104 : _GEN_6008; // @[rob.scala 346:69]
  wire  _GEN_6201 = io_wb_resps_3_valid ? _GEN_6105 : _GEN_6009; // @[rob.scala 346:69]
  wire  _GEN_6202 = io_wb_resps_3_valid ? _GEN_6106 : _GEN_6010; // @[rob.scala 346:69]
  wire  _GEN_6203 = io_wb_resps_3_valid ? _GEN_6107 : _GEN_6011; // @[rob.scala 346:69]
  wire  _GEN_6204 = io_wb_resps_3_valid ? _GEN_6108 : _GEN_6012; // @[rob.scala 346:69]
  wire  _GEN_6205 = io_wb_resps_3_valid ? _GEN_6109 : _GEN_6013; // @[rob.scala 346:69]
  wire  _GEN_6206 = io_wb_resps_3_valid ? _GEN_6110 : _GEN_6014; // @[rob.scala 346:69]
  wire  _GEN_6207 = io_wb_resps_3_valid ? _GEN_6111 : _GEN_6015; // @[rob.scala 346:69]
  wire  _GEN_6208 = io_wb_resps_3_valid ? _GEN_6112 : _GEN_6016; // @[rob.scala 346:69]
  wire  _GEN_6209 = io_wb_resps_3_valid ? _GEN_6113 : _GEN_6017; // @[rob.scala 346:69]
  wire  _GEN_6210 = io_wb_resps_3_valid ? _GEN_6114 : _GEN_6018; // @[rob.scala 346:69]
  wire  _GEN_6211 = io_wb_resps_3_valid ? _GEN_6115 : _GEN_6019; // @[rob.scala 346:69]
  wire  _GEN_6212 = io_wb_resps_3_valid ? _GEN_6116 : _GEN_6020; // @[rob.scala 346:69]
  wire  _GEN_6213 = io_wb_resps_3_valid ? _GEN_6117 : _GEN_6021; // @[rob.scala 346:69]
  wire  _GEN_6214 = io_wb_resps_3_valid ? _GEN_6118 : _GEN_6022; // @[rob.scala 346:69]
  wire  _GEN_6215 = io_wb_resps_3_valid ? _GEN_6119 : _GEN_6023; // @[rob.scala 346:69]
  wire  _GEN_6216 = io_wb_resps_3_valid ? _GEN_6120 : _GEN_6024; // @[rob.scala 346:69]
  wire  _GEN_6217 = io_wb_resps_3_valid ? _GEN_6121 : _GEN_6025; // @[rob.scala 346:69]
  wire  _GEN_6218 = io_wb_resps_3_valid ? _GEN_6122 : _GEN_6026; // @[rob.scala 346:69]
  wire  _GEN_6251 = 5'h0 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6155; // @[rob.scala 363:{26,26}]
  wire  _GEN_6252 = 5'h1 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6156; // @[rob.scala 363:{26,26}]
  wire  _GEN_6253 = 5'h2 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6157; // @[rob.scala 363:{26,26}]
  wire  _GEN_6254 = 5'h3 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6158; // @[rob.scala 363:{26,26}]
  wire  _GEN_6255 = 5'h4 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6159; // @[rob.scala 363:{26,26}]
  wire  _GEN_6256 = 5'h5 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6160; // @[rob.scala 363:{26,26}]
  wire  _GEN_6257 = 5'h6 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6161; // @[rob.scala 363:{26,26}]
  wire  _GEN_6258 = 5'h7 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6162; // @[rob.scala 363:{26,26}]
  wire  _GEN_6259 = 5'h8 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6163; // @[rob.scala 363:{26,26}]
  wire  _GEN_6260 = 5'h9 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6164; // @[rob.scala 363:{26,26}]
  wire  _GEN_6261 = 5'ha == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6165; // @[rob.scala 363:{26,26}]
  wire  _GEN_6262 = 5'hb == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6166; // @[rob.scala 363:{26,26}]
  wire  _GEN_6263 = 5'hc == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6167; // @[rob.scala 363:{26,26}]
  wire  _GEN_6264 = 5'hd == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6168; // @[rob.scala 363:{26,26}]
  wire  _GEN_6265 = 5'he == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6169; // @[rob.scala 363:{26,26}]
  wire  _GEN_6266 = 5'hf == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6170; // @[rob.scala 363:{26,26}]
  wire  _GEN_6267 = 5'h10 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6171; // @[rob.scala 363:{26,26}]
  wire  _GEN_6268 = 5'h11 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6172; // @[rob.scala 363:{26,26}]
  wire  _GEN_6269 = 5'h12 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6173; // @[rob.scala 363:{26,26}]
  wire  _GEN_6270 = 5'h13 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6174; // @[rob.scala 363:{26,26}]
  wire  _GEN_6271 = 5'h14 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6175; // @[rob.scala 363:{26,26}]
  wire  _GEN_6272 = 5'h15 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6176; // @[rob.scala 363:{26,26}]
  wire  _GEN_6273 = 5'h16 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6177; // @[rob.scala 363:{26,26}]
  wire  _GEN_6274 = 5'h17 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6178; // @[rob.scala 363:{26,26}]
  wire  _GEN_6275 = 5'h18 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6179; // @[rob.scala 363:{26,26}]
  wire  _GEN_6276 = 5'h19 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6180; // @[rob.scala 363:{26,26}]
  wire  _GEN_6277 = 5'h1a == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6181; // @[rob.scala 363:{26,26}]
  wire  _GEN_6278 = 5'h1b == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6182; // @[rob.scala 363:{26,26}]
  wire  _GEN_6279 = 5'h1c == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6183; // @[rob.scala 363:{26,26}]
  wire  _GEN_6280 = 5'h1d == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6184; // @[rob.scala 363:{26,26}]
  wire  _GEN_6281 = 5'h1e == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6185; // @[rob.scala 363:{26,26}]
  wire  _GEN_6282 = 5'h1f == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6186; // @[rob.scala 363:{26,26}]
  wire  _GEN_6283 = 5'h0 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6187; // @[rob.scala 364:{26,26}]
  wire  _GEN_6284 = 5'h1 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6188; // @[rob.scala 364:{26,26}]
  wire  _GEN_6285 = 5'h2 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6189; // @[rob.scala 364:{26,26}]
  wire  _GEN_6286 = 5'h3 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6190; // @[rob.scala 364:{26,26}]
  wire  _GEN_6287 = 5'h4 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6191; // @[rob.scala 364:{26,26}]
  wire  _GEN_6288 = 5'h5 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6192; // @[rob.scala 364:{26,26}]
  wire  _GEN_6289 = 5'h6 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6193; // @[rob.scala 364:{26,26}]
  wire  _GEN_6290 = 5'h7 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6194; // @[rob.scala 364:{26,26}]
  wire  _GEN_6291 = 5'h8 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6195; // @[rob.scala 364:{26,26}]
  wire  _GEN_6292 = 5'h9 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6196; // @[rob.scala 364:{26,26}]
  wire  _GEN_6293 = 5'ha == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6197; // @[rob.scala 364:{26,26}]
  wire  _GEN_6294 = 5'hb == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6198; // @[rob.scala 364:{26,26}]
  wire  _GEN_6295 = 5'hc == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6199; // @[rob.scala 364:{26,26}]
  wire  _GEN_6296 = 5'hd == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6200; // @[rob.scala 364:{26,26}]
  wire  _GEN_6297 = 5'he == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6201; // @[rob.scala 364:{26,26}]
  wire  _GEN_6298 = 5'hf == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6202; // @[rob.scala 364:{26,26}]
  wire  _GEN_6299 = 5'h10 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6203; // @[rob.scala 364:{26,26}]
  wire  _GEN_6300 = 5'h11 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6204; // @[rob.scala 364:{26,26}]
  wire  _GEN_6301 = 5'h12 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6205; // @[rob.scala 364:{26,26}]
  wire  _GEN_6302 = 5'h13 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6206; // @[rob.scala 364:{26,26}]
  wire  _GEN_6303 = 5'h14 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6207; // @[rob.scala 364:{26,26}]
  wire  _GEN_6304 = 5'h15 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6208; // @[rob.scala 364:{26,26}]
  wire  _GEN_6305 = 5'h16 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6209; // @[rob.scala 364:{26,26}]
  wire  _GEN_6306 = 5'h17 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6210; // @[rob.scala 364:{26,26}]
  wire  _GEN_6307 = 5'h18 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6211; // @[rob.scala 364:{26,26}]
  wire  _GEN_6308 = 5'h19 == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6212; // @[rob.scala 364:{26,26}]
  wire  _GEN_6309 = 5'h1a == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6213; // @[rob.scala 364:{26,26}]
  wire  _GEN_6310 = 5'h1b == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6214; // @[rob.scala 364:{26,26}]
  wire  _GEN_6311 = 5'h1c == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6215; // @[rob.scala 364:{26,26}]
  wire  _GEN_6312 = 5'h1d == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6216; // @[rob.scala 364:{26,26}]
  wire  _GEN_6313 = 5'h1e == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6217; // @[rob.scala 364:{26,26}]
  wire  _GEN_6314 = 5'h1f == io_lsu_clr_bsy_0_bits ? 1'h0 : _GEN_6218; // @[rob.scala 364:{26,26}]
  wire  _GEN_6316 = 5'h1 == io_lsu_clr_bsy_0_bits ? rob_val_1 : rob_val_0; // @[rob.scala 365:{31,31}]
  wire  _GEN_6317 = 5'h2 == io_lsu_clr_bsy_0_bits ? rob_val_2 : _GEN_6316; // @[rob.scala 365:{31,31}]
  wire  _GEN_6318 = 5'h3 == io_lsu_clr_bsy_0_bits ? rob_val_3 : _GEN_6317; // @[rob.scala 365:{31,31}]
  wire  _GEN_6319 = 5'h4 == io_lsu_clr_bsy_0_bits ? rob_val_4 : _GEN_6318; // @[rob.scala 365:{31,31}]
  wire  _GEN_6320 = 5'h5 == io_lsu_clr_bsy_0_bits ? rob_val_5 : _GEN_6319; // @[rob.scala 365:{31,31}]
  wire  _GEN_6321 = 5'h6 == io_lsu_clr_bsy_0_bits ? rob_val_6 : _GEN_6320; // @[rob.scala 365:{31,31}]
  wire  _GEN_6322 = 5'h7 == io_lsu_clr_bsy_0_bits ? rob_val_7 : _GEN_6321; // @[rob.scala 365:{31,31}]
  wire  _GEN_6323 = 5'h8 == io_lsu_clr_bsy_0_bits ? rob_val_8 : _GEN_6322; // @[rob.scala 365:{31,31}]
  wire  _GEN_6324 = 5'h9 == io_lsu_clr_bsy_0_bits ? rob_val_9 : _GEN_6323; // @[rob.scala 365:{31,31}]
  wire  _GEN_6325 = 5'ha == io_lsu_clr_bsy_0_bits ? rob_val_10 : _GEN_6324; // @[rob.scala 365:{31,31}]
  wire  _GEN_6326 = 5'hb == io_lsu_clr_bsy_0_bits ? rob_val_11 : _GEN_6325; // @[rob.scala 365:{31,31}]
  wire  _GEN_6327 = 5'hc == io_lsu_clr_bsy_0_bits ? rob_val_12 : _GEN_6326; // @[rob.scala 365:{31,31}]
  wire  _GEN_6328 = 5'hd == io_lsu_clr_bsy_0_bits ? rob_val_13 : _GEN_6327; // @[rob.scala 365:{31,31}]
  wire  _GEN_6329 = 5'he == io_lsu_clr_bsy_0_bits ? rob_val_14 : _GEN_6328; // @[rob.scala 365:{31,31}]
  wire  _GEN_6330 = 5'hf == io_lsu_clr_bsy_0_bits ? rob_val_15 : _GEN_6329; // @[rob.scala 365:{31,31}]
  wire  _GEN_6331 = 5'h10 == io_lsu_clr_bsy_0_bits ? rob_val_16 : _GEN_6330; // @[rob.scala 365:{31,31}]
  wire  _GEN_6332 = 5'h11 == io_lsu_clr_bsy_0_bits ? rob_val_17 : _GEN_6331; // @[rob.scala 365:{31,31}]
  wire  _GEN_6333 = 5'h12 == io_lsu_clr_bsy_0_bits ? rob_val_18 : _GEN_6332; // @[rob.scala 365:{31,31}]
  wire  _GEN_6334 = 5'h13 == io_lsu_clr_bsy_0_bits ? rob_val_19 : _GEN_6333; // @[rob.scala 365:{31,31}]
  wire  _GEN_6335 = 5'h14 == io_lsu_clr_bsy_0_bits ? rob_val_20 : _GEN_6334; // @[rob.scala 365:{31,31}]
  wire  _GEN_6336 = 5'h15 == io_lsu_clr_bsy_0_bits ? rob_val_21 : _GEN_6335; // @[rob.scala 365:{31,31}]
  wire  _GEN_6337 = 5'h16 == io_lsu_clr_bsy_0_bits ? rob_val_22 : _GEN_6336; // @[rob.scala 365:{31,31}]
  wire  _GEN_6338 = 5'h17 == io_lsu_clr_bsy_0_bits ? rob_val_23 : _GEN_6337; // @[rob.scala 365:{31,31}]
  wire  _GEN_6339 = 5'h18 == io_lsu_clr_bsy_0_bits ? rob_val_24 : _GEN_6338; // @[rob.scala 365:{31,31}]
  wire  _GEN_6340 = 5'h19 == io_lsu_clr_bsy_0_bits ? rob_val_25 : _GEN_6339; // @[rob.scala 365:{31,31}]
  wire  _GEN_6341 = 5'h1a == io_lsu_clr_bsy_0_bits ? rob_val_26 : _GEN_6340; // @[rob.scala 365:{31,31}]
  wire  _GEN_6342 = 5'h1b == io_lsu_clr_bsy_0_bits ? rob_val_27 : _GEN_6341; // @[rob.scala 365:{31,31}]
  wire  _GEN_6343 = 5'h1c == io_lsu_clr_bsy_0_bits ? rob_val_28 : _GEN_6342; // @[rob.scala 365:{31,31}]
  wire  _GEN_6344 = 5'h1d == io_lsu_clr_bsy_0_bits ? rob_val_29 : _GEN_6343; // @[rob.scala 365:{31,31}]
  wire  _GEN_6345 = 5'h1e == io_lsu_clr_bsy_0_bits ? rob_val_30 : _GEN_6344; // @[rob.scala 365:{31,31}]
  wire  _GEN_6346 = 5'h1f == io_lsu_clr_bsy_0_bits ? rob_val_31 : _GEN_6345; // @[rob.scala 365:{31,31}]
  wire  _GEN_6348 = 5'h1 == io_lsu_clr_bsy_0_bits ? rob_bsy_1 : rob_bsy_0; // @[rob.scala 366:{31,31}]
  wire  _GEN_6349 = 5'h2 == io_lsu_clr_bsy_0_bits ? rob_bsy_2 : _GEN_6348; // @[rob.scala 366:{31,31}]
  wire  _GEN_6350 = 5'h3 == io_lsu_clr_bsy_0_bits ? rob_bsy_3 : _GEN_6349; // @[rob.scala 366:{31,31}]
  wire  _GEN_6351 = 5'h4 == io_lsu_clr_bsy_0_bits ? rob_bsy_4 : _GEN_6350; // @[rob.scala 366:{31,31}]
  wire  _GEN_6352 = 5'h5 == io_lsu_clr_bsy_0_bits ? rob_bsy_5 : _GEN_6351; // @[rob.scala 366:{31,31}]
  wire  _GEN_6353 = 5'h6 == io_lsu_clr_bsy_0_bits ? rob_bsy_6 : _GEN_6352; // @[rob.scala 366:{31,31}]
  wire  _GEN_6354 = 5'h7 == io_lsu_clr_bsy_0_bits ? rob_bsy_7 : _GEN_6353; // @[rob.scala 366:{31,31}]
  wire  _GEN_6355 = 5'h8 == io_lsu_clr_bsy_0_bits ? rob_bsy_8 : _GEN_6354; // @[rob.scala 366:{31,31}]
  wire  _GEN_6356 = 5'h9 == io_lsu_clr_bsy_0_bits ? rob_bsy_9 : _GEN_6355; // @[rob.scala 366:{31,31}]
  wire  _GEN_6357 = 5'ha == io_lsu_clr_bsy_0_bits ? rob_bsy_10 : _GEN_6356; // @[rob.scala 366:{31,31}]
  wire  _GEN_6358 = 5'hb == io_lsu_clr_bsy_0_bits ? rob_bsy_11 : _GEN_6357; // @[rob.scala 366:{31,31}]
  wire  _GEN_6359 = 5'hc == io_lsu_clr_bsy_0_bits ? rob_bsy_12 : _GEN_6358; // @[rob.scala 366:{31,31}]
  wire  _GEN_6360 = 5'hd == io_lsu_clr_bsy_0_bits ? rob_bsy_13 : _GEN_6359; // @[rob.scala 366:{31,31}]
  wire  _GEN_6361 = 5'he == io_lsu_clr_bsy_0_bits ? rob_bsy_14 : _GEN_6360; // @[rob.scala 366:{31,31}]
  wire  _GEN_6362 = 5'hf == io_lsu_clr_bsy_0_bits ? rob_bsy_15 : _GEN_6361; // @[rob.scala 366:{31,31}]
  wire  _GEN_6363 = 5'h10 == io_lsu_clr_bsy_0_bits ? rob_bsy_16 : _GEN_6362; // @[rob.scala 366:{31,31}]
  wire  _GEN_6364 = 5'h11 == io_lsu_clr_bsy_0_bits ? rob_bsy_17 : _GEN_6363; // @[rob.scala 366:{31,31}]
  wire  _GEN_6365 = 5'h12 == io_lsu_clr_bsy_0_bits ? rob_bsy_18 : _GEN_6364; // @[rob.scala 366:{31,31}]
  wire  _GEN_6366 = 5'h13 == io_lsu_clr_bsy_0_bits ? rob_bsy_19 : _GEN_6365; // @[rob.scala 366:{31,31}]
  wire  _GEN_6367 = 5'h14 == io_lsu_clr_bsy_0_bits ? rob_bsy_20 : _GEN_6366; // @[rob.scala 366:{31,31}]
  wire  _GEN_6368 = 5'h15 == io_lsu_clr_bsy_0_bits ? rob_bsy_21 : _GEN_6367; // @[rob.scala 366:{31,31}]
  wire  _GEN_6369 = 5'h16 == io_lsu_clr_bsy_0_bits ? rob_bsy_22 : _GEN_6368; // @[rob.scala 366:{31,31}]
  wire  _GEN_6370 = 5'h17 == io_lsu_clr_bsy_0_bits ? rob_bsy_23 : _GEN_6369; // @[rob.scala 366:{31,31}]
  wire  _GEN_6371 = 5'h18 == io_lsu_clr_bsy_0_bits ? rob_bsy_24 : _GEN_6370; // @[rob.scala 366:{31,31}]
  wire  _GEN_6372 = 5'h19 == io_lsu_clr_bsy_0_bits ? rob_bsy_25 : _GEN_6371; // @[rob.scala 366:{31,31}]
  wire  _GEN_6373 = 5'h1a == io_lsu_clr_bsy_0_bits ? rob_bsy_26 : _GEN_6372; // @[rob.scala 366:{31,31}]
  wire  _GEN_6374 = 5'h1b == io_lsu_clr_bsy_0_bits ? rob_bsy_27 : _GEN_6373; // @[rob.scala 366:{31,31}]
  wire  _GEN_6375 = 5'h1c == io_lsu_clr_bsy_0_bits ? rob_bsy_28 : _GEN_6374; // @[rob.scala 366:{31,31}]
  wire  _GEN_6376 = 5'h1d == io_lsu_clr_bsy_0_bits ? rob_bsy_29 : _GEN_6375; // @[rob.scala 366:{31,31}]
  wire  _GEN_6377 = 5'h1e == io_lsu_clr_bsy_0_bits ? rob_bsy_30 : _GEN_6376; // @[rob.scala 366:{31,31}]
  wire  _GEN_6378 = 5'h1f == io_lsu_clr_bsy_0_bits ? rob_bsy_31 : _GEN_6377; // @[rob.scala 366:{31,31}]
  wire  _GEN_6379 = io_lsu_clr_bsy_0_valid ? _GEN_6251 : _GEN_6155; // @[rob.scala 361:75]
  wire  _GEN_6380 = io_lsu_clr_bsy_0_valid ? _GEN_6252 : _GEN_6156; // @[rob.scala 361:75]
  wire  _GEN_6381 = io_lsu_clr_bsy_0_valid ? _GEN_6253 : _GEN_6157; // @[rob.scala 361:75]
  wire  _GEN_6382 = io_lsu_clr_bsy_0_valid ? _GEN_6254 : _GEN_6158; // @[rob.scala 361:75]
  wire  _GEN_6383 = io_lsu_clr_bsy_0_valid ? _GEN_6255 : _GEN_6159; // @[rob.scala 361:75]
  wire  _GEN_6384 = io_lsu_clr_bsy_0_valid ? _GEN_6256 : _GEN_6160; // @[rob.scala 361:75]
  wire  _GEN_6385 = io_lsu_clr_bsy_0_valid ? _GEN_6257 : _GEN_6161; // @[rob.scala 361:75]
  wire  _GEN_6386 = io_lsu_clr_bsy_0_valid ? _GEN_6258 : _GEN_6162; // @[rob.scala 361:75]
  wire  _GEN_6387 = io_lsu_clr_bsy_0_valid ? _GEN_6259 : _GEN_6163; // @[rob.scala 361:75]
  wire  _GEN_6388 = io_lsu_clr_bsy_0_valid ? _GEN_6260 : _GEN_6164; // @[rob.scala 361:75]
  wire  _GEN_6389 = io_lsu_clr_bsy_0_valid ? _GEN_6261 : _GEN_6165; // @[rob.scala 361:75]
  wire  _GEN_6390 = io_lsu_clr_bsy_0_valid ? _GEN_6262 : _GEN_6166; // @[rob.scala 361:75]
  wire  _GEN_6391 = io_lsu_clr_bsy_0_valid ? _GEN_6263 : _GEN_6167; // @[rob.scala 361:75]
  wire  _GEN_6392 = io_lsu_clr_bsy_0_valid ? _GEN_6264 : _GEN_6168; // @[rob.scala 361:75]
  wire  _GEN_6393 = io_lsu_clr_bsy_0_valid ? _GEN_6265 : _GEN_6169; // @[rob.scala 361:75]
  wire  _GEN_6394 = io_lsu_clr_bsy_0_valid ? _GEN_6266 : _GEN_6170; // @[rob.scala 361:75]
  wire  _GEN_6395 = io_lsu_clr_bsy_0_valid ? _GEN_6267 : _GEN_6171; // @[rob.scala 361:75]
  wire  _GEN_6396 = io_lsu_clr_bsy_0_valid ? _GEN_6268 : _GEN_6172; // @[rob.scala 361:75]
  wire  _GEN_6397 = io_lsu_clr_bsy_0_valid ? _GEN_6269 : _GEN_6173; // @[rob.scala 361:75]
  wire  _GEN_6398 = io_lsu_clr_bsy_0_valid ? _GEN_6270 : _GEN_6174; // @[rob.scala 361:75]
  wire  _GEN_6399 = io_lsu_clr_bsy_0_valid ? _GEN_6271 : _GEN_6175; // @[rob.scala 361:75]
  wire  _GEN_6400 = io_lsu_clr_bsy_0_valid ? _GEN_6272 : _GEN_6176; // @[rob.scala 361:75]
  wire  _GEN_6401 = io_lsu_clr_bsy_0_valid ? _GEN_6273 : _GEN_6177; // @[rob.scala 361:75]
  wire  _GEN_6402 = io_lsu_clr_bsy_0_valid ? _GEN_6274 : _GEN_6178; // @[rob.scala 361:75]
  wire  _GEN_6403 = io_lsu_clr_bsy_0_valid ? _GEN_6275 : _GEN_6179; // @[rob.scala 361:75]
  wire  _GEN_6404 = io_lsu_clr_bsy_0_valid ? _GEN_6276 : _GEN_6180; // @[rob.scala 361:75]
  wire  _GEN_6405 = io_lsu_clr_bsy_0_valid ? _GEN_6277 : _GEN_6181; // @[rob.scala 361:75]
  wire  _GEN_6406 = io_lsu_clr_bsy_0_valid ? _GEN_6278 : _GEN_6182; // @[rob.scala 361:75]
  wire  _GEN_6407 = io_lsu_clr_bsy_0_valid ? _GEN_6279 : _GEN_6183; // @[rob.scala 361:75]
  wire  _GEN_6408 = io_lsu_clr_bsy_0_valid ? _GEN_6280 : _GEN_6184; // @[rob.scala 361:75]
  wire  _GEN_6409 = io_lsu_clr_bsy_0_valid ? _GEN_6281 : _GEN_6185; // @[rob.scala 361:75]
  wire  _GEN_6410 = io_lsu_clr_bsy_0_valid ? _GEN_6282 : _GEN_6186; // @[rob.scala 361:75]
  wire  _GEN_6411 = io_lsu_clr_bsy_0_valid ? _GEN_6283 : _GEN_6187; // @[rob.scala 361:75]
  wire  _GEN_6412 = io_lsu_clr_bsy_0_valid ? _GEN_6284 : _GEN_6188; // @[rob.scala 361:75]
  wire  _GEN_6413 = io_lsu_clr_bsy_0_valid ? _GEN_6285 : _GEN_6189; // @[rob.scala 361:75]
  wire  _GEN_6414 = io_lsu_clr_bsy_0_valid ? _GEN_6286 : _GEN_6190; // @[rob.scala 361:75]
  wire  _GEN_6415 = io_lsu_clr_bsy_0_valid ? _GEN_6287 : _GEN_6191; // @[rob.scala 361:75]
  wire  _GEN_6416 = io_lsu_clr_bsy_0_valid ? _GEN_6288 : _GEN_6192; // @[rob.scala 361:75]
  wire  _GEN_6417 = io_lsu_clr_bsy_0_valid ? _GEN_6289 : _GEN_6193; // @[rob.scala 361:75]
  wire  _GEN_6418 = io_lsu_clr_bsy_0_valid ? _GEN_6290 : _GEN_6194; // @[rob.scala 361:75]
  wire  _GEN_6419 = io_lsu_clr_bsy_0_valid ? _GEN_6291 : _GEN_6195; // @[rob.scala 361:75]
  wire  _GEN_6420 = io_lsu_clr_bsy_0_valid ? _GEN_6292 : _GEN_6196; // @[rob.scala 361:75]
  wire  _GEN_6421 = io_lsu_clr_bsy_0_valid ? _GEN_6293 : _GEN_6197; // @[rob.scala 361:75]
  wire  _GEN_6422 = io_lsu_clr_bsy_0_valid ? _GEN_6294 : _GEN_6198; // @[rob.scala 361:75]
  wire  _GEN_6423 = io_lsu_clr_bsy_0_valid ? _GEN_6295 : _GEN_6199; // @[rob.scala 361:75]
  wire  _GEN_6424 = io_lsu_clr_bsy_0_valid ? _GEN_6296 : _GEN_6200; // @[rob.scala 361:75]
  wire  _GEN_6425 = io_lsu_clr_bsy_0_valid ? _GEN_6297 : _GEN_6201; // @[rob.scala 361:75]
  wire  _GEN_6426 = io_lsu_clr_bsy_0_valid ? _GEN_6298 : _GEN_6202; // @[rob.scala 361:75]
  wire  _GEN_6427 = io_lsu_clr_bsy_0_valid ? _GEN_6299 : _GEN_6203; // @[rob.scala 361:75]
  wire  _GEN_6428 = io_lsu_clr_bsy_0_valid ? _GEN_6300 : _GEN_6204; // @[rob.scala 361:75]
  wire  _GEN_6429 = io_lsu_clr_bsy_0_valid ? _GEN_6301 : _GEN_6205; // @[rob.scala 361:75]
  wire  _GEN_6430 = io_lsu_clr_bsy_0_valid ? _GEN_6302 : _GEN_6206; // @[rob.scala 361:75]
  wire  _GEN_6431 = io_lsu_clr_bsy_0_valid ? _GEN_6303 : _GEN_6207; // @[rob.scala 361:75]
  wire  _GEN_6432 = io_lsu_clr_bsy_0_valid ? _GEN_6304 : _GEN_6208; // @[rob.scala 361:75]
  wire  _GEN_6433 = io_lsu_clr_bsy_0_valid ? _GEN_6305 : _GEN_6209; // @[rob.scala 361:75]
  wire  _GEN_6434 = io_lsu_clr_bsy_0_valid ? _GEN_6306 : _GEN_6210; // @[rob.scala 361:75]
  wire  _GEN_6435 = io_lsu_clr_bsy_0_valid ? _GEN_6307 : _GEN_6211; // @[rob.scala 361:75]
  wire  _GEN_6436 = io_lsu_clr_bsy_0_valid ? _GEN_6308 : _GEN_6212; // @[rob.scala 361:75]
  wire  _GEN_6437 = io_lsu_clr_bsy_0_valid ? _GEN_6309 : _GEN_6213; // @[rob.scala 361:75]
  wire  _GEN_6438 = io_lsu_clr_bsy_0_valid ? _GEN_6310 : _GEN_6214; // @[rob.scala 361:75]
  wire  _GEN_6439 = io_lsu_clr_bsy_0_valid ? _GEN_6311 : _GEN_6215; // @[rob.scala 361:75]
  wire  _GEN_6440 = io_lsu_clr_bsy_0_valid ? _GEN_6312 : _GEN_6216; // @[rob.scala 361:75]
  wire  _GEN_6441 = io_lsu_clr_bsy_0_valid ? _GEN_6313 : _GEN_6217; // @[rob.scala 361:75]
  wire  _GEN_6442 = io_lsu_clr_bsy_0_valid ? _GEN_6314 : _GEN_6218; // @[rob.scala 361:75]
  wire  _GEN_6475 = 5'h0 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6411; // @[rob.scala 364:{26,26}]
  wire  _GEN_6476 = 5'h1 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6412; // @[rob.scala 364:{26,26}]
  wire  _GEN_6477 = 5'h2 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6413; // @[rob.scala 364:{26,26}]
  wire  _GEN_6478 = 5'h3 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6414; // @[rob.scala 364:{26,26}]
  wire  _GEN_6479 = 5'h4 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6415; // @[rob.scala 364:{26,26}]
  wire  _GEN_6480 = 5'h5 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6416; // @[rob.scala 364:{26,26}]
  wire  _GEN_6481 = 5'h6 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6417; // @[rob.scala 364:{26,26}]
  wire  _GEN_6482 = 5'h7 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6418; // @[rob.scala 364:{26,26}]
  wire  _GEN_6483 = 5'h8 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6419; // @[rob.scala 364:{26,26}]
  wire  _GEN_6484 = 5'h9 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6420; // @[rob.scala 364:{26,26}]
  wire  _GEN_6485 = 5'ha == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6421; // @[rob.scala 364:{26,26}]
  wire  _GEN_6486 = 5'hb == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6422; // @[rob.scala 364:{26,26}]
  wire  _GEN_6487 = 5'hc == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6423; // @[rob.scala 364:{26,26}]
  wire  _GEN_6488 = 5'hd == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6424; // @[rob.scala 364:{26,26}]
  wire  _GEN_6489 = 5'he == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6425; // @[rob.scala 364:{26,26}]
  wire  _GEN_6490 = 5'hf == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6426; // @[rob.scala 364:{26,26}]
  wire  _GEN_6491 = 5'h10 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6427; // @[rob.scala 364:{26,26}]
  wire  _GEN_6492 = 5'h11 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6428; // @[rob.scala 364:{26,26}]
  wire  _GEN_6493 = 5'h12 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6429; // @[rob.scala 364:{26,26}]
  wire  _GEN_6494 = 5'h13 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6430; // @[rob.scala 364:{26,26}]
  wire  _GEN_6495 = 5'h14 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6431; // @[rob.scala 364:{26,26}]
  wire  _GEN_6496 = 5'h15 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6432; // @[rob.scala 364:{26,26}]
  wire  _GEN_6497 = 5'h16 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6433; // @[rob.scala 364:{26,26}]
  wire  _GEN_6498 = 5'h17 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6434; // @[rob.scala 364:{26,26}]
  wire  _GEN_6499 = 5'h18 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6435; // @[rob.scala 364:{26,26}]
  wire  _GEN_6500 = 5'h19 == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6436; // @[rob.scala 364:{26,26}]
  wire  _GEN_6501 = 5'h1a == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6437; // @[rob.scala 364:{26,26}]
  wire  _GEN_6502 = 5'h1b == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6438; // @[rob.scala 364:{26,26}]
  wire  _GEN_6503 = 5'h1c == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6439; // @[rob.scala 364:{26,26}]
  wire  _GEN_6504 = 5'h1d == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6440; // @[rob.scala 364:{26,26}]
  wire  _GEN_6505 = 5'h1e == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6441; // @[rob.scala 364:{26,26}]
  wire  _GEN_6506 = 5'h1f == io_lsu_clr_bsy_1_bits ? 1'h0 : _GEN_6442; // @[rob.scala 364:{26,26}]
  wire  _GEN_6508 = 5'h1 == io_lsu_clr_bsy_1_bits ? rob_val_1 : rob_val_0; // @[rob.scala 365:{31,31}]
  wire  _GEN_6509 = 5'h2 == io_lsu_clr_bsy_1_bits ? rob_val_2 : _GEN_6508; // @[rob.scala 365:{31,31}]
  wire  _GEN_6510 = 5'h3 == io_lsu_clr_bsy_1_bits ? rob_val_3 : _GEN_6509; // @[rob.scala 365:{31,31}]
  wire  _GEN_6511 = 5'h4 == io_lsu_clr_bsy_1_bits ? rob_val_4 : _GEN_6510; // @[rob.scala 365:{31,31}]
  wire  _GEN_6512 = 5'h5 == io_lsu_clr_bsy_1_bits ? rob_val_5 : _GEN_6511; // @[rob.scala 365:{31,31}]
  wire  _GEN_6513 = 5'h6 == io_lsu_clr_bsy_1_bits ? rob_val_6 : _GEN_6512; // @[rob.scala 365:{31,31}]
  wire  _GEN_6514 = 5'h7 == io_lsu_clr_bsy_1_bits ? rob_val_7 : _GEN_6513; // @[rob.scala 365:{31,31}]
  wire  _GEN_6515 = 5'h8 == io_lsu_clr_bsy_1_bits ? rob_val_8 : _GEN_6514; // @[rob.scala 365:{31,31}]
  wire  _GEN_6516 = 5'h9 == io_lsu_clr_bsy_1_bits ? rob_val_9 : _GEN_6515; // @[rob.scala 365:{31,31}]
  wire  _GEN_6517 = 5'ha == io_lsu_clr_bsy_1_bits ? rob_val_10 : _GEN_6516; // @[rob.scala 365:{31,31}]
  wire  _GEN_6518 = 5'hb == io_lsu_clr_bsy_1_bits ? rob_val_11 : _GEN_6517; // @[rob.scala 365:{31,31}]
  wire  _GEN_6519 = 5'hc == io_lsu_clr_bsy_1_bits ? rob_val_12 : _GEN_6518; // @[rob.scala 365:{31,31}]
  wire  _GEN_6520 = 5'hd == io_lsu_clr_bsy_1_bits ? rob_val_13 : _GEN_6519; // @[rob.scala 365:{31,31}]
  wire  _GEN_6521 = 5'he == io_lsu_clr_bsy_1_bits ? rob_val_14 : _GEN_6520; // @[rob.scala 365:{31,31}]
  wire  _GEN_6522 = 5'hf == io_lsu_clr_bsy_1_bits ? rob_val_15 : _GEN_6521; // @[rob.scala 365:{31,31}]
  wire  _GEN_6523 = 5'h10 == io_lsu_clr_bsy_1_bits ? rob_val_16 : _GEN_6522; // @[rob.scala 365:{31,31}]
  wire  _GEN_6524 = 5'h11 == io_lsu_clr_bsy_1_bits ? rob_val_17 : _GEN_6523; // @[rob.scala 365:{31,31}]
  wire  _GEN_6525 = 5'h12 == io_lsu_clr_bsy_1_bits ? rob_val_18 : _GEN_6524; // @[rob.scala 365:{31,31}]
  wire  _GEN_6526 = 5'h13 == io_lsu_clr_bsy_1_bits ? rob_val_19 : _GEN_6525; // @[rob.scala 365:{31,31}]
  wire  _GEN_6527 = 5'h14 == io_lsu_clr_bsy_1_bits ? rob_val_20 : _GEN_6526; // @[rob.scala 365:{31,31}]
  wire  _GEN_6528 = 5'h15 == io_lsu_clr_bsy_1_bits ? rob_val_21 : _GEN_6527; // @[rob.scala 365:{31,31}]
  wire  _GEN_6529 = 5'h16 == io_lsu_clr_bsy_1_bits ? rob_val_22 : _GEN_6528; // @[rob.scala 365:{31,31}]
  wire  _GEN_6530 = 5'h17 == io_lsu_clr_bsy_1_bits ? rob_val_23 : _GEN_6529; // @[rob.scala 365:{31,31}]
  wire  _GEN_6531 = 5'h18 == io_lsu_clr_bsy_1_bits ? rob_val_24 : _GEN_6530; // @[rob.scala 365:{31,31}]
  wire  _GEN_6532 = 5'h19 == io_lsu_clr_bsy_1_bits ? rob_val_25 : _GEN_6531; // @[rob.scala 365:{31,31}]
  wire  _GEN_6533 = 5'h1a == io_lsu_clr_bsy_1_bits ? rob_val_26 : _GEN_6532; // @[rob.scala 365:{31,31}]
  wire  _GEN_6534 = 5'h1b == io_lsu_clr_bsy_1_bits ? rob_val_27 : _GEN_6533; // @[rob.scala 365:{31,31}]
  wire  _GEN_6535 = 5'h1c == io_lsu_clr_bsy_1_bits ? rob_val_28 : _GEN_6534; // @[rob.scala 365:{31,31}]
  wire  _GEN_6536 = 5'h1d == io_lsu_clr_bsy_1_bits ? rob_val_29 : _GEN_6535; // @[rob.scala 365:{31,31}]
  wire  _GEN_6537 = 5'h1e == io_lsu_clr_bsy_1_bits ? rob_val_30 : _GEN_6536; // @[rob.scala 365:{31,31}]
  wire  _GEN_6538 = 5'h1f == io_lsu_clr_bsy_1_bits ? rob_val_31 : _GEN_6537; // @[rob.scala 365:{31,31}]
  wire  _GEN_6540 = 5'h1 == io_lsu_clr_bsy_1_bits ? rob_bsy_1 : rob_bsy_0; // @[rob.scala 366:{31,31}]
  wire  _GEN_6541 = 5'h2 == io_lsu_clr_bsy_1_bits ? rob_bsy_2 : _GEN_6540; // @[rob.scala 366:{31,31}]
  wire  _GEN_6542 = 5'h3 == io_lsu_clr_bsy_1_bits ? rob_bsy_3 : _GEN_6541; // @[rob.scala 366:{31,31}]
  wire  _GEN_6543 = 5'h4 == io_lsu_clr_bsy_1_bits ? rob_bsy_4 : _GEN_6542; // @[rob.scala 366:{31,31}]
  wire  _GEN_6544 = 5'h5 == io_lsu_clr_bsy_1_bits ? rob_bsy_5 : _GEN_6543; // @[rob.scala 366:{31,31}]
  wire  _GEN_6545 = 5'h6 == io_lsu_clr_bsy_1_bits ? rob_bsy_6 : _GEN_6544; // @[rob.scala 366:{31,31}]
  wire  _GEN_6546 = 5'h7 == io_lsu_clr_bsy_1_bits ? rob_bsy_7 : _GEN_6545; // @[rob.scala 366:{31,31}]
  wire  _GEN_6547 = 5'h8 == io_lsu_clr_bsy_1_bits ? rob_bsy_8 : _GEN_6546; // @[rob.scala 366:{31,31}]
  wire  _GEN_6548 = 5'h9 == io_lsu_clr_bsy_1_bits ? rob_bsy_9 : _GEN_6547; // @[rob.scala 366:{31,31}]
  wire  _GEN_6549 = 5'ha == io_lsu_clr_bsy_1_bits ? rob_bsy_10 : _GEN_6548; // @[rob.scala 366:{31,31}]
  wire  _GEN_6550 = 5'hb == io_lsu_clr_bsy_1_bits ? rob_bsy_11 : _GEN_6549; // @[rob.scala 366:{31,31}]
  wire  _GEN_6551 = 5'hc == io_lsu_clr_bsy_1_bits ? rob_bsy_12 : _GEN_6550; // @[rob.scala 366:{31,31}]
  wire  _GEN_6552 = 5'hd == io_lsu_clr_bsy_1_bits ? rob_bsy_13 : _GEN_6551; // @[rob.scala 366:{31,31}]
  wire  _GEN_6553 = 5'he == io_lsu_clr_bsy_1_bits ? rob_bsy_14 : _GEN_6552; // @[rob.scala 366:{31,31}]
  wire  _GEN_6554 = 5'hf == io_lsu_clr_bsy_1_bits ? rob_bsy_15 : _GEN_6553; // @[rob.scala 366:{31,31}]
  wire  _GEN_6555 = 5'h10 == io_lsu_clr_bsy_1_bits ? rob_bsy_16 : _GEN_6554; // @[rob.scala 366:{31,31}]
  wire  _GEN_6556 = 5'h11 == io_lsu_clr_bsy_1_bits ? rob_bsy_17 : _GEN_6555; // @[rob.scala 366:{31,31}]
  wire  _GEN_6557 = 5'h12 == io_lsu_clr_bsy_1_bits ? rob_bsy_18 : _GEN_6556; // @[rob.scala 366:{31,31}]
  wire  _GEN_6558 = 5'h13 == io_lsu_clr_bsy_1_bits ? rob_bsy_19 : _GEN_6557; // @[rob.scala 366:{31,31}]
  wire  _GEN_6559 = 5'h14 == io_lsu_clr_bsy_1_bits ? rob_bsy_20 : _GEN_6558; // @[rob.scala 366:{31,31}]
  wire  _GEN_6560 = 5'h15 == io_lsu_clr_bsy_1_bits ? rob_bsy_21 : _GEN_6559; // @[rob.scala 366:{31,31}]
  wire  _GEN_6561 = 5'h16 == io_lsu_clr_bsy_1_bits ? rob_bsy_22 : _GEN_6560; // @[rob.scala 366:{31,31}]
  wire  _GEN_6562 = 5'h17 == io_lsu_clr_bsy_1_bits ? rob_bsy_23 : _GEN_6561; // @[rob.scala 366:{31,31}]
  wire  _GEN_6563 = 5'h18 == io_lsu_clr_bsy_1_bits ? rob_bsy_24 : _GEN_6562; // @[rob.scala 366:{31,31}]
  wire  _GEN_6564 = 5'h19 == io_lsu_clr_bsy_1_bits ? rob_bsy_25 : _GEN_6563; // @[rob.scala 366:{31,31}]
  wire  _GEN_6565 = 5'h1a == io_lsu_clr_bsy_1_bits ? rob_bsy_26 : _GEN_6564; // @[rob.scala 366:{31,31}]
  wire  _GEN_6566 = 5'h1b == io_lsu_clr_bsy_1_bits ? rob_bsy_27 : _GEN_6565; // @[rob.scala 366:{31,31}]
  wire  _GEN_6567 = 5'h1c == io_lsu_clr_bsy_1_bits ? rob_bsy_28 : _GEN_6566; // @[rob.scala 366:{31,31}]
  wire  _GEN_6568 = 5'h1d == io_lsu_clr_bsy_1_bits ? rob_bsy_29 : _GEN_6567; // @[rob.scala 366:{31,31}]
  wire  _GEN_6569 = 5'h1e == io_lsu_clr_bsy_1_bits ? rob_bsy_30 : _GEN_6568; // @[rob.scala 366:{31,31}]
  wire  _GEN_6570 = 5'h1f == io_lsu_clr_bsy_1_bits ? rob_bsy_31 : _GEN_6569; // @[rob.scala 366:{31,31}]
  wire  _GEN_6603 = io_lsu_clr_bsy_1_valid ? _GEN_6475 : _GEN_6411; // @[rob.scala 361:75]
  wire  _GEN_6604 = io_lsu_clr_bsy_1_valid ? _GEN_6476 : _GEN_6412; // @[rob.scala 361:75]
  wire  _GEN_6605 = io_lsu_clr_bsy_1_valid ? _GEN_6477 : _GEN_6413; // @[rob.scala 361:75]
  wire  _GEN_6606 = io_lsu_clr_bsy_1_valid ? _GEN_6478 : _GEN_6414; // @[rob.scala 361:75]
  wire  _GEN_6607 = io_lsu_clr_bsy_1_valid ? _GEN_6479 : _GEN_6415; // @[rob.scala 361:75]
  wire  _GEN_6608 = io_lsu_clr_bsy_1_valid ? _GEN_6480 : _GEN_6416; // @[rob.scala 361:75]
  wire  _GEN_6609 = io_lsu_clr_bsy_1_valid ? _GEN_6481 : _GEN_6417; // @[rob.scala 361:75]
  wire  _GEN_6610 = io_lsu_clr_bsy_1_valid ? _GEN_6482 : _GEN_6418; // @[rob.scala 361:75]
  wire  _GEN_6611 = io_lsu_clr_bsy_1_valid ? _GEN_6483 : _GEN_6419; // @[rob.scala 361:75]
  wire  _GEN_6612 = io_lsu_clr_bsy_1_valid ? _GEN_6484 : _GEN_6420; // @[rob.scala 361:75]
  wire  _GEN_6613 = io_lsu_clr_bsy_1_valid ? _GEN_6485 : _GEN_6421; // @[rob.scala 361:75]
  wire  _GEN_6614 = io_lsu_clr_bsy_1_valid ? _GEN_6486 : _GEN_6422; // @[rob.scala 361:75]
  wire  _GEN_6615 = io_lsu_clr_bsy_1_valid ? _GEN_6487 : _GEN_6423; // @[rob.scala 361:75]
  wire  _GEN_6616 = io_lsu_clr_bsy_1_valid ? _GEN_6488 : _GEN_6424; // @[rob.scala 361:75]
  wire  _GEN_6617 = io_lsu_clr_bsy_1_valid ? _GEN_6489 : _GEN_6425; // @[rob.scala 361:75]
  wire  _GEN_6618 = io_lsu_clr_bsy_1_valid ? _GEN_6490 : _GEN_6426; // @[rob.scala 361:75]
  wire  _GEN_6619 = io_lsu_clr_bsy_1_valid ? _GEN_6491 : _GEN_6427; // @[rob.scala 361:75]
  wire  _GEN_6620 = io_lsu_clr_bsy_1_valid ? _GEN_6492 : _GEN_6428; // @[rob.scala 361:75]
  wire  _GEN_6621 = io_lsu_clr_bsy_1_valid ? _GEN_6493 : _GEN_6429; // @[rob.scala 361:75]
  wire  _GEN_6622 = io_lsu_clr_bsy_1_valid ? _GEN_6494 : _GEN_6430; // @[rob.scala 361:75]
  wire  _GEN_6623 = io_lsu_clr_bsy_1_valid ? _GEN_6495 : _GEN_6431; // @[rob.scala 361:75]
  wire  _GEN_6624 = io_lsu_clr_bsy_1_valid ? _GEN_6496 : _GEN_6432; // @[rob.scala 361:75]
  wire  _GEN_6625 = io_lsu_clr_bsy_1_valid ? _GEN_6497 : _GEN_6433; // @[rob.scala 361:75]
  wire  _GEN_6626 = io_lsu_clr_bsy_1_valid ? _GEN_6498 : _GEN_6434; // @[rob.scala 361:75]
  wire  _GEN_6627 = io_lsu_clr_bsy_1_valid ? _GEN_6499 : _GEN_6435; // @[rob.scala 361:75]
  wire  _GEN_6628 = io_lsu_clr_bsy_1_valid ? _GEN_6500 : _GEN_6436; // @[rob.scala 361:75]
  wire  _GEN_6629 = io_lsu_clr_bsy_1_valid ? _GEN_6501 : _GEN_6437; // @[rob.scala 361:75]
  wire  _GEN_6630 = io_lsu_clr_bsy_1_valid ? _GEN_6502 : _GEN_6438; // @[rob.scala 361:75]
  wire  _GEN_6631 = io_lsu_clr_bsy_1_valid ? _GEN_6503 : _GEN_6439; // @[rob.scala 361:75]
  wire  _GEN_6632 = io_lsu_clr_bsy_1_valid ? _GEN_6504 : _GEN_6440; // @[rob.scala 361:75]
  wire  _GEN_6633 = io_lsu_clr_bsy_1_valid ? _GEN_6505 : _GEN_6441; // @[rob.scala 361:75]
  wire  _GEN_6634 = io_lsu_clr_bsy_1_valid ? _GEN_6506 : _GEN_6442; // @[rob.scala 361:75]
  wire  _GEN_6709 = 5'h0 == io_lxcpt_bits_uop_rob_idx | _GEN_5414; // @[rob.scala 391:{59,59}]
  wire  _GEN_6710 = 5'h1 == io_lxcpt_bits_uop_rob_idx | _GEN_5415; // @[rob.scala 391:{59,59}]
  wire  _GEN_6711 = 5'h2 == io_lxcpt_bits_uop_rob_idx | _GEN_5416; // @[rob.scala 391:{59,59}]
  wire  _GEN_6712 = 5'h3 == io_lxcpt_bits_uop_rob_idx | _GEN_5417; // @[rob.scala 391:{59,59}]
  wire  _GEN_6713 = 5'h4 == io_lxcpt_bits_uop_rob_idx | _GEN_5418; // @[rob.scala 391:{59,59}]
  wire  _GEN_6714 = 5'h5 == io_lxcpt_bits_uop_rob_idx | _GEN_5419; // @[rob.scala 391:{59,59}]
  wire  _GEN_6715 = 5'h6 == io_lxcpt_bits_uop_rob_idx | _GEN_5420; // @[rob.scala 391:{59,59}]
  wire  _GEN_6716 = 5'h7 == io_lxcpt_bits_uop_rob_idx | _GEN_5421; // @[rob.scala 391:{59,59}]
  wire  _GEN_6717 = 5'h8 == io_lxcpt_bits_uop_rob_idx | _GEN_5422; // @[rob.scala 391:{59,59}]
  wire  _GEN_6718 = 5'h9 == io_lxcpt_bits_uop_rob_idx | _GEN_5423; // @[rob.scala 391:{59,59}]
  wire  _GEN_6719 = 5'ha == io_lxcpt_bits_uop_rob_idx | _GEN_5424; // @[rob.scala 391:{59,59}]
  wire  _GEN_6720 = 5'hb == io_lxcpt_bits_uop_rob_idx | _GEN_5425; // @[rob.scala 391:{59,59}]
  wire  _GEN_6721 = 5'hc == io_lxcpt_bits_uop_rob_idx | _GEN_5426; // @[rob.scala 391:{59,59}]
  wire  _GEN_6722 = 5'hd == io_lxcpt_bits_uop_rob_idx | _GEN_5427; // @[rob.scala 391:{59,59}]
  wire  _GEN_6723 = 5'he == io_lxcpt_bits_uop_rob_idx | _GEN_5428; // @[rob.scala 391:{59,59}]
  wire  _GEN_6724 = 5'hf == io_lxcpt_bits_uop_rob_idx | _GEN_5429; // @[rob.scala 391:{59,59}]
  wire  _GEN_6725 = 5'h10 == io_lxcpt_bits_uop_rob_idx | _GEN_5430; // @[rob.scala 391:{59,59}]
  wire  _GEN_6726 = 5'h11 == io_lxcpt_bits_uop_rob_idx | _GEN_5431; // @[rob.scala 391:{59,59}]
  wire  _GEN_6727 = 5'h12 == io_lxcpt_bits_uop_rob_idx | _GEN_5432; // @[rob.scala 391:{59,59}]
  wire  _GEN_6728 = 5'h13 == io_lxcpt_bits_uop_rob_idx | _GEN_5433; // @[rob.scala 391:{59,59}]
  wire  _GEN_6729 = 5'h14 == io_lxcpt_bits_uop_rob_idx | _GEN_5434; // @[rob.scala 391:{59,59}]
  wire  _GEN_6730 = 5'h15 == io_lxcpt_bits_uop_rob_idx | _GEN_5435; // @[rob.scala 391:{59,59}]
  wire  _GEN_6731 = 5'h16 == io_lxcpt_bits_uop_rob_idx | _GEN_5436; // @[rob.scala 391:{59,59}]
  wire  _GEN_6732 = 5'h17 == io_lxcpt_bits_uop_rob_idx | _GEN_5437; // @[rob.scala 391:{59,59}]
  wire  _GEN_6733 = 5'h18 == io_lxcpt_bits_uop_rob_idx | _GEN_5438; // @[rob.scala 391:{59,59}]
  wire  _GEN_6734 = 5'h19 == io_lxcpt_bits_uop_rob_idx | _GEN_5439; // @[rob.scala 391:{59,59}]
  wire  _GEN_6735 = 5'h1a == io_lxcpt_bits_uop_rob_idx | _GEN_5440; // @[rob.scala 391:{59,59}]
  wire  _GEN_6736 = 5'h1b == io_lxcpt_bits_uop_rob_idx | _GEN_5441; // @[rob.scala 391:{59,59}]
  wire  _GEN_6737 = 5'h1c == io_lxcpt_bits_uop_rob_idx | _GEN_5442; // @[rob.scala 391:{59,59}]
  wire  _GEN_6738 = 5'h1d == io_lxcpt_bits_uop_rob_idx | _GEN_5443; // @[rob.scala 391:{59,59}]
  wire  _GEN_6739 = 5'h1e == io_lxcpt_bits_uop_rob_idx | _GEN_5444; // @[rob.scala 391:{59,59}]
  wire  _GEN_6740 = 5'h1f == io_lxcpt_bits_uop_rob_idx | _GEN_5445; // @[rob.scala 391:{59,59}]
  wire  _T_65 = io_lxcpt_bits_cause != 5'h10; // @[rob.scala 392:33]
  wire  _GEN_6742 = 5'h1 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_1 : rob_unsafe_0; // @[rob.scala 394:{15,15}]
  wire  _GEN_6743 = 5'h2 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_2 : _GEN_6742; // @[rob.scala 394:{15,15}]
  wire  _GEN_6744 = 5'h3 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_3 : _GEN_6743; // @[rob.scala 394:{15,15}]
  wire  _GEN_6745 = 5'h4 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_4 : _GEN_6744; // @[rob.scala 394:{15,15}]
  wire  _GEN_6746 = 5'h5 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_5 : _GEN_6745; // @[rob.scala 394:{15,15}]
  wire  _GEN_6747 = 5'h6 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_6 : _GEN_6746; // @[rob.scala 394:{15,15}]
  wire  _GEN_6748 = 5'h7 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_7 : _GEN_6747; // @[rob.scala 394:{15,15}]
  wire  _GEN_6749 = 5'h8 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_8 : _GEN_6748; // @[rob.scala 394:{15,15}]
  wire  _GEN_6750 = 5'h9 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_9 : _GEN_6749; // @[rob.scala 394:{15,15}]
  wire  _GEN_6751 = 5'ha == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_10 : _GEN_6750; // @[rob.scala 394:{15,15}]
  wire  _GEN_6752 = 5'hb == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_11 : _GEN_6751; // @[rob.scala 394:{15,15}]
  wire  _GEN_6753 = 5'hc == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_12 : _GEN_6752; // @[rob.scala 394:{15,15}]
  wire  _GEN_6754 = 5'hd == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_13 : _GEN_6753; // @[rob.scala 394:{15,15}]
  wire  _GEN_6755 = 5'he == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_14 : _GEN_6754; // @[rob.scala 394:{15,15}]
  wire  _GEN_6756 = 5'hf == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_15 : _GEN_6755; // @[rob.scala 394:{15,15}]
  wire  _GEN_6757 = 5'h10 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_16 : _GEN_6756; // @[rob.scala 394:{15,15}]
  wire  _GEN_6758 = 5'h11 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_17 : _GEN_6757; // @[rob.scala 394:{15,15}]
  wire  _GEN_6759 = 5'h12 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_18 : _GEN_6758; // @[rob.scala 394:{15,15}]
  wire  _GEN_6760 = 5'h13 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_19 : _GEN_6759; // @[rob.scala 394:{15,15}]
  wire  _GEN_6761 = 5'h14 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_20 : _GEN_6760; // @[rob.scala 394:{15,15}]
  wire  _GEN_6762 = 5'h15 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_21 : _GEN_6761; // @[rob.scala 394:{15,15}]
  wire  _GEN_6763 = 5'h16 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_22 : _GEN_6762; // @[rob.scala 394:{15,15}]
  wire  _GEN_6764 = 5'h17 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_23 : _GEN_6763; // @[rob.scala 394:{15,15}]
  wire  _GEN_6765 = 5'h18 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_24 : _GEN_6764; // @[rob.scala 394:{15,15}]
  wire  _GEN_6766 = 5'h19 == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_25 : _GEN_6765; // @[rob.scala 394:{15,15}]
  wire  _GEN_6767 = 5'h1a == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_26 : _GEN_6766; // @[rob.scala 394:{15,15}]
  wire  _GEN_6768 = 5'h1b == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_27 : _GEN_6767; // @[rob.scala 394:{15,15}]
  wire  _GEN_6769 = 5'h1c == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_28 : _GEN_6768; // @[rob.scala 394:{15,15}]
  wire  _GEN_6770 = 5'h1d == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_29 : _GEN_6769; // @[rob.scala 394:{15,15}]
  wire  _GEN_6771 = 5'h1e == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_30 : _GEN_6770; // @[rob.scala 394:{15,15}]
  wire  _GEN_6772 = 5'h1f == io_lxcpt_bits_uop_rob_idx ? rob_unsafe_31 : _GEN_6771; // @[rob.scala 394:{15,15}]
  wire  _GEN_6773 = io_lxcpt_valid ? _GEN_6709 : _GEN_5414; // @[rob.scala 390:79]
  wire  _GEN_6774 = io_lxcpt_valid ? _GEN_6710 : _GEN_5415; // @[rob.scala 390:79]
  wire  _GEN_6775 = io_lxcpt_valid ? _GEN_6711 : _GEN_5416; // @[rob.scala 390:79]
  wire  _GEN_6776 = io_lxcpt_valid ? _GEN_6712 : _GEN_5417; // @[rob.scala 390:79]
  wire  _GEN_6777 = io_lxcpt_valid ? _GEN_6713 : _GEN_5418; // @[rob.scala 390:79]
  wire  _GEN_6778 = io_lxcpt_valid ? _GEN_6714 : _GEN_5419; // @[rob.scala 390:79]
  wire  _GEN_6779 = io_lxcpt_valid ? _GEN_6715 : _GEN_5420; // @[rob.scala 390:79]
  wire  _GEN_6780 = io_lxcpt_valid ? _GEN_6716 : _GEN_5421; // @[rob.scala 390:79]
  wire  _GEN_6781 = io_lxcpt_valid ? _GEN_6717 : _GEN_5422; // @[rob.scala 390:79]
  wire  _GEN_6782 = io_lxcpt_valid ? _GEN_6718 : _GEN_5423; // @[rob.scala 390:79]
  wire  _GEN_6783 = io_lxcpt_valid ? _GEN_6719 : _GEN_5424; // @[rob.scala 390:79]
  wire  _GEN_6784 = io_lxcpt_valid ? _GEN_6720 : _GEN_5425; // @[rob.scala 390:79]
  wire  _GEN_6785 = io_lxcpt_valid ? _GEN_6721 : _GEN_5426; // @[rob.scala 390:79]
  wire  _GEN_6786 = io_lxcpt_valid ? _GEN_6722 : _GEN_5427; // @[rob.scala 390:79]
  wire  _GEN_6787 = io_lxcpt_valid ? _GEN_6723 : _GEN_5428; // @[rob.scala 390:79]
  wire  _GEN_6788 = io_lxcpt_valid ? _GEN_6724 : _GEN_5429; // @[rob.scala 390:79]
  wire  _GEN_6789 = io_lxcpt_valid ? _GEN_6725 : _GEN_5430; // @[rob.scala 390:79]
  wire  _GEN_6790 = io_lxcpt_valid ? _GEN_6726 : _GEN_5431; // @[rob.scala 390:79]
  wire  _GEN_6791 = io_lxcpt_valid ? _GEN_6727 : _GEN_5432; // @[rob.scala 390:79]
  wire  _GEN_6792 = io_lxcpt_valid ? _GEN_6728 : _GEN_5433; // @[rob.scala 390:79]
  wire  _GEN_6793 = io_lxcpt_valid ? _GEN_6729 : _GEN_5434; // @[rob.scala 390:79]
  wire  _GEN_6794 = io_lxcpt_valid ? _GEN_6730 : _GEN_5435; // @[rob.scala 390:79]
  wire  _GEN_6795 = io_lxcpt_valid ? _GEN_6731 : _GEN_5436; // @[rob.scala 390:79]
  wire  _GEN_6796 = io_lxcpt_valid ? _GEN_6732 : _GEN_5437; // @[rob.scala 390:79]
  wire  _GEN_6797 = io_lxcpt_valid ? _GEN_6733 : _GEN_5438; // @[rob.scala 390:79]
  wire  _GEN_6798 = io_lxcpt_valid ? _GEN_6734 : _GEN_5439; // @[rob.scala 390:79]
  wire  _GEN_6799 = io_lxcpt_valid ? _GEN_6735 : _GEN_5440; // @[rob.scala 390:79]
  wire  _GEN_6800 = io_lxcpt_valid ? _GEN_6736 : _GEN_5441; // @[rob.scala 390:79]
  wire  _GEN_6801 = io_lxcpt_valid ? _GEN_6737 : _GEN_5442; // @[rob.scala 390:79]
  wire  _GEN_6802 = io_lxcpt_valid ? _GEN_6738 : _GEN_5443; // @[rob.scala 390:79]
  wire  _GEN_6803 = io_lxcpt_valid ? _GEN_6739 : _GEN_5444; // @[rob.scala 390:79]
  wire  _GEN_6804 = io_lxcpt_valid ? _GEN_6740 : _GEN_5445; // @[rob.scala 390:79]
  wire  _GEN_6902 = 5'h1 == com_idx ? rob_predicated_1 : rob_predicated_0; // @[rob.scala 410:{51,51}]
  wire  _GEN_6903 = 5'h2 == com_idx ? rob_predicated_2 : _GEN_6902; // @[rob.scala 410:{51,51}]
  wire  _GEN_6904 = 5'h3 == com_idx ? rob_predicated_3 : _GEN_6903; // @[rob.scala 410:{51,51}]
  wire  _GEN_6905 = 5'h4 == com_idx ? rob_predicated_4 : _GEN_6904; // @[rob.scala 410:{51,51}]
  wire  _GEN_6906 = 5'h5 == com_idx ? rob_predicated_5 : _GEN_6905; // @[rob.scala 410:{51,51}]
  wire  _GEN_6907 = 5'h6 == com_idx ? rob_predicated_6 : _GEN_6906; // @[rob.scala 410:{51,51}]
  wire  _GEN_6908 = 5'h7 == com_idx ? rob_predicated_7 : _GEN_6907; // @[rob.scala 410:{51,51}]
  wire  _GEN_6909 = 5'h8 == com_idx ? rob_predicated_8 : _GEN_6908; // @[rob.scala 410:{51,51}]
  wire  _GEN_6910 = 5'h9 == com_idx ? rob_predicated_9 : _GEN_6909; // @[rob.scala 410:{51,51}]
  wire  _GEN_6911 = 5'ha == com_idx ? rob_predicated_10 : _GEN_6910; // @[rob.scala 410:{51,51}]
  wire  _GEN_6912 = 5'hb == com_idx ? rob_predicated_11 : _GEN_6911; // @[rob.scala 410:{51,51}]
  wire  _GEN_6913 = 5'hc == com_idx ? rob_predicated_12 : _GEN_6912; // @[rob.scala 410:{51,51}]
  wire  _GEN_6914 = 5'hd == com_idx ? rob_predicated_13 : _GEN_6913; // @[rob.scala 410:{51,51}]
  wire  _GEN_6915 = 5'he == com_idx ? rob_predicated_14 : _GEN_6914; // @[rob.scala 410:{51,51}]
  wire  _GEN_6916 = 5'hf == com_idx ? rob_predicated_15 : _GEN_6915; // @[rob.scala 410:{51,51}]
  wire  _GEN_6917 = 5'h10 == com_idx ? rob_predicated_16 : _GEN_6916; // @[rob.scala 410:{51,51}]
  wire  _GEN_6918 = 5'h11 == com_idx ? rob_predicated_17 : _GEN_6917; // @[rob.scala 410:{51,51}]
  wire  _GEN_6919 = 5'h12 == com_idx ? rob_predicated_18 : _GEN_6918; // @[rob.scala 410:{51,51}]
  wire  _GEN_6920 = 5'h13 == com_idx ? rob_predicated_19 : _GEN_6919; // @[rob.scala 410:{51,51}]
  wire  _GEN_6921 = 5'h14 == com_idx ? rob_predicated_20 : _GEN_6920; // @[rob.scala 410:{51,51}]
  wire  _GEN_6922 = 5'h15 == com_idx ? rob_predicated_21 : _GEN_6921; // @[rob.scala 410:{51,51}]
  wire  _GEN_6923 = 5'h16 == com_idx ? rob_predicated_22 : _GEN_6922; // @[rob.scala 410:{51,51}]
  wire  _GEN_6924 = 5'h17 == com_idx ? rob_predicated_23 : _GEN_6923; // @[rob.scala 410:{51,51}]
  wire  _GEN_6925 = 5'h18 == com_idx ? rob_predicated_24 : _GEN_6924; // @[rob.scala 410:{51,51}]
  wire  _GEN_6926 = 5'h19 == com_idx ? rob_predicated_25 : _GEN_6925; // @[rob.scala 410:{51,51}]
  wire  _GEN_6927 = 5'h1a == com_idx ? rob_predicated_26 : _GEN_6926; // @[rob.scala 410:{51,51}]
  wire  _GEN_6928 = 5'h1b == com_idx ? rob_predicated_27 : _GEN_6927; // @[rob.scala 410:{51,51}]
  wire  _GEN_6929 = 5'h1c == com_idx ? rob_predicated_28 : _GEN_6928; // @[rob.scala 410:{51,51}]
  wire  _GEN_6930 = 5'h1d == com_idx ? rob_predicated_29 : _GEN_6929; // @[rob.scala 410:{51,51}]
  wire  _GEN_6931 = 5'h1e == com_idx ? rob_predicated_30 : _GEN_6930; // @[rob.scala 410:{51,51}]
  wire  _GEN_6932 = 5'h1f == com_idx ? rob_predicated_31 : _GEN_6931; // @[rob.scala 410:{51,51}]
  wire [1:0] _GEN_6934 = 5'h1 == com_idx ? rob_uop_1_debug_tsrc : rob_uop_0_debug_tsrc; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6935 = 5'h2 == com_idx ? rob_uop_2_debug_tsrc : _GEN_6934; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6936 = 5'h3 == com_idx ? rob_uop_3_debug_tsrc : _GEN_6935; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6937 = 5'h4 == com_idx ? rob_uop_4_debug_tsrc : _GEN_6936; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6938 = 5'h5 == com_idx ? rob_uop_5_debug_tsrc : _GEN_6937; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6939 = 5'h6 == com_idx ? rob_uop_6_debug_tsrc : _GEN_6938; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6940 = 5'h7 == com_idx ? rob_uop_7_debug_tsrc : _GEN_6939; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6941 = 5'h8 == com_idx ? rob_uop_8_debug_tsrc : _GEN_6940; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6942 = 5'h9 == com_idx ? rob_uop_9_debug_tsrc : _GEN_6941; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6943 = 5'ha == com_idx ? rob_uop_10_debug_tsrc : _GEN_6942; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6944 = 5'hb == com_idx ? rob_uop_11_debug_tsrc : _GEN_6943; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6945 = 5'hc == com_idx ? rob_uop_12_debug_tsrc : _GEN_6944; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6946 = 5'hd == com_idx ? rob_uop_13_debug_tsrc : _GEN_6945; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6947 = 5'he == com_idx ? rob_uop_14_debug_tsrc : _GEN_6946; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6948 = 5'hf == com_idx ? rob_uop_15_debug_tsrc : _GEN_6947; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6949 = 5'h10 == com_idx ? rob_uop_16_debug_tsrc : _GEN_6948; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6950 = 5'h11 == com_idx ? rob_uop_17_debug_tsrc : _GEN_6949; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6951 = 5'h12 == com_idx ? rob_uop_18_debug_tsrc : _GEN_6950; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6952 = 5'h13 == com_idx ? rob_uop_19_debug_tsrc : _GEN_6951; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6953 = 5'h14 == com_idx ? rob_uop_20_debug_tsrc : _GEN_6952; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6954 = 5'h15 == com_idx ? rob_uop_21_debug_tsrc : _GEN_6953; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6955 = 5'h16 == com_idx ? rob_uop_22_debug_tsrc : _GEN_6954; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6956 = 5'h17 == com_idx ? rob_uop_23_debug_tsrc : _GEN_6955; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6957 = 5'h18 == com_idx ? rob_uop_24_debug_tsrc : _GEN_6956; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6958 = 5'h19 == com_idx ? rob_uop_25_debug_tsrc : _GEN_6957; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6959 = 5'h1a == com_idx ? rob_uop_26_debug_tsrc : _GEN_6958; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6960 = 5'h1b == com_idx ? rob_uop_27_debug_tsrc : _GEN_6959; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6961 = 5'h1c == com_idx ? rob_uop_28_debug_tsrc : _GEN_6960; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6962 = 5'h1d == com_idx ? rob_uop_29_debug_tsrc : _GEN_6961; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6963 = 5'h1e == com_idx ? rob_uop_30_debug_tsrc : _GEN_6962; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6966 = 5'h1 == com_idx ? rob_uop_1_debug_fsrc : rob_uop_0_debug_fsrc; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6967 = 5'h2 == com_idx ? rob_uop_2_debug_fsrc : _GEN_6966; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6968 = 5'h3 == com_idx ? rob_uop_3_debug_fsrc : _GEN_6967; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6969 = 5'h4 == com_idx ? rob_uop_4_debug_fsrc : _GEN_6968; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6970 = 5'h5 == com_idx ? rob_uop_5_debug_fsrc : _GEN_6969; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6971 = 5'h6 == com_idx ? rob_uop_6_debug_fsrc : _GEN_6970; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6972 = 5'h7 == com_idx ? rob_uop_7_debug_fsrc : _GEN_6971; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6973 = 5'h8 == com_idx ? rob_uop_8_debug_fsrc : _GEN_6972; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6974 = 5'h9 == com_idx ? rob_uop_9_debug_fsrc : _GEN_6973; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6975 = 5'ha == com_idx ? rob_uop_10_debug_fsrc : _GEN_6974; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6976 = 5'hb == com_idx ? rob_uop_11_debug_fsrc : _GEN_6975; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6977 = 5'hc == com_idx ? rob_uop_12_debug_fsrc : _GEN_6976; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6978 = 5'hd == com_idx ? rob_uop_13_debug_fsrc : _GEN_6977; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6979 = 5'he == com_idx ? rob_uop_14_debug_fsrc : _GEN_6978; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6980 = 5'hf == com_idx ? rob_uop_15_debug_fsrc : _GEN_6979; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6981 = 5'h10 == com_idx ? rob_uop_16_debug_fsrc : _GEN_6980; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6982 = 5'h11 == com_idx ? rob_uop_17_debug_fsrc : _GEN_6981; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6983 = 5'h12 == com_idx ? rob_uop_18_debug_fsrc : _GEN_6982; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6984 = 5'h13 == com_idx ? rob_uop_19_debug_fsrc : _GEN_6983; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6985 = 5'h14 == com_idx ? rob_uop_20_debug_fsrc : _GEN_6984; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6986 = 5'h15 == com_idx ? rob_uop_21_debug_fsrc : _GEN_6985; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6987 = 5'h16 == com_idx ? rob_uop_22_debug_fsrc : _GEN_6986; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6988 = 5'h17 == com_idx ? rob_uop_23_debug_fsrc : _GEN_6987; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6989 = 5'h18 == com_idx ? rob_uop_24_debug_fsrc : _GEN_6988; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6990 = 5'h19 == com_idx ? rob_uop_25_debug_fsrc : _GEN_6989; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6991 = 5'h1a == com_idx ? rob_uop_26_debug_fsrc : _GEN_6990; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6992 = 5'h1b == com_idx ? rob_uop_27_debug_fsrc : _GEN_6991; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6993 = 5'h1c == com_idx ? rob_uop_28_debug_fsrc : _GEN_6992; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6994 = 5'h1d == com_idx ? rob_uop_29_debug_fsrc : _GEN_6993; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6995 = 5'h1e == com_idx ? rob_uop_30_debug_fsrc : _GEN_6994; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_6996 = 5'h1f == com_idx ? rob_uop_31_debug_fsrc : _GEN_6995; // @[rob.scala 411:{25,25}]
  wire  _GEN_6998 = 5'h1 == com_idx ? rob_uop_1_bp_xcpt_if : rob_uop_0_bp_xcpt_if; // @[rob.scala 411:{25,25}]
  wire  _GEN_6999 = 5'h2 == com_idx ? rob_uop_2_bp_xcpt_if : _GEN_6998; // @[rob.scala 411:{25,25}]
  wire  _GEN_7000 = 5'h3 == com_idx ? rob_uop_3_bp_xcpt_if : _GEN_6999; // @[rob.scala 411:{25,25}]
  wire  _GEN_7001 = 5'h4 == com_idx ? rob_uop_4_bp_xcpt_if : _GEN_7000; // @[rob.scala 411:{25,25}]
  wire  _GEN_7002 = 5'h5 == com_idx ? rob_uop_5_bp_xcpt_if : _GEN_7001; // @[rob.scala 411:{25,25}]
  wire  _GEN_7003 = 5'h6 == com_idx ? rob_uop_6_bp_xcpt_if : _GEN_7002; // @[rob.scala 411:{25,25}]
  wire  _GEN_7004 = 5'h7 == com_idx ? rob_uop_7_bp_xcpt_if : _GEN_7003; // @[rob.scala 411:{25,25}]
  wire  _GEN_7005 = 5'h8 == com_idx ? rob_uop_8_bp_xcpt_if : _GEN_7004; // @[rob.scala 411:{25,25}]
  wire  _GEN_7006 = 5'h9 == com_idx ? rob_uop_9_bp_xcpt_if : _GEN_7005; // @[rob.scala 411:{25,25}]
  wire  _GEN_7007 = 5'ha == com_idx ? rob_uop_10_bp_xcpt_if : _GEN_7006; // @[rob.scala 411:{25,25}]
  wire  _GEN_7008 = 5'hb == com_idx ? rob_uop_11_bp_xcpt_if : _GEN_7007; // @[rob.scala 411:{25,25}]
  wire  _GEN_7009 = 5'hc == com_idx ? rob_uop_12_bp_xcpt_if : _GEN_7008; // @[rob.scala 411:{25,25}]
  wire  _GEN_7010 = 5'hd == com_idx ? rob_uop_13_bp_xcpt_if : _GEN_7009; // @[rob.scala 411:{25,25}]
  wire  _GEN_7011 = 5'he == com_idx ? rob_uop_14_bp_xcpt_if : _GEN_7010; // @[rob.scala 411:{25,25}]
  wire  _GEN_7012 = 5'hf == com_idx ? rob_uop_15_bp_xcpt_if : _GEN_7011; // @[rob.scala 411:{25,25}]
  wire  _GEN_7013 = 5'h10 == com_idx ? rob_uop_16_bp_xcpt_if : _GEN_7012; // @[rob.scala 411:{25,25}]
  wire  _GEN_7014 = 5'h11 == com_idx ? rob_uop_17_bp_xcpt_if : _GEN_7013; // @[rob.scala 411:{25,25}]
  wire  _GEN_7015 = 5'h12 == com_idx ? rob_uop_18_bp_xcpt_if : _GEN_7014; // @[rob.scala 411:{25,25}]
  wire  _GEN_7016 = 5'h13 == com_idx ? rob_uop_19_bp_xcpt_if : _GEN_7015; // @[rob.scala 411:{25,25}]
  wire  _GEN_7017 = 5'h14 == com_idx ? rob_uop_20_bp_xcpt_if : _GEN_7016; // @[rob.scala 411:{25,25}]
  wire  _GEN_7018 = 5'h15 == com_idx ? rob_uop_21_bp_xcpt_if : _GEN_7017; // @[rob.scala 411:{25,25}]
  wire  _GEN_7019 = 5'h16 == com_idx ? rob_uop_22_bp_xcpt_if : _GEN_7018; // @[rob.scala 411:{25,25}]
  wire  _GEN_7020 = 5'h17 == com_idx ? rob_uop_23_bp_xcpt_if : _GEN_7019; // @[rob.scala 411:{25,25}]
  wire  _GEN_7021 = 5'h18 == com_idx ? rob_uop_24_bp_xcpt_if : _GEN_7020; // @[rob.scala 411:{25,25}]
  wire  _GEN_7022 = 5'h19 == com_idx ? rob_uop_25_bp_xcpt_if : _GEN_7021; // @[rob.scala 411:{25,25}]
  wire  _GEN_7023 = 5'h1a == com_idx ? rob_uop_26_bp_xcpt_if : _GEN_7022; // @[rob.scala 411:{25,25}]
  wire  _GEN_7024 = 5'h1b == com_idx ? rob_uop_27_bp_xcpt_if : _GEN_7023; // @[rob.scala 411:{25,25}]
  wire  _GEN_7025 = 5'h1c == com_idx ? rob_uop_28_bp_xcpt_if : _GEN_7024; // @[rob.scala 411:{25,25}]
  wire  _GEN_7026 = 5'h1d == com_idx ? rob_uop_29_bp_xcpt_if : _GEN_7025; // @[rob.scala 411:{25,25}]
  wire  _GEN_7027 = 5'h1e == com_idx ? rob_uop_30_bp_xcpt_if : _GEN_7026; // @[rob.scala 411:{25,25}]
  wire  _GEN_7030 = 5'h1 == com_idx ? rob_uop_1_bp_debug_if : rob_uop_0_bp_debug_if; // @[rob.scala 411:{25,25}]
  wire  _GEN_7031 = 5'h2 == com_idx ? rob_uop_2_bp_debug_if : _GEN_7030; // @[rob.scala 411:{25,25}]
  wire  _GEN_7032 = 5'h3 == com_idx ? rob_uop_3_bp_debug_if : _GEN_7031; // @[rob.scala 411:{25,25}]
  wire  _GEN_7033 = 5'h4 == com_idx ? rob_uop_4_bp_debug_if : _GEN_7032; // @[rob.scala 411:{25,25}]
  wire  _GEN_7034 = 5'h5 == com_idx ? rob_uop_5_bp_debug_if : _GEN_7033; // @[rob.scala 411:{25,25}]
  wire  _GEN_7035 = 5'h6 == com_idx ? rob_uop_6_bp_debug_if : _GEN_7034; // @[rob.scala 411:{25,25}]
  wire  _GEN_7036 = 5'h7 == com_idx ? rob_uop_7_bp_debug_if : _GEN_7035; // @[rob.scala 411:{25,25}]
  wire  _GEN_7037 = 5'h8 == com_idx ? rob_uop_8_bp_debug_if : _GEN_7036; // @[rob.scala 411:{25,25}]
  wire  _GEN_7038 = 5'h9 == com_idx ? rob_uop_9_bp_debug_if : _GEN_7037; // @[rob.scala 411:{25,25}]
  wire  _GEN_7039 = 5'ha == com_idx ? rob_uop_10_bp_debug_if : _GEN_7038; // @[rob.scala 411:{25,25}]
  wire  _GEN_7040 = 5'hb == com_idx ? rob_uop_11_bp_debug_if : _GEN_7039; // @[rob.scala 411:{25,25}]
  wire  _GEN_7041 = 5'hc == com_idx ? rob_uop_12_bp_debug_if : _GEN_7040; // @[rob.scala 411:{25,25}]
  wire  _GEN_7042 = 5'hd == com_idx ? rob_uop_13_bp_debug_if : _GEN_7041; // @[rob.scala 411:{25,25}]
  wire  _GEN_7043 = 5'he == com_idx ? rob_uop_14_bp_debug_if : _GEN_7042; // @[rob.scala 411:{25,25}]
  wire  _GEN_7044 = 5'hf == com_idx ? rob_uop_15_bp_debug_if : _GEN_7043; // @[rob.scala 411:{25,25}]
  wire  _GEN_7045 = 5'h10 == com_idx ? rob_uop_16_bp_debug_if : _GEN_7044; // @[rob.scala 411:{25,25}]
  wire  _GEN_7046 = 5'h11 == com_idx ? rob_uop_17_bp_debug_if : _GEN_7045; // @[rob.scala 411:{25,25}]
  wire  _GEN_7047 = 5'h12 == com_idx ? rob_uop_18_bp_debug_if : _GEN_7046; // @[rob.scala 411:{25,25}]
  wire  _GEN_7048 = 5'h13 == com_idx ? rob_uop_19_bp_debug_if : _GEN_7047; // @[rob.scala 411:{25,25}]
  wire  _GEN_7049 = 5'h14 == com_idx ? rob_uop_20_bp_debug_if : _GEN_7048; // @[rob.scala 411:{25,25}]
  wire  _GEN_7050 = 5'h15 == com_idx ? rob_uop_21_bp_debug_if : _GEN_7049; // @[rob.scala 411:{25,25}]
  wire  _GEN_7051 = 5'h16 == com_idx ? rob_uop_22_bp_debug_if : _GEN_7050; // @[rob.scala 411:{25,25}]
  wire  _GEN_7052 = 5'h17 == com_idx ? rob_uop_23_bp_debug_if : _GEN_7051; // @[rob.scala 411:{25,25}]
  wire  _GEN_7053 = 5'h18 == com_idx ? rob_uop_24_bp_debug_if : _GEN_7052; // @[rob.scala 411:{25,25}]
  wire  _GEN_7054 = 5'h19 == com_idx ? rob_uop_25_bp_debug_if : _GEN_7053; // @[rob.scala 411:{25,25}]
  wire  _GEN_7055 = 5'h1a == com_idx ? rob_uop_26_bp_debug_if : _GEN_7054; // @[rob.scala 411:{25,25}]
  wire  _GEN_7056 = 5'h1b == com_idx ? rob_uop_27_bp_debug_if : _GEN_7055; // @[rob.scala 411:{25,25}]
  wire  _GEN_7057 = 5'h1c == com_idx ? rob_uop_28_bp_debug_if : _GEN_7056; // @[rob.scala 411:{25,25}]
  wire  _GEN_7058 = 5'h1d == com_idx ? rob_uop_29_bp_debug_if : _GEN_7057; // @[rob.scala 411:{25,25}]
  wire  _GEN_7059 = 5'h1e == com_idx ? rob_uop_30_bp_debug_if : _GEN_7058; // @[rob.scala 411:{25,25}]
  wire  _GEN_7062 = 5'h1 == com_idx ? rob_uop_1_xcpt_ma_if : rob_uop_0_xcpt_ma_if; // @[rob.scala 411:{25,25}]
  wire  _GEN_7063 = 5'h2 == com_idx ? rob_uop_2_xcpt_ma_if : _GEN_7062; // @[rob.scala 411:{25,25}]
  wire  _GEN_7064 = 5'h3 == com_idx ? rob_uop_3_xcpt_ma_if : _GEN_7063; // @[rob.scala 411:{25,25}]
  wire  _GEN_7065 = 5'h4 == com_idx ? rob_uop_4_xcpt_ma_if : _GEN_7064; // @[rob.scala 411:{25,25}]
  wire  _GEN_7066 = 5'h5 == com_idx ? rob_uop_5_xcpt_ma_if : _GEN_7065; // @[rob.scala 411:{25,25}]
  wire  _GEN_7067 = 5'h6 == com_idx ? rob_uop_6_xcpt_ma_if : _GEN_7066; // @[rob.scala 411:{25,25}]
  wire  _GEN_7068 = 5'h7 == com_idx ? rob_uop_7_xcpt_ma_if : _GEN_7067; // @[rob.scala 411:{25,25}]
  wire  _GEN_7069 = 5'h8 == com_idx ? rob_uop_8_xcpt_ma_if : _GEN_7068; // @[rob.scala 411:{25,25}]
  wire  _GEN_7070 = 5'h9 == com_idx ? rob_uop_9_xcpt_ma_if : _GEN_7069; // @[rob.scala 411:{25,25}]
  wire  _GEN_7071 = 5'ha == com_idx ? rob_uop_10_xcpt_ma_if : _GEN_7070; // @[rob.scala 411:{25,25}]
  wire  _GEN_7072 = 5'hb == com_idx ? rob_uop_11_xcpt_ma_if : _GEN_7071; // @[rob.scala 411:{25,25}]
  wire  _GEN_7073 = 5'hc == com_idx ? rob_uop_12_xcpt_ma_if : _GEN_7072; // @[rob.scala 411:{25,25}]
  wire  _GEN_7074 = 5'hd == com_idx ? rob_uop_13_xcpt_ma_if : _GEN_7073; // @[rob.scala 411:{25,25}]
  wire  _GEN_7075 = 5'he == com_idx ? rob_uop_14_xcpt_ma_if : _GEN_7074; // @[rob.scala 411:{25,25}]
  wire  _GEN_7076 = 5'hf == com_idx ? rob_uop_15_xcpt_ma_if : _GEN_7075; // @[rob.scala 411:{25,25}]
  wire  _GEN_7077 = 5'h10 == com_idx ? rob_uop_16_xcpt_ma_if : _GEN_7076; // @[rob.scala 411:{25,25}]
  wire  _GEN_7078 = 5'h11 == com_idx ? rob_uop_17_xcpt_ma_if : _GEN_7077; // @[rob.scala 411:{25,25}]
  wire  _GEN_7079 = 5'h12 == com_idx ? rob_uop_18_xcpt_ma_if : _GEN_7078; // @[rob.scala 411:{25,25}]
  wire  _GEN_7080 = 5'h13 == com_idx ? rob_uop_19_xcpt_ma_if : _GEN_7079; // @[rob.scala 411:{25,25}]
  wire  _GEN_7081 = 5'h14 == com_idx ? rob_uop_20_xcpt_ma_if : _GEN_7080; // @[rob.scala 411:{25,25}]
  wire  _GEN_7082 = 5'h15 == com_idx ? rob_uop_21_xcpt_ma_if : _GEN_7081; // @[rob.scala 411:{25,25}]
  wire  _GEN_7083 = 5'h16 == com_idx ? rob_uop_22_xcpt_ma_if : _GEN_7082; // @[rob.scala 411:{25,25}]
  wire  _GEN_7084 = 5'h17 == com_idx ? rob_uop_23_xcpt_ma_if : _GEN_7083; // @[rob.scala 411:{25,25}]
  wire  _GEN_7085 = 5'h18 == com_idx ? rob_uop_24_xcpt_ma_if : _GEN_7084; // @[rob.scala 411:{25,25}]
  wire  _GEN_7086 = 5'h19 == com_idx ? rob_uop_25_xcpt_ma_if : _GEN_7085; // @[rob.scala 411:{25,25}]
  wire  _GEN_7087 = 5'h1a == com_idx ? rob_uop_26_xcpt_ma_if : _GEN_7086; // @[rob.scala 411:{25,25}]
  wire  _GEN_7088 = 5'h1b == com_idx ? rob_uop_27_xcpt_ma_if : _GEN_7087; // @[rob.scala 411:{25,25}]
  wire  _GEN_7089 = 5'h1c == com_idx ? rob_uop_28_xcpt_ma_if : _GEN_7088; // @[rob.scala 411:{25,25}]
  wire  _GEN_7090 = 5'h1d == com_idx ? rob_uop_29_xcpt_ma_if : _GEN_7089; // @[rob.scala 411:{25,25}]
  wire  _GEN_7091 = 5'h1e == com_idx ? rob_uop_30_xcpt_ma_if : _GEN_7090; // @[rob.scala 411:{25,25}]
  wire  _GEN_7094 = 5'h1 == com_idx ? rob_uop_1_xcpt_ae_if : rob_uop_0_xcpt_ae_if; // @[rob.scala 411:{25,25}]
  wire  _GEN_7095 = 5'h2 == com_idx ? rob_uop_2_xcpt_ae_if : _GEN_7094; // @[rob.scala 411:{25,25}]
  wire  _GEN_7096 = 5'h3 == com_idx ? rob_uop_3_xcpt_ae_if : _GEN_7095; // @[rob.scala 411:{25,25}]
  wire  _GEN_7097 = 5'h4 == com_idx ? rob_uop_4_xcpt_ae_if : _GEN_7096; // @[rob.scala 411:{25,25}]
  wire  _GEN_7098 = 5'h5 == com_idx ? rob_uop_5_xcpt_ae_if : _GEN_7097; // @[rob.scala 411:{25,25}]
  wire  _GEN_7099 = 5'h6 == com_idx ? rob_uop_6_xcpt_ae_if : _GEN_7098; // @[rob.scala 411:{25,25}]
  wire  _GEN_7100 = 5'h7 == com_idx ? rob_uop_7_xcpt_ae_if : _GEN_7099; // @[rob.scala 411:{25,25}]
  wire  _GEN_7101 = 5'h8 == com_idx ? rob_uop_8_xcpt_ae_if : _GEN_7100; // @[rob.scala 411:{25,25}]
  wire  _GEN_7102 = 5'h9 == com_idx ? rob_uop_9_xcpt_ae_if : _GEN_7101; // @[rob.scala 411:{25,25}]
  wire  _GEN_7103 = 5'ha == com_idx ? rob_uop_10_xcpt_ae_if : _GEN_7102; // @[rob.scala 411:{25,25}]
  wire  _GEN_7104 = 5'hb == com_idx ? rob_uop_11_xcpt_ae_if : _GEN_7103; // @[rob.scala 411:{25,25}]
  wire  _GEN_7105 = 5'hc == com_idx ? rob_uop_12_xcpt_ae_if : _GEN_7104; // @[rob.scala 411:{25,25}]
  wire  _GEN_7106 = 5'hd == com_idx ? rob_uop_13_xcpt_ae_if : _GEN_7105; // @[rob.scala 411:{25,25}]
  wire  _GEN_7107 = 5'he == com_idx ? rob_uop_14_xcpt_ae_if : _GEN_7106; // @[rob.scala 411:{25,25}]
  wire  _GEN_7108 = 5'hf == com_idx ? rob_uop_15_xcpt_ae_if : _GEN_7107; // @[rob.scala 411:{25,25}]
  wire  _GEN_7109 = 5'h10 == com_idx ? rob_uop_16_xcpt_ae_if : _GEN_7108; // @[rob.scala 411:{25,25}]
  wire  _GEN_7110 = 5'h11 == com_idx ? rob_uop_17_xcpt_ae_if : _GEN_7109; // @[rob.scala 411:{25,25}]
  wire  _GEN_7111 = 5'h12 == com_idx ? rob_uop_18_xcpt_ae_if : _GEN_7110; // @[rob.scala 411:{25,25}]
  wire  _GEN_7112 = 5'h13 == com_idx ? rob_uop_19_xcpt_ae_if : _GEN_7111; // @[rob.scala 411:{25,25}]
  wire  _GEN_7113 = 5'h14 == com_idx ? rob_uop_20_xcpt_ae_if : _GEN_7112; // @[rob.scala 411:{25,25}]
  wire  _GEN_7114 = 5'h15 == com_idx ? rob_uop_21_xcpt_ae_if : _GEN_7113; // @[rob.scala 411:{25,25}]
  wire  _GEN_7115 = 5'h16 == com_idx ? rob_uop_22_xcpt_ae_if : _GEN_7114; // @[rob.scala 411:{25,25}]
  wire  _GEN_7116 = 5'h17 == com_idx ? rob_uop_23_xcpt_ae_if : _GEN_7115; // @[rob.scala 411:{25,25}]
  wire  _GEN_7117 = 5'h18 == com_idx ? rob_uop_24_xcpt_ae_if : _GEN_7116; // @[rob.scala 411:{25,25}]
  wire  _GEN_7118 = 5'h19 == com_idx ? rob_uop_25_xcpt_ae_if : _GEN_7117; // @[rob.scala 411:{25,25}]
  wire  _GEN_7119 = 5'h1a == com_idx ? rob_uop_26_xcpt_ae_if : _GEN_7118; // @[rob.scala 411:{25,25}]
  wire  _GEN_7120 = 5'h1b == com_idx ? rob_uop_27_xcpt_ae_if : _GEN_7119; // @[rob.scala 411:{25,25}]
  wire  _GEN_7121 = 5'h1c == com_idx ? rob_uop_28_xcpt_ae_if : _GEN_7120; // @[rob.scala 411:{25,25}]
  wire  _GEN_7122 = 5'h1d == com_idx ? rob_uop_29_xcpt_ae_if : _GEN_7121; // @[rob.scala 411:{25,25}]
  wire  _GEN_7123 = 5'h1e == com_idx ? rob_uop_30_xcpt_ae_if : _GEN_7122; // @[rob.scala 411:{25,25}]
  wire  _GEN_7126 = 5'h1 == com_idx ? rob_uop_1_xcpt_pf_if : rob_uop_0_xcpt_pf_if; // @[rob.scala 411:{25,25}]
  wire  _GEN_7127 = 5'h2 == com_idx ? rob_uop_2_xcpt_pf_if : _GEN_7126; // @[rob.scala 411:{25,25}]
  wire  _GEN_7128 = 5'h3 == com_idx ? rob_uop_3_xcpt_pf_if : _GEN_7127; // @[rob.scala 411:{25,25}]
  wire  _GEN_7129 = 5'h4 == com_idx ? rob_uop_4_xcpt_pf_if : _GEN_7128; // @[rob.scala 411:{25,25}]
  wire  _GEN_7130 = 5'h5 == com_idx ? rob_uop_5_xcpt_pf_if : _GEN_7129; // @[rob.scala 411:{25,25}]
  wire  _GEN_7131 = 5'h6 == com_idx ? rob_uop_6_xcpt_pf_if : _GEN_7130; // @[rob.scala 411:{25,25}]
  wire  _GEN_7132 = 5'h7 == com_idx ? rob_uop_7_xcpt_pf_if : _GEN_7131; // @[rob.scala 411:{25,25}]
  wire  _GEN_7133 = 5'h8 == com_idx ? rob_uop_8_xcpt_pf_if : _GEN_7132; // @[rob.scala 411:{25,25}]
  wire  _GEN_7134 = 5'h9 == com_idx ? rob_uop_9_xcpt_pf_if : _GEN_7133; // @[rob.scala 411:{25,25}]
  wire  _GEN_7135 = 5'ha == com_idx ? rob_uop_10_xcpt_pf_if : _GEN_7134; // @[rob.scala 411:{25,25}]
  wire  _GEN_7136 = 5'hb == com_idx ? rob_uop_11_xcpt_pf_if : _GEN_7135; // @[rob.scala 411:{25,25}]
  wire  _GEN_7137 = 5'hc == com_idx ? rob_uop_12_xcpt_pf_if : _GEN_7136; // @[rob.scala 411:{25,25}]
  wire  _GEN_7138 = 5'hd == com_idx ? rob_uop_13_xcpt_pf_if : _GEN_7137; // @[rob.scala 411:{25,25}]
  wire  _GEN_7139 = 5'he == com_idx ? rob_uop_14_xcpt_pf_if : _GEN_7138; // @[rob.scala 411:{25,25}]
  wire  _GEN_7140 = 5'hf == com_idx ? rob_uop_15_xcpt_pf_if : _GEN_7139; // @[rob.scala 411:{25,25}]
  wire  _GEN_7141 = 5'h10 == com_idx ? rob_uop_16_xcpt_pf_if : _GEN_7140; // @[rob.scala 411:{25,25}]
  wire  _GEN_7142 = 5'h11 == com_idx ? rob_uop_17_xcpt_pf_if : _GEN_7141; // @[rob.scala 411:{25,25}]
  wire  _GEN_7143 = 5'h12 == com_idx ? rob_uop_18_xcpt_pf_if : _GEN_7142; // @[rob.scala 411:{25,25}]
  wire  _GEN_7144 = 5'h13 == com_idx ? rob_uop_19_xcpt_pf_if : _GEN_7143; // @[rob.scala 411:{25,25}]
  wire  _GEN_7145 = 5'h14 == com_idx ? rob_uop_20_xcpt_pf_if : _GEN_7144; // @[rob.scala 411:{25,25}]
  wire  _GEN_7146 = 5'h15 == com_idx ? rob_uop_21_xcpt_pf_if : _GEN_7145; // @[rob.scala 411:{25,25}]
  wire  _GEN_7147 = 5'h16 == com_idx ? rob_uop_22_xcpt_pf_if : _GEN_7146; // @[rob.scala 411:{25,25}]
  wire  _GEN_7148 = 5'h17 == com_idx ? rob_uop_23_xcpt_pf_if : _GEN_7147; // @[rob.scala 411:{25,25}]
  wire  _GEN_7149 = 5'h18 == com_idx ? rob_uop_24_xcpt_pf_if : _GEN_7148; // @[rob.scala 411:{25,25}]
  wire  _GEN_7150 = 5'h19 == com_idx ? rob_uop_25_xcpt_pf_if : _GEN_7149; // @[rob.scala 411:{25,25}]
  wire  _GEN_7151 = 5'h1a == com_idx ? rob_uop_26_xcpt_pf_if : _GEN_7150; // @[rob.scala 411:{25,25}]
  wire  _GEN_7152 = 5'h1b == com_idx ? rob_uop_27_xcpt_pf_if : _GEN_7151; // @[rob.scala 411:{25,25}]
  wire  _GEN_7153 = 5'h1c == com_idx ? rob_uop_28_xcpt_pf_if : _GEN_7152; // @[rob.scala 411:{25,25}]
  wire  _GEN_7154 = 5'h1d == com_idx ? rob_uop_29_xcpt_pf_if : _GEN_7153; // @[rob.scala 411:{25,25}]
  wire  _GEN_7155 = 5'h1e == com_idx ? rob_uop_30_xcpt_pf_if : _GEN_7154; // @[rob.scala 411:{25,25}]
  wire  _GEN_7158 = 5'h1 == com_idx ? rob_uop_1_fp_single : rob_uop_0_fp_single; // @[rob.scala 411:{25,25}]
  wire  _GEN_7159 = 5'h2 == com_idx ? rob_uop_2_fp_single : _GEN_7158; // @[rob.scala 411:{25,25}]
  wire  _GEN_7160 = 5'h3 == com_idx ? rob_uop_3_fp_single : _GEN_7159; // @[rob.scala 411:{25,25}]
  wire  _GEN_7161 = 5'h4 == com_idx ? rob_uop_4_fp_single : _GEN_7160; // @[rob.scala 411:{25,25}]
  wire  _GEN_7162 = 5'h5 == com_idx ? rob_uop_5_fp_single : _GEN_7161; // @[rob.scala 411:{25,25}]
  wire  _GEN_7163 = 5'h6 == com_idx ? rob_uop_6_fp_single : _GEN_7162; // @[rob.scala 411:{25,25}]
  wire  _GEN_7164 = 5'h7 == com_idx ? rob_uop_7_fp_single : _GEN_7163; // @[rob.scala 411:{25,25}]
  wire  _GEN_7165 = 5'h8 == com_idx ? rob_uop_8_fp_single : _GEN_7164; // @[rob.scala 411:{25,25}]
  wire  _GEN_7166 = 5'h9 == com_idx ? rob_uop_9_fp_single : _GEN_7165; // @[rob.scala 411:{25,25}]
  wire  _GEN_7167 = 5'ha == com_idx ? rob_uop_10_fp_single : _GEN_7166; // @[rob.scala 411:{25,25}]
  wire  _GEN_7168 = 5'hb == com_idx ? rob_uop_11_fp_single : _GEN_7167; // @[rob.scala 411:{25,25}]
  wire  _GEN_7169 = 5'hc == com_idx ? rob_uop_12_fp_single : _GEN_7168; // @[rob.scala 411:{25,25}]
  wire  _GEN_7170 = 5'hd == com_idx ? rob_uop_13_fp_single : _GEN_7169; // @[rob.scala 411:{25,25}]
  wire  _GEN_7171 = 5'he == com_idx ? rob_uop_14_fp_single : _GEN_7170; // @[rob.scala 411:{25,25}]
  wire  _GEN_7172 = 5'hf == com_idx ? rob_uop_15_fp_single : _GEN_7171; // @[rob.scala 411:{25,25}]
  wire  _GEN_7173 = 5'h10 == com_idx ? rob_uop_16_fp_single : _GEN_7172; // @[rob.scala 411:{25,25}]
  wire  _GEN_7174 = 5'h11 == com_idx ? rob_uop_17_fp_single : _GEN_7173; // @[rob.scala 411:{25,25}]
  wire  _GEN_7175 = 5'h12 == com_idx ? rob_uop_18_fp_single : _GEN_7174; // @[rob.scala 411:{25,25}]
  wire  _GEN_7176 = 5'h13 == com_idx ? rob_uop_19_fp_single : _GEN_7175; // @[rob.scala 411:{25,25}]
  wire  _GEN_7177 = 5'h14 == com_idx ? rob_uop_20_fp_single : _GEN_7176; // @[rob.scala 411:{25,25}]
  wire  _GEN_7178 = 5'h15 == com_idx ? rob_uop_21_fp_single : _GEN_7177; // @[rob.scala 411:{25,25}]
  wire  _GEN_7179 = 5'h16 == com_idx ? rob_uop_22_fp_single : _GEN_7178; // @[rob.scala 411:{25,25}]
  wire  _GEN_7180 = 5'h17 == com_idx ? rob_uop_23_fp_single : _GEN_7179; // @[rob.scala 411:{25,25}]
  wire  _GEN_7181 = 5'h18 == com_idx ? rob_uop_24_fp_single : _GEN_7180; // @[rob.scala 411:{25,25}]
  wire  _GEN_7182 = 5'h19 == com_idx ? rob_uop_25_fp_single : _GEN_7181; // @[rob.scala 411:{25,25}]
  wire  _GEN_7183 = 5'h1a == com_idx ? rob_uop_26_fp_single : _GEN_7182; // @[rob.scala 411:{25,25}]
  wire  _GEN_7184 = 5'h1b == com_idx ? rob_uop_27_fp_single : _GEN_7183; // @[rob.scala 411:{25,25}]
  wire  _GEN_7185 = 5'h1c == com_idx ? rob_uop_28_fp_single : _GEN_7184; // @[rob.scala 411:{25,25}]
  wire  _GEN_7186 = 5'h1d == com_idx ? rob_uop_29_fp_single : _GEN_7185; // @[rob.scala 411:{25,25}]
  wire  _GEN_7187 = 5'h1e == com_idx ? rob_uop_30_fp_single : _GEN_7186; // @[rob.scala 411:{25,25}]
  wire  _GEN_7190 = 5'h1 == com_idx ? rob_uop_1_fp_val : rob_uop_0_fp_val; // @[rob.scala 411:{25,25}]
  wire  _GEN_7191 = 5'h2 == com_idx ? rob_uop_2_fp_val : _GEN_7190; // @[rob.scala 411:{25,25}]
  wire  _GEN_7192 = 5'h3 == com_idx ? rob_uop_3_fp_val : _GEN_7191; // @[rob.scala 411:{25,25}]
  wire  _GEN_7193 = 5'h4 == com_idx ? rob_uop_4_fp_val : _GEN_7192; // @[rob.scala 411:{25,25}]
  wire  _GEN_7194 = 5'h5 == com_idx ? rob_uop_5_fp_val : _GEN_7193; // @[rob.scala 411:{25,25}]
  wire  _GEN_7195 = 5'h6 == com_idx ? rob_uop_6_fp_val : _GEN_7194; // @[rob.scala 411:{25,25}]
  wire  _GEN_7196 = 5'h7 == com_idx ? rob_uop_7_fp_val : _GEN_7195; // @[rob.scala 411:{25,25}]
  wire  _GEN_7197 = 5'h8 == com_idx ? rob_uop_8_fp_val : _GEN_7196; // @[rob.scala 411:{25,25}]
  wire  _GEN_7198 = 5'h9 == com_idx ? rob_uop_9_fp_val : _GEN_7197; // @[rob.scala 411:{25,25}]
  wire  _GEN_7199 = 5'ha == com_idx ? rob_uop_10_fp_val : _GEN_7198; // @[rob.scala 411:{25,25}]
  wire  _GEN_7200 = 5'hb == com_idx ? rob_uop_11_fp_val : _GEN_7199; // @[rob.scala 411:{25,25}]
  wire  _GEN_7201 = 5'hc == com_idx ? rob_uop_12_fp_val : _GEN_7200; // @[rob.scala 411:{25,25}]
  wire  _GEN_7202 = 5'hd == com_idx ? rob_uop_13_fp_val : _GEN_7201; // @[rob.scala 411:{25,25}]
  wire  _GEN_7203 = 5'he == com_idx ? rob_uop_14_fp_val : _GEN_7202; // @[rob.scala 411:{25,25}]
  wire  _GEN_7204 = 5'hf == com_idx ? rob_uop_15_fp_val : _GEN_7203; // @[rob.scala 411:{25,25}]
  wire  _GEN_7205 = 5'h10 == com_idx ? rob_uop_16_fp_val : _GEN_7204; // @[rob.scala 411:{25,25}]
  wire  _GEN_7206 = 5'h11 == com_idx ? rob_uop_17_fp_val : _GEN_7205; // @[rob.scala 411:{25,25}]
  wire  _GEN_7207 = 5'h12 == com_idx ? rob_uop_18_fp_val : _GEN_7206; // @[rob.scala 411:{25,25}]
  wire  _GEN_7208 = 5'h13 == com_idx ? rob_uop_19_fp_val : _GEN_7207; // @[rob.scala 411:{25,25}]
  wire  _GEN_7209 = 5'h14 == com_idx ? rob_uop_20_fp_val : _GEN_7208; // @[rob.scala 411:{25,25}]
  wire  _GEN_7210 = 5'h15 == com_idx ? rob_uop_21_fp_val : _GEN_7209; // @[rob.scala 411:{25,25}]
  wire  _GEN_7211 = 5'h16 == com_idx ? rob_uop_22_fp_val : _GEN_7210; // @[rob.scala 411:{25,25}]
  wire  _GEN_7212 = 5'h17 == com_idx ? rob_uop_23_fp_val : _GEN_7211; // @[rob.scala 411:{25,25}]
  wire  _GEN_7213 = 5'h18 == com_idx ? rob_uop_24_fp_val : _GEN_7212; // @[rob.scala 411:{25,25}]
  wire  _GEN_7214 = 5'h19 == com_idx ? rob_uop_25_fp_val : _GEN_7213; // @[rob.scala 411:{25,25}]
  wire  _GEN_7215 = 5'h1a == com_idx ? rob_uop_26_fp_val : _GEN_7214; // @[rob.scala 411:{25,25}]
  wire  _GEN_7216 = 5'h1b == com_idx ? rob_uop_27_fp_val : _GEN_7215; // @[rob.scala 411:{25,25}]
  wire  _GEN_7217 = 5'h1c == com_idx ? rob_uop_28_fp_val : _GEN_7216; // @[rob.scala 411:{25,25}]
  wire  _GEN_7218 = 5'h1d == com_idx ? rob_uop_29_fp_val : _GEN_7217; // @[rob.scala 411:{25,25}]
  wire  _GEN_7219 = 5'h1e == com_idx ? rob_uop_30_fp_val : _GEN_7218; // @[rob.scala 411:{25,25}]
  wire  _GEN_7222 = 5'h1 == com_idx ? rob_uop_1_frs3_en : rob_uop_0_frs3_en; // @[rob.scala 411:{25,25}]
  wire  _GEN_7223 = 5'h2 == com_idx ? rob_uop_2_frs3_en : _GEN_7222; // @[rob.scala 411:{25,25}]
  wire  _GEN_7224 = 5'h3 == com_idx ? rob_uop_3_frs3_en : _GEN_7223; // @[rob.scala 411:{25,25}]
  wire  _GEN_7225 = 5'h4 == com_idx ? rob_uop_4_frs3_en : _GEN_7224; // @[rob.scala 411:{25,25}]
  wire  _GEN_7226 = 5'h5 == com_idx ? rob_uop_5_frs3_en : _GEN_7225; // @[rob.scala 411:{25,25}]
  wire  _GEN_7227 = 5'h6 == com_idx ? rob_uop_6_frs3_en : _GEN_7226; // @[rob.scala 411:{25,25}]
  wire  _GEN_7228 = 5'h7 == com_idx ? rob_uop_7_frs3_en : _GEN_7227; // @[rob.scala 411:{25,25}]
  wire  _GEN_7229 = 5'h8 == com_idx ? rob_uop_8_frs3_en : _GEN_7228; // @[rob.scala 411:{25,25}]
  wire  _GEN_7230 = 5'h9 == com_idx ? rob_uop_9_frs3_en : _GEN_7229; // @[rob.scala 411:{25,25}]
  wire  _GEN_7231 = 5'ha == com_idx ? rob_uop_10_frs3_en : _GEN_7230; // @[rob.scala 411:{25,25}]
  wire  _GEN_7232 = 5'hb == com_idx ? rob_uop_11_frs3_en : _GEN_7231; // @[rob.scala 411:{25,25}]
  wire  _GEN_7233 = 5'hc == com_idx ? rob_uop_12_frs3_en : _GEN_7232; // @[rob.scala 411:{25,25}]
  wire  _GEN_7234 = 5'hd == com_idx ? rob_uop_13_frs3_en : _GEN_7233; // @[rob.scala 411:{25,25}]
  wire  _GEN_7235 = 5'he == com_idx ? rob_uop_14_frs3_en : _GEN_7234; // @[rob.scala 411:{25,25}]
  wire  _GEN_7236 = 5'hf == com_idx ? rob_uop_15_frs3_en : _GEN_7235; // @[rob.scala 411:{25,25}]
  wire  _GEN_7237 = 5'h10 == com_idx ? rob_uop_16_frs3_en : _GEN_7236; // @[rob.scala 411:{25,25}]
  wire  _GEN_7238 = 5'h11 == com_idx ? rob_uop_17_frs3_en : _GEN_7237; // @[rob.scala 411:{25,25}]
  wire  _GEN_7239 = 5'h12 == com_idx ? rob_uop_18_frs3_en : _GEN_7238; // @[rob.scala 411:{25,25}]
  wire  _GEN_7240 = 5'h13 == com_idx ? rob_uop_19_frs3_en : _GEN_7239; // @[rob.scala 411:{25,25}]
  wire  _GEN_7241 = 5'h14 == com_idx ? rob_uop_20_frs3_en : _GEN_7240; // @[rob.scala 411:{25,25}]
  wire  _GEN_7242 = 5'h15 == com_idx ? rob_uop_21_frs3_en : _GEN_7241; // @[rob.scala 411:{25,25}]
  wire  _GEN_7243 = 5'h16 == com_idx ? rob_uop_22_frs3_en : _GEN_7242; // @[rob.scala 411:{25,25}]
  wire  _GEN_7244 = 5'h17 == com_idx ? rob_uop_23_frs3_en : _GEN_7243; // @[rob.scala 411:{25,25}]
  wire  _GEN_7245 = 5'h18 == com_idx ? rob_uop_24_frs3_en : _GEN_7244; // @[rob.scala 411:{25,25}]
  wire  _GEN_7246 = 5'h19 == com_idx ? rob_uop_25_frs3_en : _GEN_7245; // @[rob.scala 411:{25,25}]
  wire  _GEN_7247 = 5'h1a == com_idx ? rob_uop_26_frs3_en : _GEN_7246; // @[rob.scala 411:{25,25}]
  wire  _GEN_7248 = 5'h1b == com_idx ? rob_uop_27_frs3_en : _GEN_7247; // @[rob.scala 411:{25,25}]
  wire  _GEN_7249 = 5'h1c == com_idx ? rob_uop_28_frs3_en : _GEN_7248; // @[rob.scala 411:{25,25}]
  wire  _GEN_7250 = 5'h1d == com_idx ? rob_uop_29_frs3_en : _GEN_7249; // @[rob.scala 411:{25,25}]
  wire  _GEN_7251 = 5'h1e == com_idx ? rob_uop_30_frs3_en : _GEN_7250; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7254 = 5'h1 == com_idx ? rob_uop_1_lrs2_rtype : rob_uop_0_lrs2_rtype; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7255 = 5'h2 == com_idx ? rob_uop_2_lrs2_rtype : _GEN_7254; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7256 = 5'h3 == com_idx ? rob_uop_3_lrs2_rtype : _GEN_7255; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7257 = 5'h4 == com_idx ? rob_uop_4_lrs2_rtype : _GEN_7256; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7258 = 5'h5 == com_idx ? rob_uop_5_lrs2_rtype : _GEN_7257; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7259 = 5'h6 == com_idx ? rob_uop_6_lrs2_rtype : _GEN_7258; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7260 = 5'h7 == com_idx ? rob_uop_7_lrs2_rtype : _GEN_7259; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7261 = 5'h8 == com_idx ? rob_uop_8_lrs2_rtype : _GEN_7260; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7262 = 5'h9 == com_idx ? rob_uop_9_lrs2_rtype : _GEN_7261; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7263 = 5'ha == com_idx ? rob_uop_10_lrs2_rtype : _GEN_7262; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7264 = 5'hb == com_idx ? rob_uop_11_lrs2_rtype : _GEN_7263; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7265 = 5'hc == com_idx ? rob_uop_12_lrs2_rtype : _GEN_7264; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7266 = 5'hd == com_idx ? rob_uop_13_lrs2_rtype : _GEN_7265; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7267 = 5'he == com_idx ? rob_uop_14_lrs2_rtype : _GEN_7266; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7268 = 5'hf == com_idx ? rob_uop_15_lrs2_rtype : _GEN_7267; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7269 = 5'h10 == com_idx ? rob_uop_16_lrs2_rtype : _GEN_7268; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7270 = 5'h11 == com_idx ? rob_uop_17_lrs2_rtype : _GEN_7269; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7271 = 5'h12 == com_idx ? rob_uop_18_lrs2_rtype : _GEN_7270; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7272 = 5'h13 == com_idx ? rob_uop_19_lrs2_rtype : _GEN_7271; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7273 = 5'h14 == com_idx ? rob_uop_20_lrs2_rtype : _GEN_7272; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7274 = 5'h15 == com_idx ? rob_uop_21_lrs2_rtype : _GEN_7273; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7275 = 5'h16 == com_idx ? rob_uop_22_lrs2_rtype : _GEN_7274; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7276 = 5'h17 == com_idx ? rob_uop_23_lrs2_rtype : _GEN_7275; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7277 = 5'h18 == com_idx ? rob_uop_24_lrs2_rtype : _GEN_7276; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7278 = 5'h19 == com_idx ? rob_uop_25_lrs2_rtype : _GEN_7277; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7279 = 5'h1a == com_idx ? rob_uop_26_lrs2_rtype : _GEN_7278; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7280 = 5'h1b == com_idx ? rob_uop_27_lrs2_rtype : _GEN_7279; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7281 = 5'h1c == com_idx ? rob_uop_28_lrs2_rtype : _GEN_7280; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7282 = 5'h1d == com_idx ? rob_uop_29_lrs2_rtype : _GEN_7281; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7283 = 5'h1e == com_idx ? rob_uop_30_lrs2_rtype : _GEN_7282; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7286 = 5'h1 == com_idx ? rob_uop_1_lrs1_rtype : rob_uop_0_lrs1_rtype; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7287 = 5'h2 == com_idx ? rob_uop_2_lrs1_rtype : _GEN_7286; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7288 = 5'h3 == com_idx ? rob_uop_3_lrs1_rtype : _GEN_7287; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7289 = 5'h4 == com_idx ? rob_uop_4_lrs1_rtype : _GEN_7288; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7290 = 5'h5 == com_idx ? rob_uop_5_lrs1_rtype : _GEN_7289; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7291 = 5'h6 == com_idx ? rob_uop_6_lrs1_rtype : _GEN_7290; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7292 = 5'h7 == com_idx ? rob_uop_7_lrs1_rtype : _GEN_7291; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7293 = 5'h8 == com_idx ? rob_uop_8_lrs1_rtype : _GEN_7292; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7294 = 5'h9 == com_idx ? rob_uop_9_lrs1_rtype : _GEN_7293; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7295 = 5'ha == com_idx ? rob_uop_10_lrs1_rtype : _GEN_7294; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7296 = 5'hb == com_idx ? rob_uop_11_lrs1_rtype : _GEN_7295; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7297 = 5'hc == com_idx ? rob_uop_12_lrs1_rtype : _GEN_7296; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7298 = 5'hd == com_idx ? rob_uop_13_lrs1_rtype : _GEN_7297; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7299 = 5'he == com_idx ? rob_uop_14_lrs1_rtype : _GEN_7298; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7300 = 5'hf == com_idx ? rob_uop_15_lrs1_rtype : _GEN_7299; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7301 = 5'h10 == com_idx ? rob_uop_16_lrs1_rtype : _GEN_7300; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7302 = 5'h11 == com_idx ? rob_uop_17_lrs1_rtype : _GEN_7301; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7303 = 5'h12 == com_idx ? rob_uop_18_lrs1_rtype : _GEN_7302; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7304 = 5'h13 == com_idx ? rob_uop_19_lrs1_rtype : _GEN_7303; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7305 = 5'h14 == com_idx ? rob_uop_20_lrs1_rtype : _GEN_7304; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7306 = 5'h15 == com_idx ? rob_uop_21_lrs1_rtype : _GEN_7305; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7307 = 5'h16 == com_idx ? rob_uop_22_lrs1_rtype : _GEN_7306; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7308 = 5'h17 == com_idx ? rob_uop_23_lrs1_rtype : _GEN_7307; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7309 = 5'h18 == com_idx ? rob_uop_24_lrs1_rtype : _GEN_7308; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7310 = 5'h19 == com_idx ? rob_uop_25_lrs1_rtype : _GEN_7309; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7311 = 5'h1a == com_idx ? rob_uop_26_lrs1_rtype : _GEN_7310; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7312 = 5'h1b == com_idx ? rob_uop_27_lrs1_rtype : _GEN_7311; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7313 = 5'h1c == com_idx ? rob_uop_28_lrs1_rtype : _GEN_7312; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7314 = 5'h1d == com_idx ? rob_uop_29_lrs1_rtype : _GEN_7313; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7315 = 5'h1e == com_idx ? rob_uop_30_lrs1_rtype : _GEN_7314; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7318 = 5'h1 == com_idx ? rob_uop_1_dst_rtype : rob_uop_0_dst_rtype; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7319 = 5'h2 == com_idx ? rob_uop_2_dst_rtype : _GEN_7318; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7320 = 5'h3 == com_idx ? rob_uop_3_dst_rtype : _GEN_7319; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7321 = 5'h4 == com_idx ? rob_uop_4_dst_rtype : _GEN_7320; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7322 = 5'h5 == com_idx ? rob_uop_5_dst_rtype : _GEN_7321; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7323 = 5'h6 == com_idx ? rob_uop_6_dst_rtype : _GEN_7322; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7324 = 5'h7 == com_idx ? rob_uop_7_dst_rtype : _GEN_7323; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7325 = 5'h8 == com_idx ? rob_uop_8_dst_rtype : _GEN_7324; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7326 = 5'h9 == com_idx ? rob_uop_9_dst_rtype : _GEN_7325; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7327 = 5'ha == com_idx ? rob_uop_10_dst_rtype : _GEN_7326; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7328 = 5'hb == com_idx ? rob_uop_11_dst_rtype : _GEN_7327; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7329 = 5'hc == com_idx ? rob_uop_12_dst_rtype : _GEN_7328; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7330 = 5'hd == com_idx ? rob_uop_13_dst_rtype : _GEN_7329; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7331 = 5'he == com_idx ? rob_uop_14_dst_rtype : _GEN_7330; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7332 = 5'hf == com_idx ? rob_uop_15_dst_rtype : _GEN_7331; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7333 = 5'h10 == com_idx ? rob_uop_16_dst_rtype : _GEN_7332; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7334 = 5'h11 == com_idx ? rob_uop_17_dst_rtype : _GEN_7333; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7335 = 5'h12 == com_idx ? rob_uop_18_dst_rtype : _GEN_7334; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7336 = 5'h13 == com_idx ? rob_uop_19_dst_rtype : _GEN_7335; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7337 = 5'h14 == com_idx ? rob_uop_20_dst_rtype : _GEN_7336; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7338 = 5'h15 == com_idx ? rob_uop_21_dst_rtype : _GEN_7337; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7339 = 5'h16 == com_idx ? rob_uop_22_dst_rtype : _GEN_7338; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7340 = 5'h17 == com_idx ? rob_uop_23_dst_rtype : _GEN_7339; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7341 = 5'h18 == com_idx ? rob_uop_24_dst_rtype : _GEN_7340; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7342 = 5'h19 == com_idx ? rob_uop_25_dst_rtype : _GEN_7341; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7343 = 5'h1a == com_idx ? rob_uop_26_dst_rtype : _GEN_7342; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7344 = 5'h1b == com_idx ? rob_uop_27_dst_rtype : _GEN_7343; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7345 = 5'h1c == com_idx ? rob_uop_28_dst_rtype : _GEN_7344; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7346 = 5'h1d == com_idx ? rob_uop_29_dst_rtype : _GEN_7345; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7347 = 5'h1e == com_idx ? rob_uop_30_dst_rtype : _GEN_7346; // @[rob.scala 411:{25,25}]
  wire  _GEN_7350 = 5'h1 == com_idx ? rob_uop_1_ldst_val : rob_uop_0_ldst_val; // @[rob.scala 411:{25,25}]
  wire  _GEN_7351 = 5'h2 == com_idx ? rob_uop_2_ldst_val : _GEN_7350; // @[rob.scala 411:{25,25}]
  wire  _GEN_7352 = 5'h3 == com_idx ? rob_uop_3_ldst_val : _GEN_7351; // @[rob.scala 411:{25,25}]
  wire  _GEN_7353 = 5'h4 == com_idx ? rob_uop_4_ldst_val : _GEN_7352; // @[rob.scala 411:{25,25}]
  wire  _GEN_7354 = 5'h5 == com_idx ? rob_uop_5_ldst_val : _GEN_7353; // @[rob.scala 411:{25,25}]
  wire  _GEN_7355 = 5'h6 == com_idx ? rob_uop_6_ldst_val : _GEN_7354; // @[rob.scala 411:{25,25}]
  wire  _GEN_7356 = 5'h7 == com_idx ? rob_uop_7_ldst_val : _GEN_7355; // @[rob.scala 411:{25,25}]
  wire  _GEN_7357 = 5'h8 == com_idx ? rob_uop_8_ldst_val : _GEN_7356; // @[rob.scala 411:{25,25}]
  wire  _GEN_7358 = 5'h9 == com_idx ? rob_uop_9_ldst_val : _GEN_7357; // @[rob.scala 411:{25,25}]
  wire  _GEN_7359 = 5'ha == com_idx ? rob_uop_10_ldst_val : _GEN_7358; // @[rob.scala 411:{25,25}]
  wire  _GEN_7360 = 5'hb == com_idx ? rob_uop_11_ldst_val : _GEN_7359; // @[rob.scala 411:{25,25}]
  wire  _GEN_7361 = 5'hc == com_idx ? rob_uop_12_ldst_val : _GEN_7360; // @[rob.scala 411:{25,25}]
  wire  _GEN_7362 = 5'hd == com_idx ? rob_uop_13_ldst_val : _GEN_7361; // @[rob.scala 411:{25,25}]
  wire  _GEN_7363 = 5'he == com_idx ? rob_uop_14_ldst_val : _GEN_7362; // @[rob.scala 411:{25,25}]
  wire  _GEN_7364 = 5'hf == com_idx ? rob_uop_15_ldst_val : _GEN_7363; // @[rob.scala 411:{25,25}]
  wire  _GEN_7365 = 5'h10 == com_idx ? rob_uop_16_ldst_val : _GEN_7364; // @[rob.scala 411:{25,25}]
  wire  _GEN_7366 = 5'h11 == com_idx ? rob_uop_17_ldst_val : _GEN_7365; // @[rob.scala 411:{25,25}]
  wire  _GEN_7367 = 5'h12 == com_idx ? rob_uop_18_ldst_val : _GEN_7366; // @[rob.scala 411:{25,25}]
  wire  _GEN_7368 = 5'h13 == com_idx ? rob_uop_19_ldst_val : _GEN_7367; // @[rob.scala 411:{25,25}]
  wire  _GEN_7369 = 5'h14 == com_idx ? rob_uop_20_ldst_val : _GEN_7368; // @[rob.scala 411:{25,25}]
  wire  _GEN_7370 = 5'h15 == com_idx ? rob_uop_21_ldst_val : _GEN_7369; // @[rob.scala 411:{25,25}]
  wire  _GEN_7371 = 5'h16 == com_idx ? rob_uop_22_ldst_val : _GEN_7370; // @[rob.scala 411:{25,25}]
  wire  _GEN_7372 = 5'h17 == com_idx ? rob_uop_23_ldst_val : _GEN_7371; // @[rob.scala 411:{25,25}]
  wire  _GEN_7373 = 5'h18 == com_idx ? rob_uop_24_ldst_val : _GEN_7372; // @[rob.scala 411:{25,25}]
  wire  _GEN_7374 = 5'h19 == com_idx ? rob_uop_25_ldst_val : _GEN_7373; // @[rob.scala 411:{25,25}]
  wire  _GEN_7375 = 5'h1a == com_idx ? rob_uop_26_ldst_val : _GEN_7374; // @[rob.scala 411:{25,25}]
  wire  _GEN_7376 = 5'h1b == com_idx ? rob_uop_27_ldst_val : _GEN_7375; // @[rob.scala 411:{25,25}]
  wire  _GEN_7377 = 5'h1c == com_idx ? rob_uop_28_ldst_val : _GEN_7376; // @[rob.scala 411:{25,25}]
  wire  _GEN_7378 = 5'h1d == com_idx ? rob_uop_29_ldst_val : _GEN_7377; // @[rob.scala 411:{25,25}]
  wire  _GEN_7379 = 5'h1e == com_idx ? rob_uop_30_ldst_val : _GEN_7378; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7382 = 5'h1 == com_idx ? rob_uop_1_lrs3 : rob_uop_0_lrs3; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7383 = 5'h2 == com_idx ? rob_uop_2_lrs3 : _GEN_7382; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7384 = 5'h3 == com_idx ? rob_uop_3_lrs3 : _GEN_7383; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7385 = 5'h4 == com_idx ? rob_uop_4_lrs3 : _GEN_7384; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7386 = 5'h5 == com_idx ? rob_uop_5_lrs3 : _GEN_7385; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7387 = 5'h6 == com_idx ? rob_uop_6_lrs3 : _GEN_7386; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7388 = 5'h7 == com_idx ? rob_uop_7_lrs3 : _GEN_7387; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7389 = 5'h8 == com_idx ? rob_uop_8_lrs3 : _GEN_7388; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7390 = 5'h9 == com_idx ? rob_uop_9_lrs3 : _GEN_7389; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7391 = 5'ha == com_idx ? rob_uop_10_lrs3 : _GEN_7390; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7392 = 5'hb == com_idx ? rob_uop_11_lrs3 : _GEN_7391; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7393 = 5'hc == com_idx ? rob_uop_12_lrs3 : _GEN_7392; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7394 = 5'hd == com_idx ? rob_uop_13_lrs3 : _GEN_7393; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7395 = 5'he == com_idx ? rob_uop_14_lrs3 : _GEN_7394; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7396 = 5'hf == com_idx ? rob_uop_15_lrs3 : _GEN_7395; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7397 = 5'h10 == com_idx ? rob_uop_16_lrs3 : _GEN_7396; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7398 = 5'h11 == com_idx ? rob_uop_17_lrs3 : _GEN_7397; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7399 = 5'h12 == com_idx ? rob_uop_18_lrs3 : _GEN_7398; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7400 = 5'h13 == com_idx ? rob_uop_19_lrs3 : _GEN_7399; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7401 = 5'h14 == com_idx ? rob_uop_20_lrs3 : _GEN_7400; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7402 = 5'h15 == com_idx ? rob_uop_21_lrs3 : _GEN_7401; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7403 = 5'h16 == com_idx ? rob_uop_22_lrs3 : _GEN_7402; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7404 = 5'h17 == com_idx ? rob_uop_23_lrs3 : _GEN_7403; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7405 = 5'h18 == com_idx ? rob_uop_24_lrs3 : _GEN_7404; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7406 = 5'h19 == com_idx ? rob_uop_25_lrs3 : _GEN_7405; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7407 = 5'h1a == com_idx ? rob_uop_26_lrs3 : _GEN_7406; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7408 = 5'h1b == com_idx ? rob_uop_27_lrs3 : _GEN_7407; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7409 = 5'h1c == com_idx ? rob_uop_28_lrs3 : _GEN_7408; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7410 = 5'h1d == com_idx ? rob_uop_29_lrs3 : _GEN_7409; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7411 = 5'h1e == com_idx ? rob_uop_30_lrs3 : _GEN_7410; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7414 = 5'h1 == com_idx ? rob_uop_1_lrs2 : rob_uop_0_lrs2; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7415 = 5'h2 == com_idx ? rob_uop_2_lrs2 : _GEN_7414; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7416 = 5'h3 == com_idx ? rob_uop_3_lrs2 : _GEN_7415; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7417 = 5'h4 == com_idx ? rob_uop_4_lrs2 : _GEN_7416; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7418 = 5'h5 == com_idx ? rob_uop_5_lrs2 : _GEN_7417; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7419 = 5'h6 == com_idx ? rob_uop_6_lrs2 : _GEN_7418; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7420 = 5'h7 == com_idx ? rob_uop_7_lrs2 : _GEN_7419; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7421 = 5'h8 == com_idx ? rob_uop_8_lrs2 : _GEN_7420; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7422 = 5'h9 == com_idx ? rob_uop_9_lrs2 : _GEN_7421; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7423 = 5'ha == com_idx ? rob_uop_10_lrs2 : _GEN_7422; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7424 = 5'hb == com_idx ? rob_uop_11_lrs2 : _GEN_7423; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7425 = 5'hc == com_idx ? rob_uop_12_lrs2 : _GEN_7424; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7426 = 5'hd == com_idx ? rob_uop_13_lrs2 : _GEN_7425; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7427 = 5'he == com_idx ? rob_uop_14_lrs2 : _GEN_7426; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7428 = 5'hf == com_idx ? rob_uop_15_lrs2 : _GEN_7427; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7429 = 5'h10 == com_idx ? rob_uop_16_lrs2 : _GEN_7428; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7430 = 5'h11 == com_idx ? rob_uop_17_lrs2 : _GEN_7429; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7431 = 5'h12 == com_idx ? rob_uop_18_lrs2 : _GEN_7430; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7432 = 5'h13 == com_idx ? rob_uop_19_lrs2 : _GEN_7431; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7433 = 5'h14 == com_idx ? rob_uop_20_lrs2 : _GEN_7432; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7434 = 5'h15 == com_idx ? rob_uop_21_lrs2 : _GEN_7433; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7435 = 5'h16 == com_idx ? rob_uop_22_lrs2 : _GEN_7434; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7436 = 5'h17 == com_idx ? rob_uop_23_lrs2 : _GEN_7435; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7437 = 5'h18 == com_idx ? rob_uop_24_lrs2 : _GEN_7436; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7438 = 5'h19 == com_idx ? rob_uop_25_lrs2 : _GEN_7437; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7439 = 5'h1a == com_idx ? rob_uop_26_lrs2 : _GEN_7438; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7440 = 5'h1b == com_idx ? rob_uop_27_lrs2 : _GEN_7439; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7441 = 5'h1c == com_idx ? rob_uop_28_lrs2 : _GEN_7440; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7442 = 5'h1d == com_idx ? rob_uop_29_lrs2 : _GEN_7441; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7443 = 5'h1e == com_idx ? rob_uop_30_lrs2 : _GEN_7442; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7446 = 5'h1 == com_idx ? rob_uop_1_lrs1 : rob_uop_0_lrs1; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7447 = 5'h2 == com_idx ? rob_uop_2_lrs1 : _GEN_7446; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7448 = 5'h3 == com_idx ? rob_uop_3_lrs1 : _GEN_7447; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7449 = 5'h4 == com_idx ? rob_uop_4_lrs1 : _GEN_7448; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7450 = 5'h5 == com_idx ? rob_uop_5_lrs1 : _GEN_7449; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7451 = 5'h6 == com_idx ? rob_uop_6_lrs1 : _GEN_7450; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7452 = 5'h7 == com_idx ? rob_uop_7_lrs1 : _GEN_7451; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7453 = 5'h8 == com_idx ? rob_uop_8_lrs1 : _GEN_7452; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7454 = 5'h9 == com_idx ? rob_uop_9_lrs1 : _GEN_7453; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7455 = 5'ha == com_idx ? rob_uop_10_lrs1 : _GEN_7454; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7456 = 5'hb == com_idx ? rob_uop_11_lrs1 : _GEN_7455; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7457 = 5'hc == com_idx ? rob_uop_12_lrs1 : _GEN_7456; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7458 = 5'hd == com_idx ? rob_uop_13_lrs1 : _GEN_7457; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7459 = 5'he == com_idx ? rob_uop_14_lrs1 : _GEN_7458; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7460 = 5'hf == com_idx ? rob_uop_15_lrs1 : _GEN_7459; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7461 = 5'h10 == com_idx ? rob_uop_16_lrs1 : _GEN_7460; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7462 = 5'h11 == com_idx ? rob_uop_17_lrs1 : _GEN_7461; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7463 = 5'h12 == com_idx ? rob_uop_18_lrs1 : _GEN_7462; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7464 = 5'h13 == com_idx ? rob_uop_19_lrs1 : _GEN_7463; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7465 = 5'h14 == com_idx ? rob_uop_20_lrs1 : _GEN_7464; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7466 = 5'h15 == com_idx ? rob_uop_21_lrs1 : _GEN_7465; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7467 = 5'h16 == com_idx ? rob_uop_22_lrs1 : _GEN_7466; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7468 = 5'h17 == com_idx ? rob_uop_23_lrs1 : _GEN_7467; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7469 = 5'h18 == com_idx ? rob_uop_24_lrs1 : _GEN_7468; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7470 = 5'h19 == com_idx ? rob_uop_25_lrs1 : _GEN_7469; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7471 = 5'h1a == com_idx ? rob_uop_26_lrs1 : _GEN_7470; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7472 = 5'h1b == com_idx ? rob_uop_27_lrs1 : _GEN_7471; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7473 = 5'h1c == com_idx ? rob_uop_28_lrs1 : _GEN_7472; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7474 = 5'h1d == com_idx ? rob_uop_29_lrs1 : _GEN_7473; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7475 = 5'h1e == com_idx ? rob_uop_30_lrs1 : _GEN_7474; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7478 = 5'h1 == com_idx ? rob_uop_1_ldst : rob_uop_0_ldst; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7479 = 5'h2 == com_idx ? rob_uop_2_ldst : _GEN_7478; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7480 = 5'h3 == com_idx ? rob_uop_3_ldst : _GEN_7479; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7481 = 5'h4 == com_idx ? rob_uop_4_ldst : _GEN_7480; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7482 = 5'h5 == com_idx ? rob_uop_5_ldst : _GEN_7481; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7483 = 5'h6 == com_idx ? rob_uop_6_ldst : _GEN_7482; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7484 = 5'h7 == com_idx ? rob_uop_7_ldst : _GEN_7483; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7485 = 5'h8 == com_idx ? rob_uop_8_ldst : _GEN_7484; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7486 = 5'h9 == com_idx ? rob_uop_9_ldst : _GEN_7485; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7487 = 5'ha == com_idx ? rob_uop_10_ldst : _GEN_7486; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7488 = 5'hb == com_idx ? rob_uop_11_ldst : _GEN_7487; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7489 = 5'hc == com_idx ? rob_uop_12_ldst : _GEN_7488; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7490 = 5'hd == com_idx ? rob_uop_13_ldst : _GEN_7489; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7491 = 5'he == com_idx ? rob_uop_14_ldst : _GEN_7490; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7492 = 5'hf == com_idx ? rob_uop_15_ldst : _GEN_7491; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7493 = 5'h10 == com_idx ? rob_uop_16_ldst : _GEN_7492; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7494 = 5'h11 == com_idx ? rob_uop_17_ldst : _GEN_7493; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7495 = 5'h12 == com_idx ? rob_uop_18_ldst : _GEN_7494; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7496 = 5'h13 == com_idx ? rob_uop_19_ldst : _GEN_7495; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7497 = 5'h14 == com_idx ? rob_uop_20_ldst : _GEN_7496; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7498 = 5'h15 == com_idx ? rob_uop_21_ldst : _GEN_7497; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7499 = 5'h16 == com_idx ? rob_uop_22_ldst : _GEN_7498; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7500 = 5'h17 == com_idx ? rob_uop_23_ldst : _GEN_7499; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7501 = 5'h18 == com_idx ? rob_uop_24_ldst : _GEN_7500; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7502 = 5'h19 == com_idx ? rob_uop_25_ldst : _GEN_7501; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7503 = 5'h1a == com_idx ? rob_uop_26_ldst : _GEN_7502; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7504 = 5'h1b == com_idx ? rob_uop_27_ldst : _GEN_7503; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7505 = 5'h1c == com_idx ? rob_uop_28_ldst : _GEN_7504; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7506 = 5'h1d == com_idx ? rob_uop_29_ldst : _GEN_7505; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7507 = 5'h1e == com_idx ? rob_uop_30_ldst : _GEN_7506; // @[rob.scala 411:{25,25}]
  wire  _GEN_7510 = 5'h1 == com_idx ? rob_uop_1_ldst_is_rs1 : rob_uop_0_ldst_is_rs1; // @[rob.scala 411:{25,25}]
  wire  _GEN_7511 = 5'h2 == com_idx ? rob_uop_2_ldst_is_rs1 : _GEN_7510; // @[rob.scala 411:{25,25}]
  wire  _GEN_7512 = 5'h3 == com_idx ? rob_uop_3_ldst_is_rs1 : _GEN_7511; // @[rob.scala 411:{25,25}]
  wire  _GEN_7513 = 5'h4 == com_idx ? rob_uop_4_ldst_is_rs1 : _GEN_7512; // @[rob.scala 411:{25,25}]
  wire  _GEN_7514 = 5'h5 == com_idx ? rob_uop_5_ldst_is_rs1 : _GEN_7513; // @[rob.scala 411:{25,25}]
  wire  _GEN_7515 = 5'h6 == com_idx ? rob_uop_6_ldst_is_rs1 : _GEN_7514; // @[rob.scala 411:{25,25}]
  wire  _GEN_7516 = 5'h7 == com_idx ? rob_uop_7_ldst_is_rs1 : _GEN_7515; // @[rob.scala 411:{25,25}]
  wire  _GEN_7517 = 5'h8 == com_idx ? rob_uop_8_ldst_is_rs1 : _GEN_7516; // @[rob.scala 411:{25,25}]
  wire  _GEN_7518 = 5'h9 == com_idx ? rob_uop_9_ldst_is_rs1 : _GEN_7517; // @[rob.scala 411:{25,25}]
  wire  _GEN_7519 = 5'ha == com_idx ? rob_uop_10_ldst_is_rs1 : _GEN_7518; // @[rob.scala 411:{25,25}]
  wire  _GEN_7520 = 5'hb == com_idx ? rob_uop_11_ldst_is_rs1 : _GEN_7519; // @[rob.scala 411:{25,25}]
  wire  _GEN_7521 = 5'hc == com_idx ? rob_uop_12_ldst_is_rs1 : _GEN_7520; // @[rob.scala 411:{25,25}]
  wire  _GEN_7522 = 5'hd == com_idx ? rob_uop_13_ldst_is_rs1 : _GEN_7521; // @[rob.scala 411:{25,25}]
  wire  _GEN_7523 = 5'he == com_idx ? rob_uop_14_ldst_is_rs1 : _GEN_7522; // @[rob.scala 411:{25,25}]
  wire  _GEN_7524 = 5'hf == com_idx ? rob_uop_15_ldst_is_rs1 : _GEN_7523; // @[rob.scala 411:{25,25}]
  wire  _GEN_7525 = 5'h10 == com_idx ? rob_uop_16_ldst_is_rs1 : _GEN_7524; // @[rob.scala 411:{25,25}]
  wire  _GEN_7526 = 5'h11 == com_idx ? rob_uop_17_ldst_is_rs1 : _GEN_7525; // @[rob.scala 411:{25,25}]
  wire  _GEN_7527 = 5'h12 == com_idx ? rob_uop_18_ldst_is_rs1 : _GEN_7526; // @[rob.scala 411:{25,25}]
  wire  _GEN_7528 = 5'h13 == com_idx ? rob_uop_19_ldst_is_rs1 : _GEN_7527; // @[rob.scala 411:{25,25}]
  wire  _GEN_7529 = 5'h14 == com_idx ? rob_uop_20_ldst_is_rs1 : _GEN_7528; // @[rob.scala 411:{25,25}]
  wire  _GEN_7530 = 5'h15 == com_idx ? rob_uop_21_ldst_is_rs1 : _GEN_7529; // @[rob.scala 411:{25,25}]
  wire  _GEN_7531 = 5'h16 == com_idx ? rob_uop_22_ldst_is_rs1 : _GEN_7530; // @[rob.scala 411:{25,25}]
  wire  _GEN_7532 = 5'h17 == com_idx ? rob_uop_23_ldst_is_rs1 : _GEN_7531; // @[rob.scala 411:{25,25}]
  wire  _GEN_7533 = 5'h18 == com_idx ? rob_uop_24_ldst_is_rs1 : _GEN_7532; // @[rob.scala 411:{25,25}]
  wire  _GEN_7534 = 5'h19 == com_idx ? rob_uop_25_ldst_is_rs1 : _GEN_7533; // @[rob.scala 411:{25,25}]
  wire  _GEN_7535 = 5'h1a == com_idx ? rob_uop_26_ldst_is_rs1 : _GEN_7534; // @[rob.scala 411:{25,25}]
  wire  _GEN_7536 = 5'h1b == com_idx ? rob_uop_27_ldst_is_rs1 : _GEN_7535; // @[rob.scala 411:{25,25}]
  wire  _GEN_7537 = 5'h1c == com_idx ? rob_uop_28_ldst_is_rs1 : _GEN_7536; // @[rob.scala 411:{25,25}]
  wire  _GEN_7538 = 5'h1d == com_idx ? rob_uop_29_ldst_is_rs1 : _GEN_7537; // @[rob.scala 411:{25,25}]
  wire  _GEN_7539 = 5'h1e == com_idx ? rob_uop_30_ldst_is_rs1 : _GEN_7538; // @[rob.scala 411:{25,25}]
  wire  _GEN_7542 = 5'h1 == com_idx ? rob_uop_1_flush_on_commit : rob_uop_0_flush_on_commit; // @[rob.scala 411:{25,25}]
  wire  _GEN_7543 = 5'h2 == com_idx ? rob_uop_2_flush_on_commit : _GEN_7542; // @[rob.scala 411:{25,25}]
  wire  _GEN_7544 = 5'h3 == com_idx ? rob_uop_3_flush_on_commit : _GEN_7543; // @[rob.scala 411:{25,25}]
  wire  _GEN_7545 = 5'h4 == com_idx ? rob_uop_4_flush_on_commit : _GEN_7544; // @[rob.scala 411:{25,25}]
  wire  _GEN_7546 = 5'h5 == com_idx ? rob_uop_5_flush_on_commit : _GEN_7545; // @[rob.scala 411:{25,25}]
  wire  _GEN_7547 = 5'h6 == com_idx ? rob_uop_6_flush_on_commit : _GEN_7546; // @[rob.scala 411:{25,25}]
  wire  _GEN_7548 = 5'h7 == com_idx ? rob_uop_7_flush_on_commit : _GEN_7547; // @[rob.scala 411:{25,25}]
  wire  _GEN_7549 = 5'h8 == com_idx ? rob_uop_8_flush_on_commit : _GEN_7548; // @[rob.scala 411:{25,25}]
  wire  _GEN_7550 = 5'h9 == com_idx ? rob_uop_9_flush_on_commit : _GEN_7549; // @[rob.scala 411:{25,25}]
  wire  _GEN_7551 = 5'ha == com_idx ? rob_uop_10_flush_on_commit : _GEN_7550; // @[rob.scala 411:{25,25}]
  wire  _GEN_7552 = 5'hb == com_idx ? rob_uop_11_flush_on_commit : _GEN_7551; // @[rob.scala 411:{25,25}]
  wire  _GEN_7553 = 5'hc == com_idx ? rob_uop_12_flush_on_commit : _GEN_7552; // @[rob.scala 411:{25,25}]
  wire  _GEN_7554 = 5'hd == com_idx ? rob_uop_13_flush_on_commit : _GEN_7553; // @[rob.scala 411:{25,25}]
  wire  _GEN_7555 = 5'he == com_idx ? rob_uop_14_flush_on_commit : _GEN_7554; // @[rob.scala 411:{25,25}]
  wire  _GEN_7556 = 5'hf == com_idx ? rob_uop_15_flush_on_commit : _GEN_7555; // @[rob.scala 411:{25,25}]
  wire  _GEN_7557 = 5'h10 == com_idx ? rob_uop_16_flush_on_commit : _GEN_7556; // @[rob.scala 411:{25,25}]
  wire  _GEN_7558 = 5'h11 == com_idx ? rob_uop_17_flush_on_commit : _GEN_7557; // @[rob.scala 411:{25,25}]
  wire  _GEN_7559 = 5'h12 == com_idx ? rob_uop_18_flush_on_commit : _GEN_7558; // @[rob.scala 411:{25,25}]
  wire  _GEN_7560 = 5'h13 == com_idx ? rob_uop_19_flush_on_commit : _GEN_7559; // @[rob.scala 411:{25,25}]
  wire  _GEN_7561 = 5'h14 == com_idx ? rob_uop_20_flush_on_commit : _GEN_7560; // @[rob.scala 411:{25,25}]
  wire  _GEN_7562 = 5'h15 == com_idx ? rob_uop_21_flush_on_commit : _GEN_7561; // @[rob.scala 411:{25,25}]
  wire  _GEN_7563 = 5'h16 == com_idx ? rob_uop_22_flush_on_commit : _GEN_7562; // @[rob.scala 411:{25,25}]
  wire  _GEN_7564 = 5'h17 == com_idx ? rob_uop_23_flush_on_commit : _GEN_7563; // @[rob.scala 411:{25,25}]
  wire  _GEN_7565 = 5'h18 == com_idx ? rob_uop_24_flush_on_commit : _GEN_7564; // @[rob.scala 411:{25,25}]
  wire  _GEN_7566 = 5'h19 == com_idx ? rob_uop_25_flush_on_commit : _GEN_7565; // @[rob.scala 411:{25,25}]
  wire  _GEN_7567 = 5'h1a == com_idx ? rob_uop_26_flush_on_commit : _GEN_7566; // @[rob.scala 411:{25,25}]
  wire  _GEN_7568 = 5'h1b == com_idx ? rob_uop_27_flush_on_commit : _GEN_7567; // @[rob.scala 411:{25,25}]
  wire  _GEN_7569 = 5'h1c == com_idx ? rob_uop_28_flush_on_commit : _GEN_7568; // @[rob.scala 411:{25,25}]
  wire  _GEN_7570 = 5'h1d == com_idx ? rob_uop_29_flush_on_commit : _GEN_7569; // @[rob.scala 411:{25,25}]
  wire  _GEN_7571 = 5'h1e == com_idx ? rob_uop_30_flush_on_commit : _GEN_7570; // @[rob.scala 411:{25,25}]
  wire  _GEN_7574 = 5'h1 == com_idx ? rob_uop_1_is_unique : rob_uop_0_is_unique; // @[rob.scala 411:{25,25}]
  wire  _GEN_7575 = 5'h2 == com_idx ? rob_uop_2_is_unique : _GEN_7574; // @[rob.scala 411:{25,25}]
  wire  _GEN_7576 = 5'h3 == com_idx ? rob_uop_3_is_unique : _GEN_7575; // @[rob.scala 411:{25,25}]
  wire  _GEN_7577 = 5'h4 == com_idx ? rob_uop_4_is_unique : _GEN_7576; // @[rob.scala 411:{25,25}]
  wire  _GEN_7578 = 5'h5 == com_idx ? rob_uop_5_is_unique : _GEN_7577; // @[rob.scala 411:{25,25}]
  wire  _GEN_7579 = 5'h6 == com_idx ? rob_uop_6_is_unique : _GEN_7578; // @[rob.scala 411:{25,25}]
  wire  _GEN_7580 = 5'h7 == com_idx ? rob_uop_7_is_unique : _GEN_7579; // @[rob.scala 411:{25,25}]
  wire  _GEN_7581 = 5'h8 == com_idx ? rob_uop_8_is_unique : _GEN_7580; // @[rob.scala 411:{25,25}]
  wire  _GEN_7582 = 5'h9 == com_idx ? rob_uop_9_is_unique : _GEN_7581; // @[rob.scala 411:{25,25}]
  wire  _GEN_7583 = 5'ha == com_idx ? rob_uop_10_is_unique : _GEN_7582; // @[rob.scala 411:{25,25}]
  wire  _GEN_7584 = 5'hb == com_idx ? rob_uop_11_is_unique : _GEN_7583; // @[rob.scala 411:{25,25}]
  wire  _GEN_7585 = 5'hc == com_idx ? rob_uop_12_is_unique : _GEN_7584; // @[rob.scala 411:{25,25}]
  wire  _GEN_7586 = 5'hd == com_idx ? rob_uop_13_is_unique : _GEN_7585; // @[rob.scala 411:{25,25}]
  wire  _GEN_7587 = 5'he == com_idx ? rob_uop_14_is_unique : _GEN_7586; // @[rob.scala 411:{25,25}]
  wire  _GEN_7588 = 5'hf == com_idx ? rob_uop_15_is_unique : _GEN_7587; // @[rob.scala 411:{25,25}]
  wire  _GEN_7589 = 5'h10 == com_idx ? rob_uop_16_is_unique : _GEN_7588; // @[rob.scala 411:{25,25}]
  wire  _GEN_7590 = 5'h11 == com_idx ? rob_uop_17_is_unique : _GEN_7589; // @[rob.scala 411:{25,25}]
  wire  _GEN_7591 = 5'h12 == com_idx ? rob_uop_18_is_unique : _GEN_7590; // @[rob.scala 411:{25,25}]
  wire  _GEN_7592 = 5'h13 == com_idx ? rob_uop_19_is_unique : _GEN_7591; // @[rob.scala 411:{25,25}]
  wire  _GEN_7593 = 5'h14 == com_idx ? rob_uop_20_is_unique : _GEN_7592; // @[rob.scala 411:{25,25}]
  wire  _GEN_7594 = 5'h15 == com_idx ? rob_uop_21_is_unique : _GEN_7593; // @[rob.scala 411:{25,25}]
  wire  _GEN_7595 = 5'h16 == com_idx ? rob_uop_22_is_unique : _GEN_7594; // @[rob.scala 411:{25,25}]
  wire  _GEN_7596 = 5'h17 == com_idx ? rob_uop_23_is_unique : _GEN_7595; // @[rob.scala 411:{25,25}]
  wire  _GEN_7597 = 5'h18 == com_idx ? rob_uop_24_is_unique : _GEN_7596; // @[rob.scala 411:{25,25}]
  wire  _GEN_7598 = 5'h19 == com_idx ? rob_uop_25_is_unique : _GEN_7597; // @[rob.scala 411:{25,25}]
  wire  _GEN_7599 = 5'h1a == com_idx ? rob_uop_26_is_unique : _GEN_7598; // @[rob.scala 411:{25,25}]
  wire  _GEN_7600 = 5'h1b == com_idx ? rob_uop_27_is_unique : _GEN_7599; // @[rob.scala 411:{25,25}]
  wire  _GEN_7601 = 5'h1c == com_idx ? rob_uop_28_is_unique : _GEN_7600; // @[rob.scala 411:{25,25}]
  wire  _GEN_7602 = 5'h1d == com_idx ? rob_uop_29_is_unique : _GEN_7601; // @[rob.scala 411:{25,25}]
  wire  _GEN_7603 = 5'h1e == com_idx ? rob_uop_30_is_unique : _GEN_7602; // @[rob.scala 411:{25,25}]
  wire  _GEN_7606 = 5'h1 == com_idx ? rob_uop_1_is_sys_pc2epc : rob_uop_0_is_sys_pc2epc; // @[rob.scala 411:{25,25}]
  wire  _GEN_7607 = 5'h2 == com_idx ? rob_uop_2_is_sys_pc2epc : _GEN_7606; // @[rob.scala 411:{25,25}]
  wire  _GEN_7608 = 5'h3 == com_idx ? rob_uop_3_is_sys_pc2epc : _GEN_7607; // @[rob.scala 411:{25,25}]
  wire  _GEN_7609 = 5'h4 == com_idx ? rob_uop_4_is_sys_pc2epc : _GEN_7608; // @[rob.scala 411:{25,25}]
  wire  _GEN_7610 = 5'h5 == com_idx ? rob_uop_5_is_sys_pc2epc : _GEN_7609; // @[rob.scala 411:{25,25}]
  wire  _GEN_7611 = 5'h6 == com_idx ? rob_uop_6_is_sys_pc2epc : _GEN_7610; // @[rob.scala 411:{25,25}]
  wire  _GEN_7612 = 5'h7 == com_idx ? rob_uop_7_is_sys_pc2epc : _GEN_7611; // @[rob.scala 411:{25,25}]
  wire  _GEN_7613 = 5'h8 == com_idx ? rob_uop_8_is_sys_pc2epc : _GEN_7612; // @[rob.scala 411:{25,25}]
  wire  _GEN_7614 = 5'h9 == com_idx ? rob_uop_9_is_sys_pc2epc : _GEN_7613; // @[rob.scala 411:{25,25}]
  wire  _GEN_7615 = 5'ha == com_idx ? rob_uop_10_is_sys_pc2epc : _GEN_7614; // @[rob.scala 411:{25,25}]
  wire  _GEN_7616 = 5'hb == com_idx ? rob_uop_11_is_sys_pc2epc : _GEN_7615; // @[rob.scala 411:{25,25}]
  wire  _GEN_7617 = 5'hc == com_idx ? rob_uop_12_is_sys_pc2epc : _GEN_7616; // @[rob.scala 411:{25,25}]
  wire  _GEN_7618 = 5'hd == com_idx ? rob_uop_13_is_sys_pc2epc : _GEN_7617; // @[rob.scala 411:{25,25}]
  wire  _GEN_7619 = 5'he == com_idx ? rob_uop_14_is_sys_pc2epc : _GEN_7618; // @[rob.scala 411:{25,25}]
  wire  _GEN_7620 = 5'hf == com_idx ? rob_uop_15_is_sys_pc2epc : _GEN_7619; // @[rob.scala 411:{25,25}]
  wire  _GEN_7621 = 5'h10 == com_idx ? rob_uop_16_is_sys_pc2epc : _GEN_7620; // @[rob.scala 411:{25,25}]
  wire  _GEN_7622 = 5'h11 == com_idx ? rob_uop_17_is_sys_pc2epc : _GEN_7621; // @[rob.scala 411:{25,25}]
  wire  _GEN_7623 = 5'h12 == com_idx ? rob_uop_18_is_sys_pc2epc : _GEN_7622; // @[rob.scala 411:{25,25}]
  wire  _GEN_7624 = 5'h13 == com_idx ? rob_uop_19_is_sys_pc2epc : _GEN_7623; // @[rob.scala 411:{25,25}]
  wire  _GEN_7625 = 5'h14 == com_idx ? rob_uop_20_is_sys_pc2epc : _GEN_7624; // @[rob.scala 411:{25,25}]
  wire  _GEN_7626 = 5'h15 == com_idx ? rob_uop_21_is_sys_pc2epc : _GEN_7625; // @[rob.scala 411:{25,25}]
  wire  _GEN_7627 = 5'h16 == com_idx ? rob_uop_22_is_sys_pc2epc : _GEN_7626; // @[rob.scala 411:{25,25}]
  wire  _GEN_7628 = 5'h17 == com_idx ? rob_uop_23_is_sys_pc2epc : _GEN_7627; // @[rob.scala 411:{25,25}]
  wire  _GEN_7629 = 5'h18 == com_idx ? rob_uop_24_is_sys_pc2epc : _GEN_7628; // @[rob.scala 411:{25,25}]
  wire  _GEN_7630 = 5'h19 == com_idx ? rob_uop_25_is_sys_pc2epc : _GEN_7629; // @[rob.scala 411:{25,25}]
  wire  _GEN_7631 = 5'h1a == com_idx ? rob_uop_26_is_sys_pc2epc : _GEN_7630; // @[rob.scala 411:{25,25}]
  wire  _GEN_7632 = 5'h1b == com_idx ? rob_uop_27_is_sys_pc2epc : _GEN_7631; // @[rob.scala 411:{25,25}]
  wire  _GEN_7633 = 5'h1c == com_idx ? rob_uop_28_is_sys_pc2epc : _GEN_7632; // @[rob.scala 411:{25,25}]
  wire  _GEN_7634 = 5'h1d == com_idx ? rob_uop_29_is_sys_pc2epc : _GEN_7633; // @[rob.scala 411:{25,25}]
  wire  _GEN_7635 = 5'h1e == com_idx ? rob_uop_30_is_sys_pc2epc : _GEN_7634; // @[rob.scala 411:{25,25}]
  wire  _GEN_7638 = 5'h1 == com_idx ? rob_uop_1_uses_stq : rob_uop_0_uses_stq; // @[rob.scala 411:{25,25}]
  wire  _GEN_7639 = 5'h2 == com_idx ? rob_uop_2_uses_stq : _GEN_7638; // @[rob.scala 411:{25,25}]
  wire  _GEN_7640 = 5'h3 == com_idx ? rob_uop_3_uses_stq : _GEN_7639; // @[rob.scala 411:{25,25}]
  wire  _GEN_7641 = 5'h4 == com_idx ? rob_uop_4_uses_stq : _GEN_7640; // @[rob.scala 411:{25,25}]
  wire  _GEN_7642 = 5'h5 == com_idx ? rob_uop_5_uses_stq : _GEN_7641; // @[rob.scala 411:{25,25}]
  wire  _GEN_7643 = 5'h6 == com_idx ? rob_uop_6_uses_stq : _GEN_7642; // @[rob.scala 411:{25,25}]
  wire  _GEN_7644 = 5'h7 == com_idx ? rob_uop_7_uses_stq : _GEN_7643; // @[rob.scala 411:{25,25}]
  wire  _GEN_7645 = 5'h8 == com_idx ? rob_uop_8_uses_stq : _GEN_7644; // @[rob.scala 411:{25,25}]
  wire  _GEN_7646 = 5'h9 == com_idx ? rob_uop_9_uses_stq : _GEN_7645; // @[rob.scala 411:{25,25}]
  wire  _GEN_7647 = 5'ha == com_idx ? rob_uop_10_uses_stq : _GEN_7646; // @[rob.scala 411:{25,25}]
  wire  _GEN_7648 = 5'hb == com_idx ? rob_uop_11_uses_stq : _GEN_7647; // @[rob.scala 411:{25,25}]
  wire  _GEN_7649 = 5'hc == com_idx ? rob_uop_12_uses_stq : _GEN_7648; // @[rob.scala 411:{25,25}]
  wire  _GEN_7650 = 5'hd == com_idx ? rob_uop_13_uses_stq : _GEN_7649; // @[rob.scala 411:{25,25}]
  wire  _GEN_7651 = 5'he == com_idx ? rob_uop_14_uses_stq : _GEN_7650; // @[rob.scala 411:{25,25}]
  wire  _GEN_7652 = 5'hf == com_idx ? rob_uop_15_uses_stq : _GEN_7651; // @[rob.scala 411:{25,25}]
  wire  _GEN_7653 = 5'h10 == com_idx ? rob_uop_16_uses_stq : _GEN_7652; // @[rob.scala 411:{25,25}]
  wire  _GEN_7654 = 5'h11 == com_idx ? rob_uop_17_uses_stq : _GEN_7653; // @[rob.scala 411:{25,25}]
  wire  _GEN_7655 = 5'h12 == com_idx ? rob_uop_18_uses_stq : _GEN_7654; // @[rob.scala 411:{25,25}]
  wire  _GEN_7656 = 5'h13 == com_idx ? rob_uop_19_uses_stq : _GEN_7655; // @[rob.scala 411:{25,25}]
  wire  _GEN_7657 = 5'h14 == com_idx ? rob_uop_20_uses_stq : _GEN_7656; // @[rob.scala 411:{25,25}]
  wire  _GEN_7658 = 5'h15 == com_idx ? rob_uop_21_uses_stq : _GEN_7657; // @[rob.scala 411:{25,25}]
  wire  _GEN_7659 = 5'h16 == com_idx ? rob_uop_22_uses_stq : _GEN_7658; // @[rob.scala 411:{25,25}]
  wire  _GEN_7660 = 5'h17 == com_idx ? rob_uop_23_uses_stq : _GEN_7659; // @[rob.scala 411:{25,25}]
  wire  _GEN_7661 = 5'h18 == com_idx ? rob_uop_24_uses_stq : _GEN_7660; // @[rob.scala 411:{25,25}]
  wire  _GEN_7662 = 5'h19 == com_idx ? rob_uop_25_uses_stq : _GEN_7661; // @[rob.scala 411:{25,25}]
  wire  _GEN_7663 = 5'h1a == com_idx ? rob_uop_26_uses_stq : _GEN_7662; // @[rob.scala 411:{25,25}]
  wire  _GEN_7664 = 5'h1b == com_idx ? rob_uop_27_uses_stq : _GEN_7663; // @[rob.scala 411:{25,25}]
  wire  _GEN_7665 = 5'h1c == com_idx ? rob_uop_28_uses_stq : _GEN_7664; // @[rob.scala 411:{25,25}]
  wire  _GEN_7666 = 5'h1d == com_idx ? rob_uop_29_uses_stq : _GEN_7665; // @[rob.scala 411:{25,25}]
  wire  _GEN_7667 = 5'h1e == com_idx ? rob_uop_30_uses_stq : _GEN_7666; // @[rob.scala 411:{25,25}]
  wire  _GEN_7670 = 5'h1 == com_idx ? rob_uop_1_uses_ldq : rob_uop_0_uses_ldq; // @[rob.scala 411:{25,25}]
  wire  _GEN_7671 = 5'h2 == com_idx ? rob_uop_2_uses_ldq : _GEN_7670; // @[rob.scala 411:{25,25}]
  wire  _GEN_7672 = 5'h3 == com_idx ? rob_uop_3_uses_ldq : _GEN_7671; // @[rob.scala 411:{25,25}]
  wire  _GEN_7673 = 5'h4 == com_idx ? rob_uop_4_uses_ldq : _GEN_7672; // @[rob.scala 411:{25,25}]
  wire  _GEN_7674 = 5'h5 == com_idx ? rob_uop_5_uses_ldq : _GEN_7673; // @[rob.scala 411:{25,25}]
  wire  _GEN_7675 = 5'h6 == com_idx ? rob_uop_6_uses_ldq : _GEN_7674; // @[rob.scala 411:{25,25}]
  wire  _GEN_7676 = 5'h7 == com_idx ? rob_uop_7_uses_ldq : _GEN_7675; // @[rob.scala 411:{25,25}]
  wire  _GEN_7677 = 5'h8 == com_idx ? rob_uop_8_uses_ldq : _GEN_7676; // @[rob.scala 411:{25,25}]
  wire  _GEN_7678 = 5'h9 == com_idx ? rob_uop_9_uses_ldq : _GEN_7677; // @[rob.scala 411:{25,25}]
  wire  _GEN_7679 = 5'ha == com_idx ? rob_uop_10_uses_ldq : _GEN_7678; // @[rob.scala 411:{25,25}]
  wire  _GEN_7680 = 5'hb == com_idx ? rob_uop_11_uses_ldq : _GEN_7679; // @[rob.scala 411:{25,25}]
  wire  _GEN_7681 = 5'hc == com_idx ? rob_uop_12_uses_ldq : _GEN_7680; // @[rob.scala 411:{25,25}]
  wire  _GEN_7682 = 5'hd == com_idx ? rob_uop_13_uses_ldq : _GEN_7681; // @[rob.scala 411:{25,25}]
  wire  _GEN_7683 = 5'he == com_idx ? rob_uop_14_uses_ldq : _GEN_7682; // @[rob.scala 411:{25,25}]
  wire  _GEN_7684 = 5'hf == com_idx ? rob_uop_15_uses_ldq : _GEN_7683; // @[rob.scala 411:{25,25}]
  wire  _GEN_7685 = 5'h10 == com_idx ? rob_uop_16_uses_ldq : _GEN_7684; // @[rob.scala 411:{25,25}]
  wire  _GEN_7686 = 5'h11 == com_idx ? rob_uop_17_uses_ldq : _GEN_7685; // @[rob.scala 411:{25,25}]
  wire  _GEN_7687 = 5'h12 == com_idx ? rob_uop_18_uses_ldq : _GEN_7686; // @[rob.scala 411:{25,25}]
  wire  _GEN_7688 = 5'h13 == com_idx ? rob_uop_19_uses_ldq : _GEN_7687; // @[rob.scala 411:{25,25}]
  wire  _GEN_7689 = 5'h14 == com_idx ? rob_uop_20_uses_ldq : _GEN_7688; // @[rob.scala 411:{25,25}]
  wire  _GEN_7690 = 5'h15 == com_idx ? rob_uop_21_uses_ldq : _GEN_7689; // @[rob.scala 411:{25,25}]
  wire  _GEN_7691 = 5'h16 == com_idx ? rob_uop_22_uses_ldq : _GEN_7690; // @[rob.scala 411:{25,25}]
  wire  _GEN_7692 = 5'h17 == com_idx ? rob_uop_23_uses_ldq : _GEN_7691; // @[rob.scala 411:{25,25}]
  wire  _GEN_7693 = 5'h18 == com_idx ? rob_uop_24_uses_ldq : _GEN_7692; // @[rob.scala 411:{25,25}]
  wire  _GEN_7694 = 5'h19 == com_idx ? rob_uop_25_uses_ldq : _GEN_7693; // @[rob.scala 411:{25,25}]
  wire  _GEN_7695 = 5'h1a == com_idx ? rob_uop_26_uses_ldq : _GEN_7694; // @[rob.scala 411:{25,25}]
  wire  _GEN_7696 = 5'h1b == com_idx ? rob_uop_27_uses_ldq : _GEN_7695; // @[rob.scala 411:{25,25}]
  wire  _GEN_7697 = 5'h1c == com_idx ? rob_uop_28_uses_ldq : _GEN_7696; // @[rob.scala 411:{25,25}]
  wire  _GEN_7698 = 5'h1d == com_idx ? rob_uop_29_uses_ldq : _GEN_7697; // @[rob.scala 411:{25,25}]
  wire  _GEN_7699 = 5'h1e == com_idx ? rob_uop_30_uses_ldq : _GEN_7698; // @[rob.scala 411:{25,25}]
  wire  _GEN_7702 = 5'h1 == com_idx ? rob_uop_1_is_amo : rob_uop_0_is_amo; // @[rob.scala 411:{25,25}]
  wire  _GEN_7703 = 5'h2 == com_idx ? rob_uop_2_is_amo : _GEN_7702; // @[rob.scala 411:{25,25}]
  wire  _GEN_7704 = 5'h3 == com_idx ? rob_uop_3_is_amo : _GEN_7703; // @[rob.scala 411:{25,25}]
  wire  _GEN_7705 = 5'h4 == com_idx ? rob_uop_4_is_amo : _GEN_7704; // @[rob.scala 411:{25,25}]
  wire  _GEN_7706 = 5'h5 == com_idx ? rob_uop_5_is_amo : _GEN_7705; // @[rob.scala 411:{25,25}]
  wire  _GEN_7707 = 5'h6 == com_idx ? rob_uop_6_is_amo : _GEN_7706; // @[rob.scala 411:{25,25}]
  wire  _GEN_7708 = 5'h7 == com_idx ? rob_uop_7_is_amo : _GEN_7707; // @[rob.scala 411:{25,25}]
  wire  _GEN_7709 = 5'h8 == com_idx ? rob_uop_8_is_amo : _GEN_7708; // @[rob.scala 411:{25,25}]
  wire  _GEN_7710 = 5'h9 == com_idx ? rob_uop_9_is_amo : _GEN_7709; // @[rob.scala 411:{25,25}]
  wire  _GEN_7711 = 5'ha == com_idx ? rob_uop_10_is_amo : _GEN_7710; // @[rob.scala 411:{25,25}]
  wire  _GEN_7712 = 5'hb == com_idx ? rob_uop_11_is_amo : _GEN_7711; // @[rob.scala 411:{25,25}]
  wire  _GEN_7713 = 5'hc == com_idx ? rob_uop_12_is_amo : _GEN_7712; // @[rob.scala 411:{25,25}]
  wire  _GEN_7714 = 5'hd == com_idx ? rob_uop_13_is_amo : _GEN_7713; // @[rob.scala 411:{25,25}]
  wire  _GEN_7715 = 5'he == com_idx ? rob_uop_14_is_amo : _GEN_7714; // @[rob.scala 411:{25,25}]
  wire  _GEN_7716 = 5'hf == com_idx ? rob_uop_15_is_amo : _GEN_7715; // @[rob.scala 411:{25,25}]
  wire  _GEN_7717 = 5'h10 == com_idx ? rob_uop_16_is_amo : _GEN_7716; // @[rob.scala 411:{25,25}]
  wire  _GEN_7718 = 5'h11 == com_idx ? rob_uop_17_is_amo : _GEN_7717; // @[rob.scala 411:{25,25}]
  wire  _GEN_7719 = 5'h12 == com_idx ? rob_uop_18_is_amo : _GEN_7718; // @[rob.scala 411:{25,25}]
  wire  _GEN_7720 = 5'h13 == com_idx ? rob_uop_19_is_amo : _GEN_7719; // @[rob.scala 411:{25,25}]
  wire  _GEN_7721 = 5'h14 == com_idx ? rob_uop_20_is_amo : _GEN_7720; // @[rob.scala 411:{25,25}]
  wire  _GEN_7722 = 5'h15 == com_idx ? rob_uop_21_is_amo : _GEN_7721; // @[rob.scala 411:{25,25}]
  wire  _GEN_7723 = 5'h16 == com_idx ? rob_uop_22_is_amo : _GEN_7722; // @[rob.scala 411:{25,25}]
  wire  _GEN_7724 = 5'h17 == com_idx ? rob_uop_23_is_amo : _GEN_7723; // @[rob.scala 411:{25,25}]
  wire  _GEN_7725 = 5'h18 == com_idx ? rob_uop_24_is_amo : _GEN_7724; // @[rob.scala 411:{25,25}]
  wire  _GEN_7726 = 5'h19 == com_idx ? rob_uop_25_is_amo : _GEN_7725; // @[rob.scala 411:{25,25}]
  wire  _GEN_7727 = 5'h1a == com_idx ? rob_uop_26_is_amo : _GEN_7726; // @[rob.scala 411:{25,25}]
  wire  _GEN_7728 = 5'h1b == com_idx ? rob_uop_27_is_amo : _GEN_7727; // @[rob.scala 411:{25,25}]
  wire  _GEN_7729 = 5'h1c == com_idx ? rob_uop_28_is_amo : _GEN_7728; // @[rob.scala 411:{25,25}]
  wire  _GEN_7730 = 5'h1d == com_idx ? rob_uop_29_is_amo : _GEN_7729; // @[rob.scala 411:{25,25}]
  wire  _GEN_7731 = 5'h1e == com_idx ? rob_uop_30_is_amo : _GEN_7730; // @[rob.scala 411:{25,25}]
  wire  _GEN_7734 = 5'h1 == com_idx ? rob_uop_1_is_fencei : rob_uop_0_is_fencei; // @[rob.scala 411:{25,25}]
  wire  _GEN_7735 = 5'h2 == com_idx ? rob_uop_2_is_fencei : _GEN_7734; // @[rob.scala 411:{25,25}]
  wire  _GEN_7736 = 5'h3 == com_idx ? rob_uop_3_is_fencei : _GEN_7735; // @[rob.scala 411:{25,25}]
  wire  _GEN_7737 = 5'h4 == com_idx ? rob_uop_4_is_fencei : _GEN_7736; // @[rob.scala 411:{25,25}]
  wire  _GEN_7738 = 5'h5 == com_idx ? rob_uop_5_is_fencei : _GEN_7737; // @[rob.scala 411:{25,25}]
  wire  _GEN_7739 = 5'h6 == com_idx ? rob_uop_6_is_fencei : _GEN_7738; // @[rob.scala 411:{25,25}]
  wire  _GEN_7740 = 5'h7 == com_idx ? rob_uop_7_is_fencei : _GEN_7739; // @[rob.scala 411:{25,25}]
  wire  _GEN_7741 = 5'h8 == com_idx ? rob_uop_8_is_fencei : _GEN_7740; // @[rob.scala 411:{25,25}]
  wire  _GEN_7742 = 5'h9 == com_idx ? rob_uop_9_is_fencei : _GEN_7741; // @[rob.scala 411:{25,25}]
  wire  _GEN_7743 = 5'ha == com_idx ? rob_uop_10_is_fencei : _GEN_7742; // @[rob.scala 411:{25,25}]
  wire  _GEN_7744 = 5'hb == com_idx ? rob_uop_11_is_fencei : _GEN_7743; // @[rob.scala 411:{25,25}]
  wire  _GEN_7745 = 5'hc == com_idx ? rob_uop_12_is_fencei : _GEN_7744; // @[rob.scala 411:{25,25}]
  wire  _GEN_7746 = 5'hd == com_idx ? rob_uop_13_is_fencei : _GEN_7745; // @[rob.scala 411:{25,25}]
  wire  _GEN_7747 = 5'he == com_idx ? rob_uop_14_is_fencei : _GEN_7746; // @[rob.scala 411:{25,25}]
  wire  _GEN_7748 = 5'hf == com_idx ? rob_uop_15_is_fencei : _GEN_7747; // @[rob.scala 411:{25,25}]
  wire  _GEN_7749 = 5'h10 == com_idx ? rob_uop_16_is_fencei : _GEN_7748; // @[rob.scala 411:{25,25}]
  wire  _GEN_7750 = 5'h11 == com_idx ? rob_uop_17_is_fencei : _GEN_7749; // @[rob.scala 411:{25,25}]
  wire  _GEN_7751 = 5'h12 == com_idx ? rob_uop_18_is_fencei : _GEN_7750; // @[rob.scala 411:{25,25}]
  wire  _GEN_7752 = 5'h13 == com_idx ? rob_uop_19_is_fencei : _GEN_7751; // @[rob.scala 411:{25,25}]
  wire  _GEN_7753 = 5'h14 == com_idx ? rob_uop_20_is_fencei : _GEN_7752; // @[rob.scala 411:{25,25}]
  wire  _GEN_7754 = 5'h15 == com_idx ? rob_uop_21_is_fencei : _GEN_7753; // @[rob.scala 411:{25,25}]
  wire  _GEN_7755 = 5'h16 == com_idx ? rob_uop_22_is_fencei : _GEN_7754; // @[rob.scala 411:{25,25}]
  wire  _GEN_7756 = 5'h17 == com_idx ? rob_uop_23_is_fencei : _GEN_7755; // @[rob.scala 411:{25,25}]
  wire  _GEN_7757 = 5'h18 == com_idx ? rob_uop_24_is_fencei : _GEN_7756; // @[rob.scala 411:{25,25}]
  wire  _GEN_7758 = 5'h19 == com_idx ? rob_uop_25_is_fencei : _GEN_7757; // @[rob.scala 411:{25,25}]
  wire  _GEN_7759 = 5'h1a == com_idx ? rob_uop_26_is_fencei : _GEN_7758; // @[rob.scala 411:{25,25}]
  wire  _GEN_7760 = 5'h1b == com_idx ? rob_uop_27_is_fencei : _GEN_7759; // @[rob.scala 411:{25,25}]
  wire  _GEN_7761 = 5'h1c == com_idx ? rob_uop_28_is_fencei : _GEN_7760; // @[rob.scala 411:{25,25}]
  wire  _GEN_7762 = 5'h1d == com_idx ? rob_uop_29_is_fencei : _GEN_7761; // @[rob.scala 411:{25,25}]
  wire  _GEN_7763 = 5'h1e == com_idx ? rob_uop_30_is_fencei : _GEN_7762; // @[rob.scala 411:{25,25}]
  wire  _GEN_7766 = 5'h1 == com_idx ? rob_uop_1_is_fence : rob_uop_0_is_fence; // @[rob.scala 411:{25,25}]
  wire  _GEN_7767 = 5'h2 == com_idx ? rob_uop_2_is_fence : _GEN_7766; // @[rob.scala 411:{25,25}]
  wire  _GEN_7768 = 5'h3 == com_idx ? rob_uop_3_is_fence : _GEN_7767; // @[rob.scala 411:{25,25}]
  wire  _GEN_7769 = 5'h4 == com_idx ? rob_uop_4_is_fence : _GEN_7768; // @[rob.scala 411:{25,25}]
  wire  _GEN_7770 = 5'h5 == com_idx ? rob_uop_5_is_fence : _GEN_7769; // @[rob.scala 411:{25,25}]
  wire  _GEN_7771 = 5'h6 == com_idx ? rob_uop_6_is_fence : _GEN_7770; // @[rob.scala 411:{25,25}]
  wire  _GEN_7772 = 5'h7 == com_idx ? rob_uop_7_is_fence : _GEN_7771; // @[rob.scala 411:{25,25}]
  wire  _GEN_7773 = 5'h8 == com_idx ? rob_uop_8_is_fence : _GEN_7772; // @[rob.scala 411:{25,25}]
  wire  _GEN_7774 = 5'h9 == com_idx ? rob_uop_9_is_fence : _GEN_7773; // @[rob.scala 411:{25,25}]
  wire  _GEN_7775 = 5'ha == com_idx ? rob_uop_10_is_fence : _GEN_7774; // @[rob.scala 411:{25,25}]
  wire  _GEN_7776 = 5'hb == com_idx ? rob_uop_11_is_fence : _GEN_7775; // @[rob.scala 411:{25,25}]
  wire  _GEN_7777 = 5'hc == com_idx ? rob_uop_12_is_fence : _GEN_7776; // @[rob.scala 411:{25,25}]
  wire  _GEN_7778 = 5'hd == com_idx ? rob_uop_13_is_fence : _GEN_7777; // @[rob.scala 411:{25,25}]
  wire  _GEN_7779 = 5'he == com_idx ? rob_uop_14_is_fence : _GEN_7778; // @[rob.scala 411:{25,25}]
  wire  _GEN_7780 = 5'hf == com_idx ? rob_uop_15_is_fence : _GEN_7779; // @[rob.scala 411:{25,25}]
  wire  _GEN_7781 = 5'h10 == com_idx ? rob_uop_16_is_fence : _GEN_7780; // @[rob.scala 411:{25,25}]
  wire  _GEN_7782 = 5'h11 == com_idx ? rob_uop_17_is_fence : _GEN_7781; // @[rob.scala 411:{25,25}]
  wire  _GEN_7783 = 5'h12 == com_idx ? rob_uop_18_is_fence : _GEN_7782; // @[rob.scala 411:{25,25}]
  wire  _GEN_7784 = 5'h13 == com_idx ? rob_uop_19_is_fence : _GEN_7783; // @[rob.scala 411:{25,25}]
  wire  _GEN_7785 = 5'h14 == com_idx ? rob_uop_20_is_fence : _GEN_7784; // @[rob.scala 411:{25,25}]
  wire  _GEN_7786 = 5'h15 == com_idx ? rob_uop_21_is_fence : _GEN_7785; // @[rob.scala 411:{25,25}]
  wire  _GEN_7787 = 5'h16 == com_idx ? rob_uop_22_is_fence : _GEN_7786; // @[rob.scala 411:{25,25}]
  wire  _GEN_7788 = 5'h17 == com_idx ? rob_uop_23_is_fence : _GEN_7787; // @[rob.scala 411:{25,25}]
  wire  _GEN_7789 = 5'h18 == com_idx ? rob_uop_24_is_fence : _GEN_7788; // @[rob.scala 411:{25,25}]
  wire  _GEN_7790 = 5'h19 == com_idx ? rob_uop_25_is_fence : _GEN_7789; // @[rob.scala 411:{25,25}]
  wire  _GEN_7791 = 5'h1a == com_idx ? rob_uop_26_is_fence : _GEN_7790; // @[rob.scala 411:{25,25}]
  wire  _GEN_7792 = 5'h1b == com_idx ? rob_uop_27_is_fence : _GEN_7791; // @[rob.scala 411:{25,25}]
  wire  _GEN_7793 = 5'h1c == com_idx ? rob_uop_28_is_fence : _GEN_7792; // @[rob.scala 411:{25,25}]
  wire  _GEN_7794 = 5'h1d == com_idx ? rob_uop_29_is_fence : _GEN_7793; // @[rob.scala 411:{25,25}]
  wire  _GEN_7795 = 5'h1e == com_idx ? rob_uop_30_is_fence : _GEN_7794; // @[rob.scala 411:{25,25}]
  wire  _GEN_7798 = 5'h1 == com_idx ? rob_uop_1_mem_signed : rob_uop_0_mem_signed; // @[rob.scala 411:{25,25}]
  wire  _GEN_7799 = 5'h2 == com_idx ? rob_uop_2_mem_signed : _GEN_7798; // @[rob.scala 411:{25,25}]
  wire  _GEN_7800 = 5'h3 == com_idx ? rob_uop_3_mem_signed : _GEN_7799; // @[rob.scala 411:{25,25}]
  wire  _GEN_7801 = 5'h4 == com_idx ? rob_uop_4_mem_signed : _GEN_7800; // @[rob.scala 411:{25,25}]
  wire  _GEN_7802 = 5'h5 == com_idx ? rob_uop_5_mem_signed : _GEN_7801; // @[rob.scala 411:{25,25}]
  wire  _GEN_7803 = 5'h6 == com_idx ? rob_uop_6_mem_signed : _GEN_7802; // @[rob.scala 411:{25,25}]
  wire  _GEN_7804 = 5'h7 == com_idx ? rob_uop_7_mem_signed : _GEN_7803; // @[rob.scala 411:{25,25}]
  wire  _GEN_7805 = 5'h8 == com_idx ? rob_uop_8_mem_signed : _GEN_7804; // @[rob.scala 411:{25,25}]
  wire  _GEN_7806 = 5'h9 == com_idx ? rob_uop_9_mem_signed : _GEN_7805; // @[rob.scala 411:{25,25}]
  wire  _GEN_7807 = 5'ha == com_idx ? rob_uop_10_mem_signed : _GEN_7806; // @[rob.scala 411:{25,25}]
  wire  _GEN_7808 = 5'hb == com_idx ? rob_uop_11_mem_signed : _GEN_7807; // @[rob.scala 411:{25,25}]
  wire  _GEN_7809 = 5'hc == com_idx ? rob_uop_12_mem_signed : _GEN_7808; // @[rob.scala 411:{25,25}]
  wire  _GEN_7810 = 5'hd == com_idx ? rob_uop_13_mem_signed : _GEN_7809; // @[rob.scala 411:{25,25}]
  wire  _GEN_7811 = 5'he == com_idx ? rob_uop_14_mem_signed : _GEN_7810; // @[rob.scala 411:{25,25}]
  wire  _GEN_7812 = 5'hf == com_idx ? rob_uop_15_mem_signed : _GEN_7811; // @[rob.scala 411:{25,25}]
  wire  _GEN_7813 = 5'h10 == com_idx ? rob_uop_16_mem_signed : _GEN_7812; // @[rob.scala 411:{25,25}]
  wire  _GEN_7814 = 5'h11 == com_idx ? rob_uop_17_mem_signed : _GEN_7813; // @[rob.scala 411:{25,25}]
  wire  _GEN_7815 = 5'h12 == com_idx ? rob_uop_18_mem_signed : _GEN_7814; // @[rob.scala 411:{25,25}]
  wire  _GEN_7816 = 5'h13 == com_idx ? rob_uop_19_mem_signed : _GEN_7815; // @[rob.scala 411:{25,25}]
  wire  _GEN_7817 = 5'h14 == com_idx ? rob_uop_20_mem_signed : _GEN_7816; // @[rob.scala 411:{25,25}]
  wire  _GEN_7818 = 5'h15 == com_idx ? rob_uop_21_mem_signed : _GEN_7817; // @[rob.scala 411:{25,25}]
  wire  _GEN_7819 = 5'h16 == com_idx ? rob_uop_22_mem_signed : _GEN_7818; // @[rob.scala 411:{25,25}]
  wire  _GEN_7820 = 5'h17 == com_idx ? rob_uop_23_mem_signed : _GEN_7819; // @[rob.scala 411:{25,25}]
  wire  _GEN_7821 = 5'h18 == com_idx ? rob_uop_24_mem_signed : _GEN_7820; // @[rob.scala 411:{25,25}]
  wire  _GEN_7822 = 5'h19 == com_idx ? rob_uop_25_mem_signed : _GEN_7821; // @[rob.scala 411:{25,25}]
  wire  _GEN_7823 = 5'h1a == com_idx ? rob_uop_26_mem_signed : _GEN_7822; // @[rob.scala 411:{25,25}]
  wire  _GEN_7824 = 5'h1b == com_idx ? rob_uop_27_mem_signed : _GEN_7823; // @[rob.scala 411:{25,25}]
  wire  _GEN_7825 = 5'h1c == com_idx ? rob_uop_28_mem_signed : _GEN_7824; // @[rob.scala 411:{25,25}]
  wire  _GEN_7826 = 5'h1d == com_idx ? rob_uop_29_mem_signed : _GEN_7825; // @[rob.scala 411:{25,25}]
  wire  _GEN_7827 = 5'h1e == com_idx ? rob_uop_30_mem_signed : _GEN_7826; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7830 = 5'h1 == com_idx ? rob_uop_1_mem_size : rob_uop_0_mem_size; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7831 = 5'h2 == com_idx ? rob_uop_2_mem_size : _GEN_7830; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7832 = 5'h3 == com_idx ? rob_uop_3_mem_size : _GEN_7831; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7833 = 5'h4 == com_idx ? rob_uop_4_mem_size : _GEN_7832; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7834 = 5'h5 == com_idx ? rob_uop_5_mem_size : _GEN_7833; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7835 = 5'h6 == com_idx ? rob_uop_6_mem_size : _GEN_7834; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7836 = 5'h7 == com_idx ? rob_uop_7_mem_size : _GEN_7835; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7837 = 5'h8 == com_idx ? rob_uop_8_mem_size : _GEN_7836; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7838 = 5'h9 == com_idx ? rob_uop_9_mem_size : _GEN_7837; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7839 = 5'ha == com_idx ? rob_uop_10_mem_size : _GEN_7838; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7840 = 5'hb == com_idx ? rob_uop_11_mem_size : _GEN_7839; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7841 = 5'hc == com_idx ? rob_uop_12_mem_size : _GEN_7840; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7842 = 5'hd == com_idx ? rob_uop_13_mem_size : _GEN_7841; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7843 = 5'he == com_idx ? rob_uop_14_mem_size : _GEN_7842; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7844 = 5'hf == com_idx ? rob_uop_15_mem_size : _GEN_7843; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7845 = 5'h10 == com_idx ? rob_uop_16_mem_size : _GEN_7844; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7846 = 5'h11 == com_idx ? rob_uop_17_mem_size : _GEN_7845; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7847 = 5'h12 == com_idx ? rob_uop_18_mem_size : _GEN_7846; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7848 = 5'h13 == com_idx ? rob_uop_19_mem_size : _GEN_7847; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7849 = 5'h14 == com_idx ? rob_uop_20_mem_size : _GEN_7848; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7850 = 5'h15 == com_idx ? rob_uop_21_mem_size : _GEN_7849; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7851 = 5'h16 == com_idx ? rob_uop_22_mem_size : _GEN_7850; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7852 = 5'h17 == com_idx ? rob_uop_23_mem_size : _GEN_7851; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7853 = 5'h18 == com_idx ? rob_uop_24_mem_size : _GEN_7852; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7854 = 5'h19 == com_idx ? rob_uop_25_mem_size : _GEN_7853; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7855 = 5'h1a == com_idx ? rob_uop_26_mem_size : _GEN_7854; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7856 = 5'h1b == com_idx ? rob_uop_27_mem_size : _GEN_7855; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7857 = 5'h1c == com_idx ? rob_uop_28_mem_size : _GEN_7856; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7858 = 5'h1d == com_idx ? rob_uop_29_mem_size : _GEN_7857; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_7859 = 5'h1e == com_idx ? rob_uop_30_mem_size : _GEN_7858; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7862 = 5'h1 == com_idx ? rob_uop_1_mem_cmd : rob_uop_0_mem_cmd; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7863 = 5'h2 == com_idx ? rob_uop_2_mem_cmd : _GEN_7862; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7864 = 5'h3 == com_idx ? rob_uop_3_mem_cmd : _GEN_7863; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7865 = 5'h4 == com_idx ? rob_uop_4_mem_cmd : _GEN_7864; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7866 = 5'h5 == com_idx ? rob_uop_5_mem_cmd : _GEN_7865; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7867 = 5'h6 == com_idx ? rob_uop_6_mem_cmd : _GEN_7866; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7868 = 5'h7 == com_idx ? rob_uop_7_mem_cmd : _GEN_7867; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7869 = 5'h8 == com_idx ? rob_uop_8_mem_cmd : _GEN_7868; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7870 = 5'h9 == com_idx ? rob_uop_9_mem_cmd : _GEN_7869; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7871 = 5'ha == com_idx ? rob_uop_10_mem_cmd : _GEN_7870; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7872 = 5'hb == com_idx ? rob_uop_11_mem_cmd : _GEN_7871; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7873 = 5'hc == com_idx ? rob_uop_12_mem_cmd : _GEN_7872; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7874 = 5'hd == com_idx ? rob_uop_13_mem_cmd : _GEN_7873; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7875 = 5'he == com_idx ? rob_uop_14_mem_cmd : _GEN_7874; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7876 = 5'hf == com_idx ? rob_uop_15_mem_cmd : _GEN_7875; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7877 = 5'h10 == com_idx ? rob_uop_16_mem_cmd : _GEN_7876; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7878 = 5'h11 == com_idx ? rob_uop_17_mem_cmd : _GEN_7877; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7879 = 5'h12 == com_idx ? rob_uop_18_mem_cmd : _GEN_7878; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7880 = 5'h13 == com_idx ? rob_uop_19_mem_cmd : _GEN_7879; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7881 = 5'h14 == com_idx ? rob_uop_20_mem_cmd : _GEN_7880; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7882 = 5'h15 == com_idx ? rob_uop_21_mem_cmd : _GEN_7881; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7883 = 5'h16 == com_idx ? rob_uop_22_mem_cmd : _GEN_7882; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7884 = 5'h17 == com_idx ? rob_uop_23_mem_cmd : _GEN_7883; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7885 = 5'h18 == com_idx ? rob_uop_24_mem_cmd : _GEN_7884; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7886 = 5'h19 == com_idx ? rob_uop_25_mem_cmd : _GEN_7885; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7887 = 5'h1a == com_idx ? rob_uop_26_mem_cmd : _GEN_7886; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7888 = 5'h1b == com_idx ? rob_uop_27_mem_cmd : _GEN_7887; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7889 = 5'h1c == com_idx ? rob_uop_28_mem_cmd : _GEN_7888; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7890 = 5'h1d == com_idx ? rob_uop_29_mem_cmd : _GEN_7889; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_7891 = 5'h1e == com_idx ? rob_uop_30_mem_cmd : _GEN_7890; // @[rob.scala 411:{25,25}]
  wire  _GEN_7894 = 5'h1 == com_idx ? rob_uop_1_bypassable : rob_uop_0_bypassable; // @[rob.scala 411:{25,25}]
  wire  _GEN_7895 = 5'h2 == com_idx ? rob_uop_2_bypassable : _GEN_7894; // @[rob.scala 411:{25,25}]
  wire  _GEN_7896 = 5'h3 == com_idx ? rob_uop_3_bypassable : _GEN_7895; // @[rob.scala 411:{25,25}]
  wire  _GEN_7897 = 5'h4 == com_idx ? rob_uop_4_bypassable : _GEN_7896; // @[rob.scala 411:{25,25}]
  wire  _GEN_7898 = 5'h5 == com_idx ? rob_uop_5_bypassable : _GEN_7897; // @[rob.scala 411:{25,25}]
  wire  _GEN_7899 = 5'h6 == com_idx ? rob_uop_6_bypassable : _GEN_7898; // @[rob.scala 411:{25,25}]
  wire  _GEN_7900 = 5'h7 == com_idx ? rob_uop_7_bypassable : _GEN_7899; // @[rob.scala 411:{25,25}]
  wire  _GEN_7901 = 5'h8 == com_idx ? rob_uop_8_bypassable : _GEN_7900; // @[rob.scala 411:{25,25}]
  wire  _GEN_7902 = 5'h9 == com_idx ? rob_uop_9_bypassable : _GEN_7901; // @[rob.scala 411:{25,25}]
  wire  _GEN_7903 = 5'ha == com_idx ? rob_uop_10_bypassable : _GEN_7902; // @[rob.scala 411:{25,25}]
  wire  _GEN_7904 = 5'hb == com_idx ? rob_uop_11_bypassable : _GEN_7903; // @[rob.scala 411:{25,25}]
  wire  _GEN_7905 = 5'hc == com_idx ? rob_uop_12_bypassable : _GEN_7904; // @[rob.scala 411:{25,25}]
  wire  _GEN_7906 = 5'hd == com_idx ? rob_uop_13_bypassable : _GEN_7905; // @[rob.scala 411:{25,25}]
  wire  _GEN_7907 = 5'he == com_idx ? rob_uop_14_bypassable : _GEN_7906; // @[rob.scala 411:{25,25}]
  wire  _GEN_7908 = 5'hf == com_idx ? rob_uop_15_bypassable : _GEN_7907; // @[rob.scala 411:{25,25}]
  wire  _GEN_7909 = 5'h10 == com_idx ? rob_uop_16_bypassable : _GEN_7908; // @[rob.scala 411:{25,25}]
  wire  _GEN_7910 = 5'h11 == com_idx ? rob_uop_17_bypassable : _GEN_7909; // @[rob.scala 411:{25,25}]
  wire  _GEN_7911 = 5'h12 == com_idx ? rob_uop_18_bypassable : _GEN_7910; // @[rob.scala 411:{25,25}]
  wire  _GEN_7912 = 5'h13 == com_idx ? rob_uop_19_bypassable : _GEN_7911; // @[rob.scala 411:{25,25}]
  wire  _GEN_7913 = 5'h14 == com_idx ? rob_uop_20_bypassable : _GEN_7912; // @[rob.scala 411:{25,25}]
  wire  _GEN_7914 = 5'h15 == com_idx ? rob_uop_21_bypassable : _GEN_7913; // @[rob.scala 411:{25,25}]
  wire  _GEN_7915 = 5'h16 == com_idx ? rob_uop_22_bypassable : _GEN_7914; // @[rob.scala 411:{25,25}]
  wire  _GEN_7916 = 5'h17 == com_idx ? rob_uop_23_bypassable : _GEN_7915; // @[rob.scala 411:{25,25}]
  wire  _GEN_7917 = 5'h18 == com_idx ? rob_uop_24_bypassable : _GEN_7916; // @[rob.scala 411:{25,25}]
  wire  _GEN_7918 = 5'h19 == com_idx ? rob_uop_25_bypassable : _GEN_7917; // @[rob.scala 411:{25,25}]
  wire  _GEN_7919 = 5'h1a == com_idx ? rob_uop_26_bypassable : _GEN_7918; // @[rob.scala 411:{25,25}]
  wire  _GEN_7920 = 5'h1b == com_idx ? rob_uop_27_bypassable : _GEN_7919; // @[rob.scala 411:{25,25}]
  wire  _GEN_7921 = 5'h1c == com_idx ? rob_uop_28_bypassable : _GEN_7920; // @[rob.scala 411:{25,25}]
  wire  _GEN_7922 = 5'h1d == com_idx ? rob_uop_29_bypassable : _GEN_7921; // @[rob.scala 411:{25,25}]
  wire  _GEN_7923 = 5'h1e == com_idx ? rob_uop_30_bypassable : _GEN_7922; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7926 = 5'h1 == com_idx ? rob_uop_1_exc_cause : rob_uop_0_exc_cause; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7927 = 5'h2 == com_idx ? rob_uop_2_exc_cause : _GEN_7926; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7928 = 5'h3 == com_idx ? rob_uop_3_exc_cause : _GEN_7927; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7929 = 5'h4 == com_idx ? rob_uop_4_exc_cause : _GEN_7928; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7930 = 5'h5 == com_idx ? rob_uop_5_exc_cause : _GEN_7929; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7931 = 5'h6 == com_idx ? rob_uop_6_exc_cause : _GEN_7930; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7932 = 5'h7 == com_idx ? rob_uop_7_exc_cause : _GEN_7931; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7933 = 5'h8 == com_idx ? rob_uop_8_exc_cause : _GEN_7932; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7934 = 5'h9 == com_idx ? rob_uop_9_exc_cause : _GEN_7933; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7935 = 5'ha == com_idx ? rob_uop_10_exc_cause : _GEN_7934; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7936 = 5'hb == com_idx ? rob_uop_11_exc_cause : _GEN_7935; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7937 = 5'hc == com_idx ? rob_uop_12_exc_cause : _GEN_7936; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7938 = 5'hd == com_idx ? rob_uop_13_exc_cause : _GEN_7937; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7939 = 5'he == com_idx ? rob_uop_14_exc_cause : _GEN_7938; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7940 = 5'hf == com_idx ? rob_uop_15_exc_cause : _GEN_7939; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7941 = 5'h10 == com_idx ? rob_uop_16_exc_cause : _GEN_7940; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7942 = 5'h11 == com_idx ? rob_uop_17_exc_cause : _GEN_7941; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7943 = 5'h12 == com_idx ? rob_uop_18_exc_cause : _GEN_7942; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7944 = 5'h13 == com_idx ? rob_uop_19_exc_cause : _GEN_7943; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7945 = 5'h14 == com_idx ? rob_uop_20_exc_cause : _GEN_7944; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7946 = 5'h15 == com_idx ? rob_uop_21_exc_cause : _GEN_7945; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7947 = 5'h16 == com_idx ? rob_uop_22_exc_cause : _GEN_7946; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7948 = 5'h17 == com_idx ? rob_uop_23_exc_cause : _GEN_7947; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7949 = 5'h18 == com_idx ? rob_uop_24_exc_cause : _GEN_7948; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7950 = 5'h19 == com_idx ? rob_uop_25_exc_cause : _GEN_7949; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7951 = 5'h1a == com_idx ? rob_uop_26_exc_cause : _GEN_7950; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7952 = 5'h1b == com_idx ? rob_uop_27_exc_cause : _GEN_7951; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7953 = 5'h1c == com_idx ? rob_uop_28_exc_cause : _GEN_7952; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7954 = 5'h1d == com_idx ? rob_uop_29_exc_cause : _GEN_7953; // @[rob.scala 411:{25,25}]
  wire [63:0] _GEN_7955 = 5'h1e == com_idx ? rob_uop_30_exc_cause : _GEN_7954; // @[rob.scala 411:{25,25}]
  wire  _GEN_7958 = 5'h1 == com_idx ? rob_uop_1_exception : rob_uop_0_exception; // @[rob.scala 411:{25,25}]
  wire  _GEN_7959 = 5'h2 == com_idx ? rob_uop_2_exception : _GEN_7958; // @[rob.scala 411:{25,25}]
  wire  _GEN_7960 = 5'h3 == com_idx ? rob_uop_3_exception : _GEN_7959; // @[rob.scala 411:{25,25}]
  wire  _GEN_7961 = 5'h4 == com_idx ? rob_uop_4_exception : _GEN_7960; // @[rob.scala 411:{25,25}]
  wire  _GEN_7962 = 5'h5 == com_idx ? rob_uop_5_exception : _GEN_7961; // @[rob.scala 411:{25,25}]
  wire  _GEN_7963 = 5'h6 == com_idx ? rob_uop_6_exception : _GEN_7962; // @[rob.scala 411:{25,25}]
  wire  _GEN_7964 = 5'h7 == com_idx ? rob_uop_7_exception : _GEN_7963; // @[rob.scala 411:{25,25}]
  wire  _GEN_7965 = 5'h8 == com_idx ? rob_uop_8_exception : _GEN_7964; // @[rob.scala 411:{25,25}]
  wire  _GEN_7966 = 5'h9 == com_idx ? rob_uop_9_exception : _GEN_7965; // @[rob.scala 411:{25,25}]
  wire  _GEN_7967 = 5'ha == com_idx ? rob_uop_10_exception : _GEN_7966; // @[rob.scala 411:{25,25}]
  wire  _GEN_7968 = 5'hb == com_idx ? rob_uop_11_exception : _GEN_7967; // @[rob.scala 411:{25,25}]
  wire  _GEN_7969 = 5'hc == com_idx ? rob_uop_12_exception : _GEN_7968; // @[rob.scala 411:{25,25}]
  wire  _GEN_7970 = 5'hd == com_idx ? rob_uop_13_exception : _GEN_7969; // @[rob.scala 411:{25,25}]
  wire  _GEN_7971 = 5'he == com_idx ? rob_uop_14_exception : _GEN_7970; // @[rob.scala 411:{25,25}]
  wire  _GEN_7972 = 5'hf == com_idx ? rob_uop_15_exception : _GEN_7971; // @[rob.scala 411:{25,25}]
  wire  _GEN_7973 = 5'h10 == com_idx ? rob_uop_16_exception : _GEN_7972; // @[rob.scala 411:{25,25}]
  wire  _GEN_7974 = 5'h11 == com_idx ? rob_uop_17_exception : _GEN_7973; // @[rob.scala 411:{25,25}]
  wire  _GEN_7975 = 5'h12 == com_idx ? rob_uop_18_exception : _GEN_7974; // @[rob.scala 411:{25,25}]
  wire  _GEN_7976 = 5'h13 == com_idx ? rob_uop_19_exception : _GEN_7975; // @[rob.scala 411:{25,25}]
  wire  _GEN_7977 = 5'h14 == com_idx ? rob_uop_20_exception : _GEN_7976; // @[rob.scala 411:{25,25}]
  wire  _GEN_7978 = 5'h15 == com_idx ? rob_uop_21_exception : _GEN_7977; // @[rob.scala 411:{25,25}]
  wire  _GEN_7979 = 5'h16 == com_idx ? rob_uop_22_exception : _GEN_7978; // @[rob.scala 411:{25,25}]
  wire  _GEN_7980 = 5'h17 == com_idx ? rob_uop_23_exception : _GEN_7979; // @[rob.scala 411:{25,25}]
  wire  _GEN_7981 = 5'h18 == com_idx ? rob_uop_24_exception : _GEN_7980; // @[rob.scala 411:{25,25}]
  wire  _GEN_7982 = 5'h19 == com_idx ? rob_uop_25_exception : _GEN_7981; // @[rob.scala 411:{25,25}]
  wire  _GEN_7983 = 5'h1a == com_idx ? rob_uop_26_exception : _GEN_7982; // @[rob.scala 411:{25,25}]
  wire  _GEN_7984 = 5'h1b == com_idx ? rob_uop_27_exception : _GEN_7983; // @[rob.scala 411:{25,25}]
  wire  _GEN_7985 = 5'h1c == com_idx ? rob_uop_28_exception : _GEN_7984; // @[rob.scala 411:{25,25}]
  wire  _GEN_7986 = 5'h1d == com_idx ? rob_uop_29_exception : _GEN_7985; // @[rob.scala 411:{25,25}]
  wire  _GEN_7987 = 5'h1e == com_idx ? rob_uop_30_exception : _GEN_7986; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7990 = 5'h1 == com_idx ? rob_uop_1_stale_pdst : rob_uop_0_stale_pdst; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7991 = 5'h2 == com_idx ? rob_uop_2_stale_pdst : _GEN_7990; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7992 = 5'h3 == com_idx ? rob_uop_3_stale_pdst : _GEN_7991; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7993 = 5'h4 == com_idx ? rob_uop_4_stale_pdst : _GEN_7992; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7994 = 5'h5 == com_idx ? rob_uop_5_stale_pdst : _GEN_7993; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7995 = 5'h6 == com_idx ? rob_uop_6_stale_pdst : _GEN_7994; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7996 = 5'h7 == com_idx ? rob_uop_7_stale_pdst : _GEN_7995; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7997 = 5'h8 == com_idx ? rob_uop_8_stale_pdst : _GEN_7996; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7998 = 5'h9 == com_idx ? rob_uop_9_stale_pdst : _GEN_7997; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_7999 = 5'ha == com_idx ? rob_uop_10_stale_pdst : _GEN_7998; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8000 = 5'hb == com_idx ? rob_uop_11_stale_pdst : _GEN_7999; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8001 = 5'hc == com_idx ? rob_uop_12_stale_pdst : _GEN_8000; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8002 = 5'hd == com_idx ? rob_uop_13_stale_pdst : _GEN_8001; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8003 = 5'he == com_idx ? rob_uop_14_stale_pdst : _GEN_8002; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8004 = 5'hf == com_idx ? rob_uop_15_stale_pdst : _GEN_8003; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8005 = 5'h10 == com_idx ? rob_uop_16_stale_pdst : _GEN_8004; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8006 = 5'h11 == com_idx ? rob_uop_17_stale_pdst : _GEN_8005; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8007 = 5'h12 == com_idx ? rob_uop_18_stale_pdst : _GEN_8006; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8008 = 5'h13 == com_idx ? rob_uop_19_stale_pdst : _GEN_8007; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8009 = 5'h14 == com_idx ? rob_uop_20_stale_pdst : _GEN_8008; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8010 = 5'h15 == com_idx ? rob_uop_21_stale_pdst : _GEN_8009; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8011 = 5'h16 == com_idx ? rob_uop_22_stale_pdst : _GEN_8010; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8012 = 5'h17 == com_idx ? rob_uop_23_stale_pdst : _GEN_8011; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8013 = 5'h18 == com_idx ? rob_uop_24_stale_pdst : _GEN_8012; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8014 = 5'h19 == com_idx ? rob_uop_25_stale_pdst : _GEN_8013; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8015 = 5'h1a == com_idx ? rob_uop_26_stale_pdst : _GEN_8014; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8016 = 5'h1b == com_idx ? rob_uop_27_stale_pdst : _GEN_8015; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8017 = 5'h1c == com_idx ? rob_uop_28_stale_pdst : _GEN_8016; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8018 = 5'h1d == com_idx ? rob_uop_29_stale_pdst : _GEN_8017; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8019 = 5'h1e == com_idx ? rob_uop_30_stale_pdst : _GEN_8018; // @[rob.scala 411:{25,25}]
  wire  _GEN_8022 = 5'h1 == com_idx ? rob_uop_1_ppred_busy : rob_uop_0_ppred_busy; // @[rob.scala 411:{25,25}]
  wire  _GEN_8023 = 5'h2 == com_idx ? rob_uop_2_ppred_busy : _GEN_8022; // @[rob.scala 411:{25,25}]
  wire  _GEN_8024 = 5'h3 == com_idx ? rob_uop_3_ppred_busy : _GEN_8023; // @[rob.scala 411:{25,25}]
  wire  _GEN_8025 = 5'h4 == com_idx ? rob_uop_4_ppred_busy : _GEN_8024; // @[rob.scala 411:{25,25}]
  wire  _GEN_8026 = 5'h5 == com_idx ? rob_uop_5_ppred_busy : _GEN_8025; // @[rob.scala 411:{25,25}]
  wire  _GEN_8027 = 5'h6 == com_idx ? rob_uop_6_ppred_busy : _GEN_8026; // @[rob.scala 411:{25,25}]
  wire  _GEN_8028 = 5'h7 == com_idx ? rob_uop_7_ppred_busy : _GEN_8027; // @[rob.scala 411:{25,25}]
  wire  _GEN_8029 = 5'h8 == com_idx ? rob_uop_8_ppred_busy : _GEN_8028; // @[rob.scala 411:{25,25}]
  wire  _GEN_8030 = 5'h9 == com_idx ? rob_uop_9_ppred_busy : _GEN_8029; // @[rob.scala 411:{25,25}]
  wire  _GEN_8031 = 5'ha == com_idx ? rob_uop_10_ppred_busy : _GEN_8030; // @[rob.scala 411:{25,25}]
  wire  _GEN_8032 = 5'hb == com_idx ? rob_uop_11_ppred_busy : _GEN_8031; // @[rob.scala 411:{25,25}]
  wire  _GEN_8033 = 5'hc == com_idx ? rob_uop_12_ppred_busy : _GEN_8032; // @[rob.scala 411:{25,25}]
  wire  _GEN_8034 = 5'hd == com_idx ? rob_uop_13_ppred_busy : _GEN_8033; // @[rob.scala 411:{25,25}]
  wire  _GEN_8035 = 5'he == com_idx ? rob_uop_14_ppred_busy : _GEN_8034; // @[rob.scala 411:{25,25}]
  wire  _GEN_8036 = 5'hf == com_idx ? rob_uop_15_ppred_busy : _GEN_8035; // @[rob.scala 411:{25,25}]
  wire  _GEN_8037 = 5'h10 == com_idx ? rob_uop_16_ppred_busy : _GEN_8036; // @[rob.scala 411:{25,25}]
  wire  _GEN_8038 = 5'h11 == com_idx ? rob_uop_17_ppred_busy : _GEN_8037; // @[rob.scala 411:{25,25}]
  wire  _GEN_8039 = 5'h12 == com_idx ? rob_uop_18_ppred_busy : _GEN_8038; // @[rob.scala 411:{25,25}]
  wire  _GEN_8040 = 5'h13 == com_idx ? rob_uop_19_ppred_busy : _GEN_8039; // @[rob.scala 411:{25,25}]
  wire  _GEN_8041 = 5'h14 == com_idx ? rob_uop_20_ppred_busy : _GEN_8040; // @[rob.scala 411:{25,25}]
  wire  _GEN_8042 = 5'h15 == com_idx ? rob_uop_21_ppred_busy : _GEN_8041; // @[rob.scala 411:{25,25}]
  wire  _GEN_8043 = 5'h16 == com_idx ? rob_uop_22_ppred_busy : _GEN_8042; // @[rob.scala 411:{25,25}]
  wire  _GEN_8044 = 5'h17 == com_idx ? rob_uop_23_ppred_busy : _GEN_8043; // @[rob.scala 411:{25,25}]
  wire  _GEN_8045 = 5'h18 == com_idx ? rob_uop_24_ppred_busy : _GEN_8044; // @[rob.scala 411:{25,25}]
  wire  _GEN_8046 = 5'h19 == com_idx ? rob_uop_25_ppred_busy : _GEN_8045; // @[rob.scala 411:{25,25}]
  wire  _GEN_8047 = 5'h1a == com_idx ? rob_uop_26_ppred_busy : _GEN_8046; // @[rob.scala 411:{25,25}]
  wire  _GEN_8048 = 5'h1b == com_idx ? rob_uop_27_ppred_busy : _GEN_8047; // @[rob.scala 411:{25,25}]
  wire  _GEN_8049 = 5'h1c == com_idx ? rob_uop_28_ppred_busy : _GEN_8048; // @[rob.scala 411:{25,25}]
  wire  _GEN_8050 = 5'h1d == com_idx ? rob_uop_29_ppred_busy : _GEN_8049; // @[rob.scala 411:{25,25}]
  wire  _GEN_8051 = 5'h1e == com_idx ? rob_uop_30_ppred_busy : _GEN_8050; // @[rob.scala 411:{25,25}]
  wire  _GEN_8054 = 5'h1 == com_idx ? rob_uop_1_prs3_busy : rob_uop_0_prs3_busy; // @[rob.scala 411:{25,25}]
  wire  _GEN_8055 = 5'h2 == com_idx ? rob_uop_2_prs3_busy : _GEN_8054; // @[rob.scala 411:{25,25}]
  wire  _GEN_8056 = 5'h3 == com_idx ? rob_uop_3_prs3_busy : _GEN_8055; // @[rob.scala 411:{25,25}]
  wire  _GEN_8057 = 5'h4 == com_idx ? rob_uop_4_prs3_busy : _GEN_8056; // @[rob.scala 411:{25,25}]
  wire  _GEN_8058 = 5'h5 == com_idx ? rob_uop_5_prs3_busy : _GEN_8057; // @[rob.scala 411:{25,25}]
  wire  _GEN_8059 = 5'h6 == com_idx ? rob_uop_6_prs3_busy : _GEN_8058; // @[rob.scala 411:{25,25}]
  wire  _GEN_8060 = 5'h7 == com_idx ? rob_uop_7_prs3_busy : _GEN_8059; // @[rob.scala 411:{25,25}]
  wire  _GEN_8061 = 5'h8 == com_idx ? rob_uop_8_prs3_busy : _GEN_8060; // @[rob.scala 411:{25,25}]
  wire  _GEN_8062 = 5'h9 == com_idx ? rob_uop_9_prs3_busy : _GEN_8061; // @[rob.scala 411:{25,25}]
  wire  _GEN_8063 = 5'ha == com_idx ? rob_uop_10_prs3_busy : _GEN_8062; // @[rob.scala 411:{25,25}]
  wire  _GEN_8064 = 5'hb == com_idx ? rob_uop_11_prs3_busy : _GEN_8063; // @[rob.scala 411:{25,25}]
  wire  _GEN_8065 = 5'hc == com_idx ? rob_uop_12_prs3_busy : _GEN_8064; // @[rob.scala 411:{25,25}]
  wire  _GEN_8066 = 5'hd == com_idx ? rob_uop_13_prs3_busy : _GEN_8065; // @[rob.scala 411:{25,25}]
  wire  _GEN_8067 = 5'he == com_idx ? rob_uop_14_prs3_busy : _GEN_8066; // @[rob.scala 411:{25,25}]
  wire  _GEN_8068 = 5'hf == com_idx ? rob_uop_15_prs3_busy : _GEN_8067; // @[rob.scala 411:{25,25}]
  wire  _GEN_8069 = 5'h10 == com_idx ? rob_uop_16_prs3_busy : _GEN_8068; // @[rob.scala 411:{25,25}]
  wire  _GEN_8070 = 5'h11 == com_idx ? rob_uop_17_prs3_busy : _GEN_8069; // @[rob.scala 411:{25,25}]
  wire  _GEN_8071 = 5'h12 == com_idx ? rob_uop_18_prs3_busy : _GEN_8070; // @[rob.scala 411:{25,25}]
  wire  _GEN_8072 = 5'h13 == com_idx ? rob_uop_19_prs3_busy : _GEN_8071; // @[rob.scala 411:{25,25}]
  wire  _GEN_8073 = 5'h14 == com_idx ? rob_uop_20_prs3_busy : _GEN_8072; // @[rob.scala 411:{25,25}]
  wire  _GEN_8074 = 5'h15 == com_idx ? rob_uop_21_prs3_busy : _GEN_8073; // @[rob.scala 411:{25,25}]
  wire  _GEN_8075 = 5'h16 == com_idx ? rob_uop_22_prs3_busy : _GEN_8074; // @[rob.scala 411:{25,25}]
  wire  _GEN_8076 = 5'h17 == com_idx ? rob_uop_23_prs3_busy : _GEN_8075; // @[rob.scala 411:{25,25}]
  wire  _GEN_8077 = 5'h18 == com_idx ? rob_uop_24_prs3_busy : _GEN_8076; // @[rob.scala 411:{25,25}]
  wire  _GEN_8078 = 5'h19 == com_idx ? rob_uop_25_prs3_busy : _GEN_8077; // @[rob.scala 411:{25,25}]
  wire  _GEN_8079 = 5'h1a == com_idx ? rob_uop_26_prs3_busy : _GEN_8078; // @[rob.scala 411:{25,25}]
  wire  _GEN_8080 = 5'h1b == com_idx ? rob_uop_27_prs3_busy : _GEN_8079; // @[rob.scala 411:{25,25}]
  wire  _GEN_8081 = 5'h1c == com_idx ? rob_uop_28_prs3_busy : _GEN_8080; // @[rob.scala 411:{25,25}]
  wire  _GEN_8082 = 5'h1d == com_idx ? rob_uop_29_prs3_busy : _GEN_8081; // @[rob.scala 411:{25,25}]
  wire  _GEN_8083 = 5'h1e == com_idx ? rob_uop_30_prs3_busy : _GEN_8082; // @[rob.scala 411:{25,25}]
  wire  _GEN_8086 = 5'h1 == com_idx ? rob_uop_1_prs2_busy : rob_uop_0_prs2_busy; // @[rob.scala 411:{25,25}]
  wire  _GEN_8087 = 5'h2 == com_idx ? rob_uop_2_prs2_busy : _GEN_8086; // @[rob.scala 411:{25,25}]
  wire  _GEN_8088 = 5'h3 == com_idx ? rob_uop_3_prs2_busy : _GEN_8087; // @[rob.scala 411:{25,25}]
  wire  _GEN_8089 = 5'h4 == com_idx ? rob_uop_4_prs2_busy : _GEN_8088; // @[rob.scala 411:{25,25}]
  wire  _GEN_8090 = 5'h5 == com_idx ? rob_uop_5_prs2_busy : _GEN_8089; // @[rob.scala 411:{25,25}]
  wire  _GEN_8091 = 5'h6 == com_idx ? rob_uop_6_prs2_busy : _GEN_8090; // @[rob.scala 411:{25,25}]
  wire  _GEN_8092 = 5'h7 == com_idx ? rob_uop_7_prs2_busy : _GEN_8091; // @[rob.scala 411:{25,25}]
  wire  _GEN_8093 = 5'h8 == com_idx ? rob_uop_8_prs2_busy : _GEN_8092; // @[rob.scala 411:{25,25}]
  wire  _GEN_8094 = 5'h9 == com_idx ? rob_uop_9_prs2_busy : _GEN_8093; // @[rob.scala 411:{25,25}]
  wire  _GEN_8095 = 5'ha == com_idx ? rob_uop_10_prs2_busy : _GEN_8094; // @[rob.scala 411:{25,25}]
  wire  _GEN_8096 = 5'hb == com_idx ? rob_uop_11_prs2_busy : _GEN_8095; // @[rob.scala 411:{25,25}]
  wire  _GEN_8097 = 5'hc == com_idx ? rob_uop_12_prs2_busy : _GEN_8096; // @[rob.scala 411:{25,25}]
  wire  _GEN_8098 = 5'hd == com_idx ? rob_uop_13_prs2_busy : _GEN_8097; // @[rob.scala 411:{25,25}]
  wire  _GEN_8099 = 5'he == com_idx ? rob_uop_14_prs2_busy : _GEN_8098; // @[rob.scala 411:{25,25}]
  wire  _GEN_8100 = 5'hf == com_idx ? rob_uop_15_prs2_busy : _GEN_8099; // @[rob.scala 411:{25,25}]
  wire  _GEN_8101 = 5'h10 == com_idx ? rob_uop_16_prs2_busy : _GEN_8100; // @[rob.scala 411:{25,25}]
  wire  _GEN_8102 = 5'h11 == com_idx ? rob_uop_17_prs2_busy : _GEN_8101; // @[rob.scala 411:{25,25}]
  wire  _GEN_8103 = 5'h12 == com_idx ? rob_uop_18_prs2_busy : _GEN_8102; // @[rob.scala 411:{25,25}]
  wire  _GEN_8104 = 5'h13 == com_idx ? rob_uop_19_prs2_busy : _GEN_8103; // @[rob.scala 411:{25,25}]
  wire  _GEN_8105 = 5'h14 == com_idx ? rob_uop_20_prs2_busy : _GEN_8104; // @[rob.scala 411:{25,25}]
  wire  _GEN_8106 = 5'h15 == com_idx ? rob_uop_21_prs2_busy : _GEN_8105; // @[rob.scala 411:{25,25}]
  wire  _GEN_8107 = 5'h16 == com_idx ? rob_uop_22_prs2_busy : _GEN_8106; // @[rob.scala 411:{25,25}]
  wire  _GEN_8108 = 5'h17 == com_idx ? rob_uop_23_prs2_busy : _GEN_8107; // @[rob.scala 411:{25,25}]
  wire  _GEN_8109 = 5'h18 == com_idx ? rob_uop_24_prs2_busy : _GEN_8108; // @[rob.scala 411:{25,25}]
  wire  _GEN_8110 = 5'h19 == com_idx ? rob_uop_25_prs2_busy : _GEN_8109; // @[rob.scala 411:{25,25}]
  wire  _GEN_8111 = 5'h1a == com_idx ? rob_uop_26_prs2_busy : _GEN_8110; // @[rob.scala 411:{25,25}]
  wire  _GEN_8112 = 5'h1b == com_idx ? rob_uop_27_prs2_busy : _GEN_8111; // @[rob.scala 411:{25,25}]
  wire  _GEN_8113 = 5'h1c == com_idx ? rob_uop_28_prs2_busy : _GEN_8112; // @[rob.scala 411:{25,25}]
  wire  _GEN_8114 = 5'h1d == com_idx ? rob_uop_29_prs2_busy : _GEN_8113; // @[rob.scala 411:{25,25}]
  wire  _GEN_8115 = 5'h1e == com_idx ? rob_uop_30_prs2_busy : _GEN_8114; // @[rob.scala 411:{25,25}]
  wire  _GEN_8118 = 5'h1 == com_idx ? rob_uop_1_prs1_busy : rob_uop_0_prs1_busy; // @[rob.scala 411:{25,25}]
  wire  _GEN_8119 = 5'h2 == com_idx ? rob_uop_2_prs1_busy : _GEN_8118; // @[rob.scala 411:{25,25}]
  wire  _GEN_8120 = 5'h3 == com_idx ? rob_uop_3_prs1_busy : _GEN_8119; // @[rob.scala 411:{25,25}]
  wire  _GEN_8121 = 5'h4 == com_idx ? rob_uop_4_prs1_busy : _GEN_8120; // @[rob.scala 411:{25,25}]
  wire  _GEN_8122 = 5'h5 == com_idx ? rob_uop_5_prs1_busy : _GEN_8121; // @[rob.scala 411:{25,25}]
  wire  _GEN_8123 = 5'h6 == com_idx ? rob_uop_6_prs1_busy : _GEN_8122; // @[rob.scala 411:{25,25}]
  wire  _GEN_8124 = 5'h7 == com_idx ? rob_uop_7_prs1_busy : _GEN_8123; // @[rob.scala 411:{25,25}]
  wire  _GEN_8125 = 5'h8 == com_idx ? rob_uop_8_prs1_busy : _GEN_8124; // @[rob.scala 411:{25,25}]
  wire  _GEN_8126 = 5'h9 == com_idx ? rob_uop_9_prs1_busy : _GEN_8125; // @[rob.scala 411:{25,25}]
  wire  _GEN_8127 = 5'ha == com_idx ? rob_uop_10_prs1_busy : _GEN_8126; // @[rob.scala 411:{25,25}]
  wire  _GEN_8128 = 5'hb == com_idx ? rob_uop_11_prs1_busy : _GEN_8127; // @[rob.scala 411:{25,25}]
  wire  _GEN_8129 = 5'hc == com_idx ? rob_uop_12_prs1_busy : _GEN_8128; // @[rob.scala 411:{25,25}]
  wire  _GEN_8130 = 5'hd == com_idx ? rob_uop_13_prs1_busy : _GEN_8129; // @[rob.scala 411:{25,25}]
  wire  _GEN_8131 = 5'he == com_idx ? rob_uop_14_prs1_busy : _GEN_8130; // @[rob.scala 411:{25,25}]
  wire  _GEN_8132 = 5'hf == com_idx ? rob_uop_15_prs1_busy : _GEN_8131; // @[rob.scala 411:{25,25}]
  wire  _GEN_8133 = 5'h10 == com_idx ? rob_uop_16_prs1_busy : _GEN_8132; // @[rob.scala 411:{25,25}]
  wire  _GEN_8134 = 5'h11 == com_idx ? rob_uop_17_prs1_busy : _GEN_8133; // @[rob.scala 411:{25,25}]
  wire  _GEN_8135 = 5'h12 == com_idx ? rob_uop_18_prs1_busy : _GEN_8134; // @[rob.scala 411:{25,25}]
  wire  _GEN_8136 = 5'h13 == com_idx ? rob_uop_19_prs1_busy : _GEN_8135; // @[rob.scala 411:{25,25}]
  wire  _GEN_8137 = 5'h14 == com_idx ? rob_uop_20_prs1_busy : _GEN_8136; // @[rob.scala 411:{25,25}]
  wire  _GEN_8138 = 5'h15 == com_idx ? rob_uop_21_prs1_busy : _GEN_8137; // @[rob.scala 411:{25,25}]
  wire  _GEN_8139 = 5'h16 == com_idx ? rob_uop_22_prs1_busy : _GEN_8138; // @[rob.scala 411:{25,25}]
  wire  _GEN_8140 = 5'h17 == com_idx ? rob_uop_23_prs1_busy : _GEN_8139; // @[rob.scala 411:{25,25}]
  wire  _GEN_8141 = 5'h18 == com_idx ? rob_uop_24_prs1_busy : _GEN_8140; // @[rob.scala 411:{25,25}]
  wire  _GEN_8142 = 5'h19 == com_idx ? rob_uop_25_prs1_busy : _GEN_8141; // @[rob.scala 411:{25,25}]
  wire  _GEN_8143 = 5'h1a == com_idx ? rob_uop_26_prs1_busy : _GEN_8142; // @[rob.scala 411:{25,25}]
  wire  _GEN_8144 = 5'h1b == com_idx ? rob_uop_27_prs1_busy : _GEN_8143; // @[rob.scala 411:{25,25}]
  wire  _GEN_8145 = 5'h1c == com_idx ? rob_uop_28_prs1_busy : _GEN_8144; // @[rob.scala 411:{25,25}]
  wire  _GEN_8146 = 5'h1d == com_idx ? rob_uop_29_prs1_busy : _GEN_8145; // @[rob.scala 411:{25,25}]
  wire  _GEN_8147 = 5'h1e == com_idx ? rob_uop_30_prs1_busy : _GEN_8146; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8150 = 5'h1 == com_idx ? rob_uop_1_ppred : rob_uop_0_ppred; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8151 = 5'h2 == com_idx ? rob_uop_2_ppred : _GEN_8150; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8152 = 5'h3 == com_idx ? rob_uop_3_ppred : _GEN_8151; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8153 = 5'h4 == com_idx ? rob_uop_4_ppred : _GEN_8152; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8154 = 5'h5 == com_idx ? rob_uop_5_ppred : _GEN_8153; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8155 = 5'h6 == com_idx ? rob_uop_6_ppred : _GEN_8154; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8156 = 5'h7 == com_idx ? rob_uop_7_ppred : _GEN_8155; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8157 = 5'h8 == com_idx ? rob_uop_8_ppred : _GEN_8156; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8158 = 5'h9 == com_idx ? rob_uop_9_ppred : _GEN_8157; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8159 = 5'ha == com_idx ? rob_uop_10_ppred : _GEN_8158; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8160 = 5'hb == com_idx ? rob_uop_11_ppred : _GEN_8159; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8161 = 5'hc == com_idx ? rob_uop_12_ppred : _GEN_8160; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8162 = 5'hd == com_idx ? rob_uop_13_ppred : _GEN_8161; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8163 = 5'he == com_idx ? rob_uop_14_ppred : _GEN_8162; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8164 = 5'hf == com_idx ? rob_uop_15_ppred : _GEN_8163; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8165 = 5'h10 == com_idx ? rob_uop_16_ppred : _GEN_8164; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8166 = 5'h11 == com_idx ? rob_uop_17_ppred : _GEN_8165; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8167 = 5'h12 == com_idx ? rob_uop_18_ppred : _GEN_8166; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8168 = 5'h13 == com_idx ? rob_uop_19_ppred : _GEN_8167; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8169 = 5'h14 == com_idx ? rob_uop_20_ppred : _GEN_8168; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8170 = 5'h15 == com_idx ? rob_uop_21_ppred : _GEN_8169; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8171 = 5'h16 == com_idx ? rob_uop_22_ppred : _GEN_8170; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8172 = 5'h17 == com_idx ? rob_uop_23_ppred : _GEN_8171; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8173 = 5'h18 == com_idx ? rob_uop_24_ppred : _GEN_8172; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8174 = 5'h19 == com_idx ? rob_uop_25_ppred : _GEN_8173; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8175 = 5'h1a == com_idx ? rob_uop_26_ppred : _GEN_8174; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8176 = 5'h1b == com_idx ? rob_uop_27_ppred : _GEN_8175; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8177 = 5'h1c == com_idx ? rob_uop_28_ppred : _GEN_8176; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8178 = 5'h1d == com_idx ? rob_uop_29_ppred : _GEN_8177; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8179 = 5'h1e == com_idx ? rob_uop_30_ppred : _GEN_8178; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8182 = 5'h1 == com_idx ? rob_uop_1_prs3 : rob_uop_0_prs3; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8183 = 5'h2 == com_idx ? rob_uop_2_prs3 : _GEN_8182; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8184 = 5'h3 == com_idx ? rob_uop_3_prs3 : _GEN_8183; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8185 = 5'h4 == com_idx ? rob_uop_4_prs3 : _GEN_8184; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8186 = 5'h5 == com_idx ? rob_uop_5_prs3 : _GEN_8185; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8187 = 5'h6 == com_idx ? rob_uop_6_prs3 : _GEN_8186; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8188 = 5'h7 == com_idx ? rob_uop_7_prs3 : _GEN_8187; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8189 = 5'h8 == com_idx ? rob_uop_8_prs3 : _GEN_8188; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8190 = 5'h9 == com_idx ? rob_uop_9_prs3 : _GEN_8189; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8191 = 5'ha == com_idx ? rob_uop_10_prs3 : _GEN_8190; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8192 = 5'hb == com_idx ? rob_uop_11_prs3 : _GEN_8191; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8193 = 5'hc == com_idx ? rob_uop_12_prs3 : _GEN_8192; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8194 = 5'hd == com_idx ? rob_uop_13_prs3 : _GEN_8193; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8195 = 5'he == com_idx ? rob_uop_14_prs3 : _GEN_8194; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8196 = 5'hf == com_idx ? rob_uop_15_prs3 : _GEN_8195; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8197 = 5'h10 == com_idx ? rob_uop_16_prs3 : _GEN_8196; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8198 = 5'h11 == com_idx ? rob_uop_17_prs3 : _GEN_8197; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8199 = 5'h12 == com_idx ? rob_uop_18_prs3 : _GEN_8198; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8200 = 5'h13 == com_idx ? rob_uop_19_prs3 : _GEN_8199; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8201 = 5'h14 == com_idx ? rob_uop_20_prs3 : _GEN_8200; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8202 = 5'h15 == com_idx ? rob_uop_21_prs3 : _GEN_8201; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8203 = 5'h16 == com_idx ? rob_uop_22_prs3 : _GEN_8202; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8204 = 5'h17 == com_idx ? rob_uop_23_prs3 : _GEN_8203; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8205 = 5'h18 == com_idx ? rob_uop_24_prs3 : _GEN_8204; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8206 = 5'h19 == com_idx ? rob_uop_25_prs3 : _GEN_8205; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8207 = 5'h1a == com_idx ? rob_uop_26_prs3 : _GEN_8206; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8208 = 5'h1b == com_idx ? rob_uop_27_prs3 : _GEN_8207; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8209 = 5'h1c == com_idx ? rob_uop_28_prs3 : _GEN_8208; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8210 = 5'h1d == com_idx ? rob_uop_29_prs3 : _GEN_8209; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8211 = 5'h1e == com_idx ? rob_uop_30_prs3 : _GEN_8210; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8214 = 5'h1 == com_idx ? rob_uop_1_prs2 : rob_uop_0_prs2; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8215 = 5'h2 == com_idx ? rob_uop_2_prs2 : _GEN_8214; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8216 = 5'h3 == com_idx ? rob_uop_3_prs2 : _GEN_8215; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8217 = 5'h4 == com_idx ? rob_uop_4_prs2 : _GEN_8216; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8218 = 5'h5 == com_idx ? rob_uop_5_prs2 : _GEN_8217; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8219 = 5'h6 == com_idx ? rob_uop_6_prs2 : _GEN_8218; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8220 = 5'h7 == com_idx ? rob_uop_7_prs2 : _GEN_8219; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8221 = 5'h8 == com_idx ? rob_uop_8_prs2 : _GEN_8220; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8222 = 5'h9 == com_idx ? rob_uop_9_prs2 : _GEN_8221; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8223 = 5'ha == com_idx ? rob_uop_10_prs2 : _GEN_8222; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8224 = 5'hb == com_idx ? rob_uop_11_prs2 : _GEN_8223; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8225 = 5'hc == com_idx ? rob_uop_12_prs2 : _GEN_8224; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8226 = 5'hd == com_idx ? rob_uop_13_prs2 : _GEN_8225; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8227 = 5'he == com_idx ? rob_uop_14_prs2 : _GEN_8226; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8228 = 5'hf == com_idx ? rob_uop_15_prs2 : _GEN_8227; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8229 = 5'h10 == com_idx ? rob_uop_16_prs2 : _GEN_8228; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8230 = 5'h11 == com_idx ? rob_uop_17_prs2 : _GEN_8229; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8231 = 5'h12 == com_idx ? rob_uop_18_prs2 : _GEN_8230; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8232 = 5'h13 == com_idx ? rob_uop_19_prs2 : _GEN_8231; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8233 = 5'h14 == com_idx ? rob_uop_20_prs2 : _GEN_8232; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8234 = 5'h15 == com_idx ? rob_uop_21_prs2 : _GEN_8233; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8235 = 5'h16 == com_idx ? rob_uop_22_prs2 : _GEN_8234; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8236 = 5'h17 == com_idx ? rob_uop_23_prs2 : _GEN_8235; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8237 = 5'h18 == com_idx ? rob_uop_24_prs2 : _GEN_8236; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8238 = 5'h19 == com_idx ? rob_uop_25_prs2 : _GEN_8237; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8239 = 5'h1a == com_idx ? rob_uop_26_prs2 : _GEN_8238; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8240 = 5'h1b == com_idx ? rob_uop_27_prs2 : _GEN_8239; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8241 = 5'h1c == com_idx ? rob_uop_28_prs2 : _GEN_8240; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8242 = 5'h1d == com_idx ? rob_uop_29_prs2 : _GEN_8241; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8243 = 5'h1e == com_idx ? rob_uop_30_prs2 : _GEN_8242; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8246 = 5'h1 == com_idx ? rob_uop_1_prs1 : rob_uop_0_prs1; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8247 = 5'h2 == com_idx ? rob_uop_2_prs1 : _GEN_8246; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8248 = 5'h3 == com_idx ? rob_uop_3_prs1 : _GEN_8247; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8249 = 5'h4 == com_idx ? rob_uop_4_prs1 : _GEN_8248; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8250 = 5'h5 == com_idx ? rob_uop_5_prs1 : _GEN_8249; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8251 = 5'h6 == com_idx ? rob_uop_6_prs1 : _GEN_8250; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8252 = 5'h7 == com_idx ? rob_uop_7_prs1 : _GEN_8251; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8253 = 5'h8 == com_idx ? rob_uop_8_prs1 : _GEN_8252; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8254 = 5'h9 == com_idx ? rob_uop_9_prs1 : _GEN_8253; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8255 = 5'ha == com_idx ? rob_uop_10_prs1 : _GEN_8254; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8256 = 5'hb == com_idx ? rob_uop_11_prs1 : _GEN_8255; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8257 = 5'hc == com_idx ? rob_uop_12_prs1 : _GEN_8256; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8258 = 5'hd == com_idx ? rob_uop_13_prs1 : _GEN_8257; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8259 = 5'he == com_idx ? rob_uop_14_prs1 : _GEN_8258; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8260 = 5'hf == com_idx ? rob_uop_15_prs1 : _GEN_8259; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8261 = 5'h10 == com_idx ? rob_uop_16_prs1 : _GEN_8260; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8262 = 5'h11 == com_idx ? rob_uop_17_prs1 : _GEN_8261; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8263 = 5'h12 == com_idx ? rob_uop_18_prs1 : _GEN_8262; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8264 = 5'h13 == com_idx ? rob_uop_19_prs1 : _GEN_8263; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8265 = 5'h14 == com_idx ? rob_uop_20_prs1 : _GEN_8264; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8266 = 5'h15 == com_idx ? rob_uop_21_prs1 : _GEN_8265; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8267 = 5'h16 == com_idx ? rob_uop_22_prs1 : _GEN_8266; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8268 = 5'h17 == com_idx ? rob_uop_23_prs1 : _GEN_8267; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8269 = 5'h18 == com_idx ? rob_uop_24_prs1 : _GEN_8268; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8270 = 5'h19 == com_idx ? rob_uop_25_prs1 : _GEN_8269; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8271 = 5'h1a == com_idx ? rob_uop_26_prs1 : _GEN_8270; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8272 = 5'h1b == com_idx ? rob_uop_27_prs1 : _GEN_8271; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8273 = 5'h1c == com_idx ? rob_uop_28_prs1 : _GEN_8272; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8274 = 5'h1d == com_idx ? rob_uop_29_prs1 : _GEN_8273; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8275 = 5'h1e == com_idx ? rob_uop_30_prs1 : _GEN_8274; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8278 = 5'h1 == com_idx ? rob_uop_1_pdst : rob_uop_0_pdst; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8279 = 5'h2 == com_idx ? rob_uop_2_pdst : _GEN_8278; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8280 = 5'h3 == com_idx ? rob_uop_3_pdst : _GEN_8279; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8281 = 5'h4 == com_idx ? rob_uop_4_pdst : _GEN_8280; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8282 = 5'h5 == com_idx ? rob_uop_5_pdst : _GEN_8281; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8283 = 5'h6 == com_idx ? rob_uop_6_pdst : _GEN_8282; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8284 = 5'h7 == com_idx ? rob_uop_7_pdst : _GEN_8283; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8285 = 5'h8 == com_idx ? rob_uop_8_pdst : _GEN_8284; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8286 = 5'h9 == com_idx ? rob_uop_9_pdst : _GEN_8285; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8287 = 5'ha == com_idx ? rob_uop_10_pdst : _GEN_8286; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8288 = 5'hb == com_idx ? rob_uop_11_pdst : _GEN_8287; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8289 = 5'hc == com_idx ? rob_uop_12_pdst : _GEN_8288; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8290 = 5'hd == com_idx ? rob_uop_13_pdst : _GEN_8289; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8291 = 5'he == com_idx ? rob_uop_14_pdst : _GEN_8290; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8292 = 5'hf == com_idx ? rob_uop_15_pdst : _GEN_8291; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8293 = 5'h10 == com_idx ? rob_uop_16_pdst : _GEN_8292; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8294 = 5'h11 == com_idx ? rob_uop_17_pdst : _GEN_8293; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8295 = 5'h12 == com_idx ? rob_uop_18_pdst : _GEN_8294; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8296 = 5'h13 == com_idx ? rob_uop_19_pdst : _GEN_8295; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8297 = 5'h14 == com_idx ? rob_uop_20_pdst : _GEN_8296; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8298 = 5'h15 == com_idx ? rob_uop_21_pdst : _GEN_8297; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8299 = 5'h16 == com_idx ? rob_uop_22_pdst : _GEN_8298; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8300 = 5'h17 == com_idx ? rob_uop_23_pdst : _GEN_8299; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8301 = 5'h18 == com_idx ? rob_uop_24_pdst : _GEN_8300; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8302 = 5'h19 == com_idx ? rob_uop_25_pdst : _GEN_8301; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8303 = 5'h1a == com_idx ? rob_uop_26_pdst : _GEN_8302; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8304 = 5'h1b == com_idx ? rob_uop_27_pdst : _GEN_8303; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8305 = 5'h1c == com_idx ? rob_uop_28_pdst : _GEN_8304; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8306 = 5'h1d == com_idx ? rob_uop_29_pdst : _GEN_8305; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8307 = 5'h1e == com_idx ? rob_uop_30_pdst : _GEN_8306; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8310 = 5'h1 == com_idx ? rob_uop_1_rxq_idx : rob_uop_0_rxq_idx; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8311 = 5'h2 == com_idx ? rob_uop_2_rxq_idx : _GEN_8310; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8312 = 5'h3 == com_idx ? rob_uop_3_rxq_idx : _GEN_8311; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8313 = 5'h4 == com_idx ? rob_uop_4_rxq_idx : _GEN_8312; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8314 = 5'h5 == com_idx ? rob_uop_5_rxq_idx : _GEN_8313; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8315 = 5'h6 == com_idx ? rob_uop_6_rxq_idx : _GEN_8314; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8316 = 5'h7 == com_idx ? rob_uop_7_rxq_idx : _GEN_8315; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8317 = 5'h8 == com_idx ? rob_uop_8_rxq_idx : _GEN_8316; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8318 = 5'h9 == com_idx ? rob_uop_9_rxq_idx : _GEN_8317; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8319 = 5'ha == com_idx ? rob_uop_10_rxq_idx : _GEN_8318; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8320 = 5'hb == com_idx ? rob_uop_11_rxq_idx : _GEN_8319; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8321 = 5'hc == com_idx ? rob_uop_12_rxq_idx : _GEN_8320; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8322 = 5'hd == com_idx ? rob_uop_13_rxq_idx : _GEN_8321; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8323 = 5'he == com_idx ? rob_uop_14_rxq_idx : _GEN_8322; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8324 = 5'hf == com_idx ? rob_uop_15_rxq_idx : _GEN_8323; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8325 = 5'h10 == com_idx ? rob_uop_16_rxq_idx : _GEN_8324; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8326 = 5'h11 == com_idx ? rob_uop_17_rxq_idx : _GEN_8325; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8327 = 5'h12 == com_idx ? rob_uop_18_rxq_idx : _GEN_8326; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8328 = 5'h13 == com_idx ? rob_uop_19_rxq_idx : _GEN_8327; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8329 = 5'h14 == com_idx ? rob_uop_20_rxq_idx : _GEN_8328; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8330 = 5'h15 == com_idx ? rob_uop_21_rxq_idx : _GEN_8329; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8331 = 5'h16 == com_idx ? rob_uop_22_rxq_idx : _GEN_8330; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8332 = 5'h17 == com_idx ? rob_uop_23_rxq_idx : _GEN_8331; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8333 = 5'h18 == com_idx ? rob_uop_24_rxq_idx : _GEN_8332; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8334 = 5'h19 == com_idx ? rob_uop_25_rxq_idx : _GEN_8333; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8335 = 5'h1a == com_idx ? rob_uop_26_rxq_idx : _GEN_8334; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8336 = 5'h1b == com_idx ? rob_uop_27_rxq_idx : _GEN_8335; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8337 = 5'h1c == com_idx ? rob_uop_28_rxq_idx : _GEN_8336; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8338 = 5'h1d == com_idx ? rob_uop_29_rxq_idx : _GEN_8337; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8339 = 5'h1e == com_idx ? rob_uop_30_rxq_idx : _GEN_8338; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8342 = 5'h1 == com_idx ? rob_uop_1_stq_idx : rob_uop_0_stq_idx; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8343 = 5'h2 == com_idx ? rob_uop_2_stq_idx : _GEN_8342; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8344 = 5'h3 == com_idx ? rob_uop_3_stq_idx : _GEN_8343; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8345 = 5'h4 == com_idx ? rob_uop_4_stq_idx : _GEN_8344; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8346 = 5'h5 == com_idx ? rob_uop_5_stq_idx : _GEN_8345; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8347 = 5'h6 == com_idx ? rob_uop_6_stq_idx : _GEN_8346; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8348 = 5'h7 == com_idx ? rob_uop_7_stq_idx : _GEN_8347; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8349 = 5'h8 == com_idx ? rob_uop_8_stq_idx : _GEN_8348; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8350 = 5'h9 == com_idx ? rob_uop_9_stq_idx : _GEN_8349; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8351 = 5'ha == com_idx ? rob_uop_10_stq_idx : _GEN_8350; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8352 = 5'hb == com_idx ? rob_uop_11_stq_idx : _GEN_8351; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8353 = 5'hc == com_idx ? rob_uop_12_stq_idx : _GEN_8352; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8354 = 5'hd == com_idx ? rob_uop_13_stq_idx : _GEN_8353; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8355 = 5'he == com_idx ? rob_uop_14_stq_idx : _GEN_8354; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8356 = 5'hf == com_idx ? rob_uop_15_stq_idx : _GEN_8355; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8357 = 5'h10 == com_idx ? rob_uop_16_stq_idx : _GEN_8356; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8358 = 5'h11 == com_idx ? rob_uop_17_stq_idx : _GEN_8357; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8359 = 5'h12 == com_idx ? rob_uop_18_stq_idx : _GEN_8358; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8360 = 5'h13 == com_idx ? rob_uop_19_stq_idx : _GEN_8359; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8361 = 5'h14 == com_idx ? rob_uop_20_stq_idx : _GEN_8360; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8362 = 5'h15 == com_idx ? rob_uop_21_stq_idx : _GEN_8361; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8363 = 5'h16 == com_idx ? rob_uop_22_stq_idx : _GEN_8362; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8364 = 5'h17 == com_idx ? rob_uop_23_stq_idx : _GEN_8363; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8365 = 5'h18 == com_idx ? rob_uop_24_stq_idx : _GEN_8364; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8366 = 5'h19 == com_idx ? rob_uop_25_stq_idx : _GEN_8365; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8367 = 5'h1a == com_idx ? rob_uop_26_stq_idx : _GEN_8366; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8368 = 5'h1b == com_idx ? rob_uop_27_stq_idx : _GEN_8367; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8369 = 5'h1c == com_idx ? rob_uop_28_stq_idx : _GEN_8368; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8370 = 5'h1d == com_idx ? rob_uop_29_stq_idx : _GEN_8369; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8371 = 5'h1e == com_idx ? rob_uop_30_stq_idx : _GEN_8370; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8374 = 5'h1 == com_idx ? rob_uop_1_ldq_idx : rob_uop_0_ldq_idx; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8375 = 5'h2 == com_idx ? rob_uop_2_ldq_idx : _GEN_8374; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8376 = 5'h3 == com_idx ? rob_uop_3_ldq_idx : _GEN_8375; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8377 = 5'h4 == com_idx ? rob_uop_4_ldq_idx : _GEN_8376; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8378 = 5'h5 == com_idx ? rob_uop_5_ldq_idx : _GEN_8377; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8379 = 5'h6 == com_idx ? rob_uop_6_ldq_idx : _GEN_8378; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8380 = 5'h7 == com_idx ? rob_uop_7_ldq_idx : _GEN_8379; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8381 = 5'h8 == com_idx ? rob_uop_8_ldq_idx : _GEN_8380; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8382 = 5'h9 == com_idx ? rob_uop_9_ldq_idx : _GEN_8381; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8383 = 5'ha == com_idx ? rob_uop_10_ldq_idx : _GEN_8382; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8384 = 5'hb == com_idx ? rob_uop_11_ldq_idx : _GEN_8383; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8385 = 5'hc == com_idx ? rob_uop_12_ldq_idx : _GEN_8384; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8386 = 5'hd == com_idx ? rob_uop_13_ldq_idx : _GEN_8385; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8387 = 5'he == com_idx ? rob_uop_14_ldq_idx : _GEN_8386; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8388 = 5'hf == com_idx ? rob_uop_15_ldq_idx : _GEN_8387; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8389 = 5'h10 == com_idx ? rob_uop_16_ldq_idx : _GEN_8388; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8390 = 5'h11 == com_idx ? rob_uop_17_ldq_idx : _GEN_8389; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8391 = 5'h12 == com_idx ? rob_uop_18_ldq_idx : _GEN_8390; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8392 = 5'h13 == com_idx ? rob_uop_19_ldq_idx : _GEN_8391; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8393 = 5'h14 == com_idx ? rob_uop_20_ldq_idx : _GEN_8392; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8394 = 5'h15 == com_idx ? rob_uop_21_ldq_idx : _GEN_8393; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8395 = 5'h16 == com_idx ? rob_uop_22_ldq_idx : _GEN_8394; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8396 = 5'h17 == com_idx ? rob_uop_23_ldq_idx : _GEN_8395; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8397 = 5'h18 == com_idx ? rob_uop_24_ldq_idx : _GEN_8396; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8398 = 5'h19 == com_idx ? rob_uop_25_ldq_idx : _GEN_8397; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8399 = 5'h1a == com_idx ? rob_uop_26_ldq_idx : _GEN_8398; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8400 = 5'h1b == com_idx ? rob_uop_27_ldq_idx : _GEN_8399; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8401 = 5'h1c == com_idx ? rob_uop_28_ldq_idx : _GEN_8400; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8402 = 5'h1d == com_idx ? rob_uop_29_ldq_idx : _GEN_8401; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8403 = 5'h1e == com_idx ? rob_uop_30_ldq_idx : _GEN_8402; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8406 = 5'h1 == com_idx ? rob_uop_1_rob_idx : rob_uop_0_rob_idx; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8407 = 5'h2 == com_idx ? rob_uop_2_rob_idx : _GEN_8406; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8408 = 5'h3 == com_idx ? rob_uop_3_rob_idx : _GEN_8407; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8409 = 5'h4 == com_idx ? rob_uop_4_rob_idx : _GEN_8408; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8410 = 5'h5 == com_idx ? rob_uop_5_rob_idx : _GEN_8409; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8411 = 5'h6 == com_idx ? rob_uop_6_rob_idx : _GEN_8410; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8412 = 5'h7 == com_idx ? rob_uop_7_rob_idx : _GEN_8411; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8413 = 5'h8 == com_idx ? rob_uop_8_rob_idx : _GEN_8412; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8414 = 5'h9 == com_idx ? rob_uop_9_rob_idx : _GEN_8413; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8415 = 5'ha == com_idx ? rob_uop_10_rob_idx : _GEN_8414; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8416 = 5'hb == com_idx ? rob_uop_11_rob_idx : _GEN_8415; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8417 = 5'hc == com_idx ? rob_uop_12_rob_idx : _GEN_8416; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8418 = 5'hd == com_idx ? rob_uop_13_rob_idx : _GEN_8417; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8419 = 5'he == com_idx ? rob_uop_14_rob_idx : _GEN_8418; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8420 = 5'hf == com_idx ? rob_uop_15_rob_idx : _GEN_8419; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8421 = 5'h10 == com_idx ? rob_uop_16_rob_idx : _GEN_8420; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8422 = 5'h11 == com_idx ? rob_uop_17_rob_idx : _GEN_8421; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8423 = 5'h12 == com_idx ? rob_uop_18_rob_idx : _GEN_8422; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8424 = 5'h13 == com_idx ? rob_uop_19_rob_idx : _GEN_8423; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8425 = 5'h14 == com_idx ? rob_uop_20_rob_idx : _GEN_8424; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8426 = 5'h15 == com_idx ? rob_uop_21_rob_idx : _GEN_8425; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8427 = 5'h16 == com_idx ? rob_uop_22_rob_idx : _GEN_8426; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8428 = 5'h17 == com_idx ? rob_uop_23_rob_idx : _GEN_8427; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8429 = 5'h18 == com_idx ? rob_uop_24_rob_idx : _GEN_8428; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8430 = 5'h19 == com_idx ? rob_uop_25_rob_idx : _GEN_8429; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8431 = 5'h1a == com_idx ? rob_uop_26_rob_idx : _GEN_8430; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8432 = 5'h1b == com_idx ? rob_uop_27_rob_idx : _GEN_8431; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8433 = 5'h1c == com_idx ? rob_uop_28_rob_idx : _GEN_8432; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8434 = 5'h1d == com_idx ? rob_uop_29_rob_idx : _GEN_8433; // @[rob.scala 411:{25,25}]
  wire [4:0] _GEN_8435 = 5'h1e == com_idx ? rob_uop_30_rob_idx : _GEN_8434; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8438 = 5'h1 == com_idx ? rob_uop_1_csr_addr : rob_uop_0_csr_addr; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8439 = 5'h2 == com_idx ? rob_uop_2_csr_addr : _GEN_8438; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8440 = 5'h3 == com_idx ? rob_uop_3_csr_addr : _GEN_8439; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8441 = 5'h4 == com_idx ? rob_uop_4_csr_addr : _GEN_8440; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8442 = 5'h5 == com_idx ? rob_uop_5_csr_addr : _GEN_8441; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8443 = 5'h6 == com_idx ? rob_uop_6_csr_addr : _GEN_8442; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8444 = 5'h7 == com_idx ? rob_uop_7_csr_addr : _GEN_8443; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8445 = 5'h8 == com_idx ? rob_uop_8_csr_addr : _GEN_8444; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8446 = 5'h9 == com_idx ? rob_uop_9_csr_addr : _GEN_8445; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8447 = 5'ha == com_idx ? rob_uop_10_csr_addr : _GEN_8446; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8448 = 5'hb == com_idx ? rob_uop_11_csr_addr : _GEN_8447; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8449 = 5'hc == com_idx ? rob_uop_12_csr_addr : _GEN_8448; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8450 = 5'hd == com_idx ? rob_uop_13_csr_addr : _GEN_8449; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8451 = 5'he == com_idx ? rob_uop_14_csr_addr : _GEN_8450; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8452 = 5'hf == com_idx ? rob_uop_15_csr_addr : _GEN_8451; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8453 = 5'h10 == com_idx ? rob_uop_16_csr_addr : _GEN_8452; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8454 = 5'h11 == com_idx ? rob_uop_17_csr_addr : _GEN_8453; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8455 = 5'h12 == com_idx ? rob_uop_18_csr_addr : _GEN_8454; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8456 = 5'h13 == com_idx ? rob_uop_19_csr_addr : _GEN_8455; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8457 = 5'h14 == com_idx ? rob_uop_20_csr_addr : _GEN_8456; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8458 = 5'h15 == com_idx ? rob_uop_21_csr_addr : _GEN_8457; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8459 = 5'h16 == com_idx ? rob_uop_22_csr_addr : _GEN_8458; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8460 = 5'h17 == com_idx ? rob_uop_23_csr_addr : _GEN_8459; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8461 = 5'h18 == com_idx ? rob_uop_24_csr_addr : _GEN_8460; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8462 = 5'h19 == com_idx ? rob_uop_25_csr_addr : _GEN_8461; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8463 = 5'h1a == com_idx ? rob_uop_26_csr_addr : _GEN_8462; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8464 = 5'h1b == com_idx ? rob_uop_27_csr_addr : _GEN_8463; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8465 = 5'h1c == com_idx ? rob_uop_28_csr_addr : _GEN_8464; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8466 = 5'h1d == com_idx ? rob_uop_29_csr_addr : _GEN_8465; // @[rob.scala 411:{25,25}]
  wire [11:0] _GEN_8467 = 5'h1e == com_idx ? rob_uop_30_csr_addr : _GEN_8466; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8470 = 5'h1 == com_idx ? rob_uop_1_imm_packed : rob_uop_0_imm_packed; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8471 = 5'h2 == com_idx ? rob_uop_2_imm_packed : _GEN_8470; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8472 = 5'h3 == com_idx ? rob_uop_3_imm_packed : _GEN_8471; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8473 = 5'h4 == com_idx ? rob_uop_4_imm_packed : _GEN_8472; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8474 = 5'h5 == com_idx ? rob_uop_5_imm_packed : _GEN_8473; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8475 = 5'h6 == com_idx ? rob_uop_6_imm_packed : _GEN_8474; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8476 = 5'h7 == com_idx ? rob_uop_7_imm_packed : _GEN_8475; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8477 = 5'h8 == com_idx ? rob_uop_8_imm_packed : _GEN_8476; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8478 = 5'h9 == com_idx ? rob_uop_9_imm_packed : _GEN_8477; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8479 = 5'ha == com_idx ? rob_uop_10_imm_packed : _GEN_8478; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8480 = 5'hb == com_idx ? rob_uop_11_imm_packed : _GEN_8479; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8481 = 5'hc == com_idx ? rob_uop_12_imm_packed : _GEN_8480; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8482 = 5'hd == com_idx ? rob_uop_13_imm_packed : _GEN_8481; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8483 = 5'he == com_idx ? rob_uop_14_imm_packed : _GEN_8482; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8484 = 5'hf == com_idx ? rob_uop_15_imm_packed : _GEN_8483; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8485 = 5'h10 == com_idx ? rob_uop_16_imm_packed : _GEN_8484; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8486 = 5'h11 == com_idx ? rob_uop_17_imm_packed : _GEN_8485; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8487 = 5'h12 == com_idx ? rob_uop_18_imm_packed : _GEN_8486; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8488 = 5'h13 == com_idx ? rob_uop_19_imm_packed : _GEN_8487; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8489 = 5'h14 == com_idx ? rob_uop_20_imm_packed : _GEN_8488; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8490 = 5'h15 == com_idx ? rob_uop_21_imm_packed : _GEN_8489; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8491 = 5'h16 == com_idx ? rob_uop_22_imm_packed : _GEN_8490; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8492 = 5'h17 == com_idx ? rob_uop_23_imm_packed : _GEN_8491; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8493 = 5'h18 == com_idx ? rob_uop_24_imm_packed : _GEN_8492; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8494 = 5'h19 == com_idx ? rob_uop_25_imm_packed : _GEN_8493; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8495 = 5'h1a == com_idx ? rob_uop_26_imm_packed : _GEN_8494; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8496 = 5'h1b == com_idx ? rob_uop_27_imm_packed : _GEN_8495; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8497 = 5'h1c == com_idx ? rob_uop_28_imm_packed : _GEN_8496; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8498 = 5'h1d == com_idx ? rob_uop_29_imm_packed : _GEN_8497; // @[rob.scala 411:{25,25}]
  wire [19:0] _GEN_8499 = 5'h1e == com_idx ? rob_uop_30_imm_packed : _GEN_8498; // @[rob.scala 411:{25,25}]
  wire  _GEN_8502 = 5'h1 == com_idx ? rob_uop_1_taken : rob_uop_0_taken; // @[rob.scala 411:{25,25}]
  wire  _GEN_8503 = 5'h2 == com_idx ? rob_uop_2_taken : _GEN_8502; // @[rob.scala 411:{25,25}]
  wire  _GEN_8504 = 5'h3 == com_idx ? rob_uop_3_taken : _GEN_8503; // @[rob.scala 411:{25,25}]
  wire  _GEN_8505 = 5'h4 == com_idx ? rob_uop_4_taken : _GEN_8504; // @[rob.scala 411:{25,25}]
  wire  _GEN_8506 = 5'h5 == com_idx ? rob_uop_5_taken : _GEN_8505; // @[rob.scala 411:{25,25}]
  wire  _GEN_8507 = 5'h6 == com_idx ? rob_uop_6_taken : _GEN_8506; // @[rob.scala 411:{25,25}]
  wire  _GEN_8508 = 5'h7 == com_idx ? rob_uop_7_taken : _GEN_8507; // @[rob.scala 411:{25,25}]
  wire  _GEN_8509 = 5'h8 == com_idx ? rob_uop_8_taken : _GEN_8508; // @[rob.scala 411:{25,25}]
  wire  _GEN_8510 = 5'h9 == com_idx ? rob_uop_9_taken : _GEN_8509; // @[rob.scala 411:{25,25}]
  wire  _GEN_8511 = 5'ha == com_idx ? rob_uop_10_taken : _GEN_8510; // @[rob.scala 411:{25,25}]
  wire  _GEN_8512 = 5'hb == com_idx ? rob_uop_11_taken : _GEN_8511; // @[rob.scala 411:{25,25}]
  wire  _GEN_8513 = 5'hc == com_idx ? rob_uop_12_taken : _GEN_8512; // @[rob.scala 411:{25,25}]
  wire  _GEN_8514 = 5'hd == com_idx ? rob_uop_13_taken : _GEN_8513; // @[rob.scala 411:{25,25}]
  wire  _GEN_8515 = 5'he == com_idx ? rob_uop_14_taken : _GEN_8514; // @[rob.scala 411:{25,25}]
  wire  _GEN_8516 = 5'hf == com_idx ? rob_uop_15_taken : _GEN_8515; // @[rob.scala 411:{25,25}]
  wire  _GEN_8517 = 5'h10 == com_idx ? rob_uop_16_taken : _GEN_8516; // @[rob.scala 411:{25,25}]
  wire  _GEN_8518 = 5'h11 == com_idx ? rob_uop_17_taken : _GEN_8517; // @[rob.scala 411:{25,25}]
  wire  _GEN_8519 = 5'h12 == com_idx ? rob_uop_18_taken : _GEN_8518; // @[rob.scala 411:{25,25}]
  wire  _GEN_8520 = 5'h13 == com_idx ? rob_uop_19_taken : _GEN_8519; // @[rob.scala 411:{25,25}]
  wire  _GEN_8521 = 5'h14 == com_idx ? rob_uop_20_taken : _GEN_8520; // @[rob.scala 411:{25,25}]
  wire  _GEN_8522 = 5'h15 == com_idx ? rob_uop_21_taken : _GEN_8521; // @[rob.scala 411:{25,25}]
  wire  _GEN_8523 = 5'h16 == com_idx ? rob_uop_22_taken : _GEN_8522; // @[rob.scala 411:{25,25}]
  wire  _GEN_8524 = 5'h17 == com_idx ? rob_uop_23_taken : _GEN_8523; // @[rob.scala 411:{25,25}]
  wire  _GEN_8525 = 5'h18 == com_idx ? rob_uop_24_taken : _GEN_8524; // @[rob.scala 411:{25,25}]
  wire  _GEN_8526 = 5'h19 == com_idx ? rob_uop_25_taken : _GEN_8525; // @[rob.scala 411:{25,25}]
  wire  _GEN_8527 = 5'h1a == com_idx ? rob_uop_26_taken : _GEN_8526; // @[rob.scala 411:{25,25}]
  wire  _GEN_8528 = 5'h1b == com_idx ? rob_uop_27_taken : _GEN_8527; // @[rob.scala 411:{25,25}]
  wire  _GEN_8529 = 5'h1c == com_idx ? rob_uop_28_taken : _GEN_8528; // @[rob.scala 411:{25,25}]
  wire  _GEN_8530 = 5'h1d == com_idx ? rob_uop_29_taken : _GEN_8529; // @[rob.scala 411:{25,25}]
  wire  _GEN_8531 = 5'h1e == com_idx ? rob_uop_30_taken : _GEN_8530; // @[rob.scala 411:{25,25}]
  wire  _GEN_8532 = 5'h1f == com_idx ? rob_uop_31_taken : _GEN_8531; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8534 = 5'h1 == com_idx ? rob_uop_1_pc_lob : rob_uop_0_pc_lob; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8535 = 5'h2 == com_idx ? rob_uop_2_pc_lob : _GEN_8534; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8536 = 5'h3 == com_idx ? rob_uop_3_pc_lob : _GEN_8535; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8537 = 5'h4 == com_idx ? rob_uop_4_pc_lob : _GEN_8536; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8538 = 5'h5 == com_idx ? rob_uop_5_pc_lob : _GEN_8537; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8539 = 5'h6 == com_idx ? rob_uop_6_pc_lob : _GEN_8538; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8540 = 5'h7 == com_idx ? rob_uop_7_pc_lob : _GEN_8539; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8541 = 5'h8 == com_idx ? rob_uop_8_pc_lob : _GEN_8540; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8542 = 5'h9 == com_idx ? rob_uop_9_pc_lob : _GEN_8541; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8543 = 5'ha == com_idx ? rob_uop_10_pc_lob : _GEN_8542; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8544 = 5'hb == com_idx ? rob_uop_11_pc_lob : _GEN_8543; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8545 = 5'hc == com_idx ? rob_uop_12_pc_lob : _GEN_8544; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8546 = 5'hd == com_idx ? rob_uop_13_pc_lob : _GEN_8545; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8547 = 5'he == com_idx ? rob_uop_14_pc_lob : _GEN_8546; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8548 = 5'hf == com_idx ? rob_uop_15_pc_lob : _GEN_8547; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8549 = 5'h10 == com_idx ? rob_uop_16_pc_lob : _GEN_8548; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8550 = 5'h11 == com_idx ? rob_uop_17_pc_lob : _GEN_8549; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8551 = 5'h12 == com_idx ? rob_uop_18_pc_lob : _GEN_8550; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8552 = 5'h13 == com_idx ? rob_uop_19_pc_lob : _GEN_8551; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8553 = 5'h14 == com_idx ? rob_uop_20_pc_lob : _GEN_8552; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8554 = 5'h15 == com_idx ? rob_uop_21_pc_lob : _GEN_8553; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8555 = 5'h16 == com_idx ? rob_uop_22_pc_lob : _GEN_8554; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8556 = 5'h17 == com_idx ? rob_uop_23_pc_lob : _GEN_8555; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8557 = 5'h18 == com_idx ? rob_uop_24_pc_lob : _GEN_8556; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8558 = 5'h19 == com_idx ? rob_uop_25_pc_lob : _GEN_8557; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8559 = 5'h1a == com_idx ? rob_uop_26_pc_lob : _GEN_8558; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8560 = 5'h1b == com_idx ? rob_uop_27_pc_lob : _GEN_8559; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8561 = 5'h1c == com_idx ? rob_uop_28_pc_lob : _GEN_8560; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8562 = 5'h1d == com_idx ? rob_uop_29_pc_lob : _GEN_8561; // @[rob.scala 411:{25,25}]
  wire [5:0] _GEN_8563 = 5'h1e == com_idx ? rob_uop_30_pc_lob : _GEN_8562; // @[rob.scala 411:{25,25}]
  wire  _GEN_8566 = 5'h1 == com_idx ? rob_uop_1_edge_inst : rob_uop_0_edge_inst; // @[rob.scala 411:{25,25}]
  wire  _GEN_8567 = 5'h2 == com_idx ? rob_uop_2_edge_inst : _GEN_8566; // @[rob.scala 411:{25,25}]
  wire  _GEN_8568 = 5'h3 == com_idx ? rob_uop_3_edge_inst : _GEN_8567; // @[rob.scala 411:{25,25}]
  wire  _GEN_8569 = 5'h4 == com_idx ? rob_uop_4_edge_inst : _GEN_8568; // @[rob.scala 411:{25,25}]
  wire  _GEN_8570 = 5'h5 == com_idx ? rob_uop_5_edge_inst : _GEN_8569; // @[rob.scala 411:{25,25}]
  wire  _GEN_8571 = 5'h6 == com_idx ? rob_uop_6_edge_inst : _GEN_8570; // @[rob.scala 411:{25,25}]
  wire  _GEN_8572 = 5'h7 == com_idx ? rob_uop_7_edge_inst : _GEN_8571; // @[rob.scala 411:{25,25}]
  wire  _GEN_8573 = 5'h8 == com_idx ? rob_uop_8_edge_inst : _GEN_8572; // @[rob.scala 411:{25,25}]
  wire  _GEN_8574 = 5'h9 == com_idx ? rob_uop_9_edge_inst : _GEN_8573; // @[rob.scala 411:{25,25}]
  wire  _GEN_8575 = 5'ha == com_idx ? rob_uop_10_edge_inst : _GEN_8574; // @[rob.scala 411:{25,25}]
  wire  _GEN_8576 = 5'hb == com_idx ? rob_uop_11_edge_inst : _GEN_8575; // @[rob.scala 411:{25,25}]
  wire  _GEN_8577 = 5'hc == com_idx ? rob_uop_12_edge_inst : _GEN_8576; // @[rob.scala 411:{25,25}]
  wire  _GEN_8578 = 5'hd == com_idx ? rob_uop_13_edge_inst : _GEN_8577; // @[rob.scala 411:{25,25}]
  wire  _GEN_8579 = 5'he == com_idx ? rob_uop_14_edge_inst : _GEN_8578; // @[rob.scala 411:{25,25}]
  wire  _GEN_8580 = 5'hf == com_idx ? rob_uop_15_edge_inst : _GEN_8579; // @[rob.scala 411:{25,25}]
  wire  _GEN_8581 = 5'h10 == com_idx ? rob_uop_16_edge_inst : _GEN_8580; // @[rob.scala 411:{25,25}]
  wire  _GEN_8582 = 5'h11 == com_idx ? rob_uop_17_edge_inst : _GEN_8581; // @[rob.scala 411:{25,25}]
  wire  _GEN_8583 = 5'h12 == com_idx ? rob_uop_18_edge_inst : _GEN_8582; // @[rob.scala 411:{25,25}]
  wire  _GEN_8584 = 5'h13 == com_idx ? rob_uop_19_edge_inst : _GEN_8583; // @[rob.scala 411:{25,25}]
  wire  _GEN_8585 = 5'h14 == com_idx ? rob_uop_20_edge_inst : _GEN_8584; // @[rob.scala 411:{25,25}]
  wire  _GEN_8586 = 5'h15 == com_idx ? rob_uop_21_edge_inst : _GEN_8585; // @[rob.scala 411:{25,25}]
  wire  _GEN_8587 = 5'h16 == com_idx ? rob_uop_22_edge_inst : _GEN_8586; // @[rob.scala 411:{25,25}]
  wire  _GEN_8588 = 5'h17 == com_idx ? rob_uop_23_edge_inst : _GEN_8587; // @[rob.scala 411:{25,25}]
  wire  _GEN_8589 = 5'h18 == com_idx ? rob_uop_24_edge_inst : _GEN_8588; // @[rob.scala 411:{25,25}]
  wire  _GEN_8590 = 5'h19 == com_idx ? rob_uop_25_edge_inst : _GEN_8589; // @[rob.scala 411:{25,25}]
  wire  _GEN_8591 = 5'h1a == com_idx ? rob_uop_26_edge_inst : _GEN_8590; // @[rob.scala 411:{25,25}]
  wire  _GEN_8592 = 5'h1b == com_idx ? rob_uop_27_edge_inst : _GEN_8591; // @[rob.scala 411:{25,25}]
  wire  _GEN_8593 = 5'h1c == com_idx ? rob_uop_28_edge_inst : _GEN_8592; // @[rob.scala 411:{25,25}]
  wire  _GEN_8594 = 5'h1d == com_idx ? rob_uop_29_edge_inst : _GEN_8593; // @[rob.scala 411:{25,25}]
  wire  _GEN_8595 = 5'h1e == com_idx ? rob_uop_30_edge_inst : _GEN_8594; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8598 = 5'h1 == com_idx ? rob_uop_1_ftq_idx : rob_uop_0_ftq_idx; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8599 = 5'h2 == com_idx ? rob_uop_2_ftq_idx : _GEN_8598; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8600 = 5'h3 == com_idx ? rob_uop_3_ftq_idx : _GEN_8599; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8601 = 5'h4 == com_idx ? rob_uop_4_ftq_idx : _GEN_8600; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8602 = 5'h5 == com_idx ? rob_uop_5_ftq_idx : _GEN_8601; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8603 = 5'h6 == com_idx ? rob_uop_6_ftq_idx : _GEN_8602; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8604 = 5'h7 == com_idx ? rob_uop_7_ftq_idx : _GEN_8603; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8605 = 5'h8 == com_idx ? rob_uop_8_ftq_idx : _GEN_8604; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8606 = 5'h9 == com_idx ? rob_uop_9_ftq_idx : _GEN_8605; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8607 = 5'ha == com_idx ? rob_uop_10_ftq_idx : _GEN_8606; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8608 = 5'hb == com_idx ? rob_uop_11_ftq_idx : _GEN_8607; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8609 = 5'hc == com_idx ? rob_uop_12_ftq_idx : _GEN_8608; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8610 = 5'hd == com_idx ? rob_uop_13_ftq_idx : _GEN_8609; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8611 = 5'he == com_idx ? rob_uop_14_ftq_idx : _GEN_8610; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8612 = 5'hf == com_idx ? rob_uop_15_ftq_idx : _GEN_8611; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8613 = 5'h10 == com_idx ? rob_uop_16_ftq_idx : _GEN_8612; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8614 = 5'h11 == com_idx ? rob_uop_17_ftq_idx : _GEN_8613; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8615 = 5'h12 == com_idx ? rob_uop_18_ftq_idx : _GEN_8614; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8616 = 5'h13 == com_idx ? rob_uop_19_ftq_idx : _GEN_8615; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8617 = 5'h14 == com_idx ? rob_uop_20_ftq_idx : _GEN_8616; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8618 = 5'h15 == com_idx ? rob_uop_21_ftq_idx : _GEN_8617; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8619 = 5'h16 == com_idx ? rob_uop_22_ftq_idx : _GEN_8618; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8620 = 5'h17 == com_idx ? rob_uop_23_ftq_idx : _GEN_8619; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8621 = 5'h18 == com_idx ? rob_uop_24_ftq_idx : _GEN_8620; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8622 = 5'h19 == com_idx ? rob_uop_25_ftq_idx : _GEN_8621; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8623 = 5'h1a == com_idx ? rob_uop_26_ftq_idx : _GEN_8622; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8624 = 5'h1b == com_idx ? rob_uop_27_ftq_idx : _GEN_8623; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8625 = 5'h1c == com_idx ? rob_uop_28_ftq_idx : _GEN_8624; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8626 = 5'h1d == com_idx ? rob_uop_29_ftq_idx : _GEN_8625; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_8627 = 5'h1e == com_idx ? rob_uop_30_ftq_idx : _GEN_8626; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8630 = 5'h1 == com_idx ? rob_uop_1_br_tag : rob_uop_0_br_tag; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8631 = 5'h2 == com_idx ? rob_uop_2_br_tag : _GEN_8630; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8632 = 5'h3 == com_idx ? rob_uop_3_br_tag : _GEN_8631; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8633 = 5'h4 == com_idx ? rob_uop_4_br_tag : _GEN_8632; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8634 = 5'h5 == com_idx ? rob_uop_5_br_tag : _GEN_8633; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8635 = 5'h6 == com_idx ? rob_uop_6_br_tag : _GEN_8634; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8636 = 5'h7 == com_idx ? rob_uop_7_br_tag : _GEN_8635; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8637 = 5'h8 == com_idx ? rob_uop_8_br_tag : _GEN_8636; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8638 = 5'h9 == com_idx ? rob_uop_9_br_tag : _GEN_8637; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8639 = 5'ha == com_idx ? rob_uop_10_br_tag : _GEN_8638; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8640 = 5'hb == com_idx ? rob_uop_11_br_tag : _GEN_8639; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8641 = 5'hc == com_idx ? rob_uop_12_br_tag : _GEN_8640; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8642 = 5'hd == com_idx ? rob_uop_13_br_tag : _GEN_8641; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8643 = 5'he == com_idx ? rob_uop_14_br_tag : _GEN_8642; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8644 = 5'hf == com_idx ? rob_uop_15_br_tag : _GEN_8643; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8645 = 5'h10 == com_idx ? rob_uop_16_br_tag : _GEN_8644; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8646 = 5'h11 == com_idx ? rob_uop_17_br_tag : _GEN_8645; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8647 = 5'h12 == com_idx ? rob_uop_18_br_tag : _GEN_8646; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8648 = 5'h13 == com_idx ? rob_uop_19_br_tag : _GEN_8647; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8649 = 5'h14 == com_idx ? rob_uop_20_br_tag : _GEN_8648; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8650 = 5'h15 == com_idx ? rob_uop_21_br_tag : _GEN_8649; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8651 = 5'h16 == com_idx ? rob_uop_22_br_tag : _GEN_8650; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8652 = 5'h17 == com_idx ? rob_uop_23_br_tag : _GEN_8651; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8653 = 5'h18 == com_idx ? rob_uop_24_br_tag : _GEN_8652; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8654 = 5'h19 == com_idx ? rob_uop_25_br_tag : _GEN_8653; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8655 = 5'h1a == com_idx ? rob_uop_26_br_tag : _GEN_8654; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8656 = 5'h1b == com_idx ? rob_uop_27_br_tag : _GEN_8655; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8657 = 5'h1c == com_idx ? rob_uop_28_br_tag : _GEN_8656; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8658 = 5'h1d == com_idx ? rob_uop_29_br_tag : _GEN_8657; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_8659 = 5'h1e == com_idx ? rob_uop_30_br_tag : _GEN_8658; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8662 = 5'h1 == com_idx ? rob_uop_1_br_mask : rob_uop_0_br_mask; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8663 = 5'h2 == com_idx ? rob_uop_2_br_mask : _GEN_8662; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8664 = 5'h3 == com_idx ? rob_uop_3_br_mask : _GEN_8663; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8665 = 5'h4 == com_idx ? rob_uop_4_br_mask : _GEN_8664; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8666 = 5'h5 == com_idx ? rob_uop_5_br_mask : _GEN_8665; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8667 = 5'h6 == com_idx ? rob_uop_6_br_mask : _GEN_8666; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8668 = 5'h7 == com_idx ? rob_uop_7_br_mask : _GEN_8667; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8669 = 5'h8 == com_idx ? rob_uop_8_br_mask : _GEN_8668; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8670 = 5'h9 == com_idx ? rob_uop_9_br_mask : _GEN_8669; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8671 = 5'ha == com_idx ? rob_uop_10_br_mask : _GEN_8670; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8672 = 5'hb == com_idx ? rob_uop_11_br_mask : _GEN_8671; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8673 = 5'hc == com_idx ? rob_uop_12_br_mask : _GEN_8672; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8674 = 5'hd == com_idx ? rob_uop_13_br_mask : _GEN_8673; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8675 = 5'he == com_idx ? rob_uop_14_br_mask : _GEN_8674; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8676 = 5'hf == com_idx ? rob_uop_15_br_mask : _GEN_8675; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8677 = 5'h10 == com_idx ? rob_uop_16_br_mask : _GEN_8676; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8678 = 5'h11 == com_idx ? rob_uop_17_br_mask : _GEN_8677; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8679 = 5'h12 == com_idx ? rob_uop_18_br_mask : _GEN_8678; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8680 = 5'h13 == com_idx ? rob_uop_19_br_mask : _GEN_8679; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8681 = 5'h14 == com_idx ? rob_uop_20_br_mask : _GEN_8680; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8682 = 5'h15 == com_idx ? rob_uop_21_br_mask : _GEN_8681; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8683 = 5'h16 == com_idx ? rob_uop_22_br_mask : _GEN_8682; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8684 = 5'h17 == com_idx ? rob_uop_23_br_mask : _GEN_8683; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8685 = 5'h18 == com_idx ? rob_uop_24_br_mask : _GEN_8684; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8686 = 5'h19 == com_idx ? rob_uop_25_br_mask : _GEN_8685; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8687 = 5'h1a == com_idx ? rob_uop_26_br_mask : _GEN_8686; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8688 = 5'h1b == com_idx ? rob_uop_27_br_mask : _GEN_8687; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8689 = 5'h1c == com_idx ? rob_uop_28_br_mask : _GEN_8688; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8690 = 5'h1d == com_idx ? rob_uop_29_br_mask : _GEN_8689; // @[rob.scala 411:{25,25}]
  wire [7:0] _GEN_8691 = 5'h1e == com_idx ? rob_uop_30_br_mask : _GEN_8690; // @[rob.scala 411:{25,25}]
  wire  _GEN_8694 = 5'h1 == com_idx ? rob_uop_1_is_sfb : rob_uop_0_is_sfb; // @[rob.scala 411:{25,25}]
  wire  _GEN_8695 = 5'h2 == com_idx ? rob_uop_2_is_sfb : _GEN_8694; // @[rob.scala 411:{25,25}]
  wire  _GEN_8696 = 5'h3 == com_idx ? rob_uop_3_is_sfb : _GEN_8695; // @[rob.scala 411:{25,25}]
  wire  _GEN_8697 = 5'h4 == com_idx ? rob_uop_4_is_sfb : _GEN_8696; // @[rob.scala 411:{25,25}]
  wire  _GEN_8698 = 5'h5 == com_idx ? rob_uop_5_is_sfb : _GEN_8697; // @[rob.scala 411:{25,25}]
  wire  _GEN_8699 = 5'h6 == com_idx ? rob_uop_6_is_sfb : _GEN_8698; // @[rob.scala 411:{25,25}]
  wire  _GEN_8700 = 5'h7 == com_idx ? rob_uop_7_is_sfb : _GEN_8699; // @[rob.scala 411:{25,25}]
  wire  _GEN_8701 = 5'h8 == com_idx ? rob_uop_8_is_sfb : _GEN_8700; // @[rob.scala 411:{25,25}]
  wire  _GEN_8702 = 5'h9 == com_idx ? rob_uop_9_is_sfb : _GEN_8701; // @[rob.scala 411:{25,25}]
  wire  _GEN_8703 = 5'ha == com_idx ? rob_uop_10_is_sfb : _GEN_8702; // @[rob.scala 411:{25,25}]
  wire  _GEN_8704 = 5'hb == com_idx ? rob_uop_11_is_sfb : _GEN_8703; // @[rob.scala 411:{25,25}]
  wire  _GEN_8705 = 5'hc == com_idx ? rob_uop_12_is_sfb : _GEN_8704; // @[rob.scala 411:{25,25}]
  wire  _GEN_8706 = 5'hd == com_idx ? rob_uop_13_is_sfb : _GEN_8705; // @[rob.scala 411:{25,25}]
  wire  _GEN_8707 = 5'he == com_idx ? rob_uop_14_is_sfb : _GEN_8706; // @[rob.scala 411:{25,25}]
  wire  _GEN_8708 = 5'hf == com_idx ? rob_uop_15_is_sfb : _GEN_8707; // @[rob.scala 411:{25,25}]
  wire  _GEN_8709 = 5'h10 == com_idx ? rob_uop_16_is_sfb : _GEN_8708; // @[rob.scala 411:{25,25}]
  wire  _GEN_8710 = 5'h11 == com_idx ? rob_uop_17_is_sfb : _GEN_8709; // @[rob.scala 411:{25,25}]
  wire  _GEN_8711 = 5'h12 == com_idx ? rob_uop_18_is_sfb : _GEN_8710; // @[rob.scala 411:{25,25}]
  wire  _GEN_8712 = 5'h13 == com_idx ? rob_uop_19_is_sfb : _GEN_8711; // @[rob.scala 411:{25,25}]
  wire  _GEN_8713 = 5'h14 == com_idx ? rob_uop_20_is_sfb : _GEN_8712; // @[rob.scala 411:{25,25}]
  wire  _GEN_8714 = 5'h15 == com_idx ? rob_uop_21_is_sfb : _GEN_8713; // @[rob.scala 411:{25,25}]
  wire  _GEN_8715 = 5'h16 == com_idx ? rob_uop_22_is_sfb : _GEN_8714; // @[rob.scala 411:{25,25}]
  wire  _GEN_8716 = 5'h17 == com_idx ? rob_uop_23_is_sfb : _GEN_8715; // @[rob.scala 411:{25,25}]
  wire  _GEN_8717 = 5'h18 == com_idx ? rob_uop_24_is_sfb : _GEN_8716; // @[rob.scala 411:{25,25}]
  wire  _GEN_8718 = 5'h19 == com_idx ? rob_uop_25_is_sfb : _GEN_8717; // @[rob.scala 411:{25,25}]
  wire  _GEN_8719 = 5'h1a == com_idx ? rob_uop_26_is_sfb : _GEN_8718; // @[rob.scala 411:{25,25}]
  wire  _GEN_8720 = 5'h1b == com_idx ? rob_uop_27_is_sfb : _GEN_8719; // @[rob.scala 411:{25,25}]
  wire  _GEN_8721 = 5'h1c == com_idx ? rob_uop_28_is_sfb : _GEN_8720; // @[rob.scala 411:{25,25}]
  wire  _GEN_8722 = 5'h1d == com_idx ? rob_uop_29_is_sfb : _GEN_8721; // @[rob.scala 411:{25,25}]
  wire  _GEN_8723 = 5'h1e == com_idx ? rob_uop_30_is_sfb : _GEN_8722; // @[rob.scala 411:{25,25}]
  wire  _GEN_8726 = 5'h1 == com_idx ? rob_uop_1_is_jal : rob_uop_0_is_jal; // @[rob.scala 411:{25,25}]
  wire  _GEN_8727 = 5'h2 == com_idx ? rob_uop_2_is_jal : _GEN_8726; // @[rob.scala 411:{25,25}]
  wire  _GEN_8728 = 5'h3 == com_idx ? rob_uop_3_is_jal : _GEN_8727; // @[rob.scala 411:{25,25}]
  wire  _GEN_8729 = 5'h4 == com_idx ? rob_uop_4_is_jal : _GEN_8728; // @[rob.scala 411:{25,25}]
  wire  _GEN_8730 = 5'h5 == com_idx ? rob_uop_5_is_jal : _GEN_8729; // @[rob.scala 411:{25,25}]
  wire  _GEN_8731 = 5'h6 == com_idx ? rob_uop_6_is_jal : _GEN_8730; // @[rob.scala 411:{25,25}]
  wire  _GEN_8732 = 5'h7 == com_idx ? rob_uop_7_is_jal : _GEN_8731; // @[rob.scala 411:{25,25}]
  wire  _GEN_8733 = 5'h8 == com_idx ? rob_uop_8_is_jal : _GEN_8732; // @[rob.scala 411:{25,25}]
  wire  _GEN_8734 = 5'h9 == com_idx ? rob_uop_9_is_jal : _GEN_8733; // @[rob.scala 411:{25,25}]
  wire  _GEN_8735 = 5'ha == com_idx ? rob_uop_10_is_jal : _GEN_8734; // @[rob.scala 411:{25,25}]
  wire  _GEN_8736 = 5'hb == com_idx ? rob_uop_11_is_jal : _GEN_8735; // @[rob.scala 411:{25,25}]
  wire  _GEN_8737 = 5'hc == com_idx ? rob_uop_12_is_jal : _GEN_8736; // @[rob.scala 411:{25,25}]
  wire  _GEN_8738 = 5'hd == com_idx ? rob_uop_13_is_jal : _GEN_8737; // @[rob.scala 411:{25,25}]
  wire  _GEN_8739 = 5'he == com_idx ? rob_uop_14_is_jal : _GEN_8738; // @[rob.scala 411:{25,25}]
  wire  _GEN_8740 = 5'hf == com_idx ? rob_uop_15_is_jal : _GEN_8739; // @[rob.scala 411:{25,25}]
  wire  _GEN_8741 = 5'h10 == com_idx ? rob_uop_16_is_jal : _GEN_8740; // @[rob.scala 411:{25,25}]
  wire  _GEN_8742 = 5'h11 == com_idx ? rob_uop_17_is_jal : _GEN_8741; // @[rob.scala 411:{25,25}]
  wire  _GEN_8743 = 5'h12 == com_idx ? rob_uop_18_is_jal : _GEN_8742; // @[rob.scala 411:{25,25}]
  wire  _GEN_8744 = 5'h13 == com_idx ? rob_uop_19_is_jal : _GEN_8743; // @[rob.scala 411:{25,25}]
  wire  _GEN_8745 = 5'h14 == com_idx ? rob_uop_20_is_jal : _GEN_8744; // @[rob.scala 411:{25,25}]
  wire  _GEN_8746 = 5'h15 == com_idx ? rob_uop_21_is_jal : _GEN_8745; // @[rob.scala 411:{25,25}]
  wire  _GEN_8747 = 5'h16 == com_idx ? rob_uop_22_is_jal : _GEN_8746; // @[rob.scala 411:{25,25}]
  wire  _GEN_8748 = 5'h17 == com_idx ? rob_uop_23_is_jal : _GEN_8747; // @[rob.scala 411:{25,25}]
  wire  _GEN_8749 = 5'h18 == com_idx ? rob_uop_24_is_jal : _GEN_8748; // @[rob.scala 411:{25,25}]
  wire  _GEN_8750 = 5'h19 == com_idx ? rob_uop_25_is_jal : _GEN_8749; // @[rob.scala 411:{25,25}]
  wire  _GEN_8751 = 5'h1a == com_idx ? rob_uop_26_is_jal : _GEN_8750; // @[rob.scala 411:{25,25}]
  wire  _GEN_8752 = 5'h1b == com_idx ? rob_uop_27_is_jal : _GEN_8751; // @[rob.scala 411:{25,25}]
  wire  _GEN_8753 = 5'h1c == com_idx ? rob_uop_28_is_jal : _GEN_8752; // @[rob.scala 411:{25,25}]
  wire  _GEN_8754 = 5'h1d == com_idx ? rob_uop_29_is_jal : _GEN_8753; // @[rob.scala 411:{25,25}]
  wire  _GEN_8755 = 5'h1e == com_idx ? rob_uop_30_is_jal : _GEN_8754; // @[rob.scala 411:{25,25}]
  wire  _GEN_8758 = 5'h1 == com_idx ? rob_uop_1_is_jalr : rob_uop_0_is_jalr; // @[rob.scala 411:{25,25}]
  wire  _GEN_8759 = 5'h2 == com_idx ? rob_uop_2_is_jalr : _GEN_8758; // @[rob.scala 411:{25,25}]
  wire  _GEN_8760 = 5'h3 == com_idx ? rob_uop_3_is_jalr : _GEN_8759; // @[rob.scala 411:{25,25}]
  wire  _GEN_8761 = 5'h4 == com_idx ? rob_uop_4_is_jalr : _GEN_8760; // @[rob.scala 411:{25,25}]
  wire  _GEN_8762 = 5'h5 == com_idx ? rob_uop_5_is_jalr : _GEN_8761; // @[rob.scala 411:{25,25}]
  wire  _GEN_8763 = 5'h6 == com_idx ? rob_uop_6_is_jalr : _GEN_8762; // @[rob.scala 411:{25,25}]
  wire  _GEN_8764 = 5'h7 == com_idx ? rob_uop_7_is_jalr : _GEN_8763; // @[rob.scala 411:{25,25}]
  wire  _GEN_8765 = 5'h8 == com_idx ? rob_uop_8_is_jalr : _GEN_8764; // @[rob.scala 411:{25,25}]
  wire  _GEN_8766 = 5'h9 == com_idx ? rob_uop_9_is_jalr : _GEN_8765; // @[rob.scala 411:{25,25}]
  wire  _GEN_8767 = 5'ha == com_idx ? rob_uop_10_is_jalr : _GEN_8766; // @[rob.scala 411:{25,25}]
  wire  _GEN_8768 = 5'hb == com_idx ? rob_uop_11_is_jalr : _GEN_8767; // @[rob.scala 411:{25,25}]
  wire  _GEN_8769 = 5'hc == com_idx ? rob_uop_12_is_jalr : _GEN_8768; // @[rob.scala 411:{25,25}]
  wire  _GEN_8770 = 5'hd == com_idx ? rob_uop_13_is_jalr : _GEN_8769; // @[rob.scala 411:{25,25}]
  wire  _GEN_8771 = 5'he == com_idx ? rob_uop_14_is_jalr : _GEN_8770; // @[rob.scala 411:{25,25}]
  wire  _GEN_8772 = 5'hf == com_idx ? rob_uop_15_is_jalr : _GEN_8771; // @[rob.scala 411:{25,25}]
  wire  _GEN_8773 = 5'h10 == com_idx ? rob_uop_16_is_jalr : _GEN_8772; // @[rob.scala 411:{25,25}]
  wire  _GEN_8774 = 5'h11 == com_idx ? rob_uop_17_is_jalr : _GEN_8773; // @[rob.scala 411:{25,25}]
  wire  _GEN_8775 = 5'h12 == com_idx ? rob_uop_18_is_jalr : _GEN_8774; // @[rob.scala 411:{25,25}]
  wire  _GEN_8776 = 5'h13 == com_idx ? rob_uop_19_is_jalr : _GEN_8775; // @[rob.scala 411:{25,25}]
  wire  _GEN_8777 = 5'h14 == com_idx ? rob_uop_20_is_jalr : _GEN_8776; // @[rob.scala 411:{25,25}]
  wire  _GEN_8778 = 5'h15 == com_idx ? rob_uop_21_is_jalr : _GEN_8777; // @[rob.scala 411:{25,25}]
  wire  _GEN_8779 = 5'h16 == com_idx ? rob_uop_22_is_jalr : _GEN_8778; // @[rob.scala 411:{25,25}]
  wire  _GEN_8780 = 5'h17 == com_idx ? rob_uop_23_is_jalr : _GEN_8779; // @[rob.scala 411:{25,25}]
  wire  _GEN_8781 = 5'h18 == com_idx ? rob_uop_24_is_jalr : _GEN_8780; // @[rob.scala 411:{25,25}]
  wire  _GEN_8782 = 5'h19 == com_idx ? rob_uop_25_is_jalr : _GEN_8781; // @[rob.scala 411:{25,25}]
  wire  _GEN_8783 = 5'h1a == com_idx ? rob_uop_26_is_jalr : _GEN_8782; // @[rob.scala 411:{25,25}]
  wire  _GEN_8784 = 5'h1b == com_idx ? rob_uop_27_is_jalr : _GEN_8783; // @[rob.scala 411:{25,25}]
  wire  _GEN_8785 = 5'h1c == com_idx ? rob_uop_28_is_jalr : _GEN_8784; // @[rob.scala 411:{25,25}]
  wire  _GEN_8786 = 5'h1d == com_idx ? rob_uop_29_is_jalr : _GEN_8785; // @[rob.scala 411:{25,25}]
  wire  _GEN_8787 = 5'h1e == com_idx ? rob_uop_30_is_jalr : _GEN_8786; // @[rob.scala 411:{25,25}]
  wire  _GEN_8790 = 5'h1 == com_idx ? rob_uop_1_is_br : rob_uop_0_is_br; // @[rob.scala 411:{25,25}]
  wire  _GEN_8791 = 5'h2 == com_idx ? rob_uop_2_is_br : _GEN_8790; // @[rob.scala 411:{25,25}]
  wire  _GEN_8792 = 5'h3 == com_idx ? rob_uop_3_is_br : _GEN_8791; // @[rob.scala 411:{25,25}]
  wire  _GEN_8793 = 5'h4 == com_idx ? rob_uop_4_is_br : _GEN_8792; // @[rob.scala 411:{25,25}]
  wire  _GEN_8794 = 5'h5 == com_idx ? rob_uop_5_is_br : _GEN_8793; // @[rob.scala 411:{25,25}]
  wire  _GEN_8795 = 5'h6 == com_idx ? rob_uop_6_is_br : _GEN_8794; // @[rob.scala 411:{25,25}]
  wire  _GEN_8796 = 5'h7 == com_idx ? rob_uop_7_is_br : _GEN_8795; // @[rob.scala 411:{25,25}]
  wire  _GEN_8797 = 5'h8 == com_idx ? rob_uop_8_is_br : _GEN_8796; // @[rob.scala 411:{25,25}]
  wire  _GEN_8798 = 5'h9 == com_idx ? rob_uop_9_is_br : _GEN_8797; // @[rob.scala 411:{25,25}]
  wire  _GEN_8799 = 5'ha == com_idx ? rob_uop_10_is_br : _GEN_8798; // @[rob.scala 411:{25,25}]
  wire  _GEN_8800 = 5'hb == com_idx ? rob_uop_11_is_br : _GEN_8799; // @[rob.scala 411:{25,25}]
  wire  _GEN_8801 = 5'hc == com_idx ? rob_uop_12_is_br : _GEN_8800; // @[rob.scala 411:{25,25}]
  wire  _GEN_8802 = 5'hd == com_idx ? rob_uop_13_is_br : _GEN_8801; // @[rob.scala 411:{25,25}]
  wire  _GEN_8803 = 5'he == com_idx ? rob_uop_14_is_br : _GEN_8802; // @[rob.scala 411:{25,25}]
  wire  _GEN_8804 = 5'hf == com_idx ? rob_uop_15_is_br : _GEN_8803; // @[rob.scala 411:{25,25}]
  wire  _GEN_8805 = 5'h10 == com_idx ? rob_uop_16_is_br : _GEN_8804; // @[rob.scala 411:{25,25}]
  wire  _GEN_8806 = 5'h11 == com_idx ? rob_uop_17_is_br : _GEN_8805; // @[rob.scala 411:{25,25}]
  wire  _GEN_8807 = 5'h12 == com_idx ? rob_uop_18_is_br : _GEN_8806; // @[rob.scala 411:{25,25}]
  wire  _GEN_8808 = 5'h13 == com_idx ? rob_uop_19_is_br : _GEN_8807; // @[rob.scala 411:{25,25}]
  wire  _GEN_8809 = 5'h14 == com_idx ? rob_uop_20_is_br : _GEN_8808; // @[rob.scala 411:{25,25}]
  wire  _GEN_8810 = 5'h15 == com_idx ? rob_uop_21_is_br : _GEN_8809; // @[rob.scala 411:{25,25}]
  wire  _GEN_8811 = 5'h16 == com_idx ? rob_uop_22_is_br : _GEN_8810; // @[rob.scala 411:{25,25}]
  wire  _GEN_8812 = 5'h17 == com_idx ? rob_uop_23_is_br : _GEN_8811; // @[rob.scala 411:{25,25}]
  wire  _GEN_8813 = 5'h18 == com_idx ? rob_uop_24_is_br : _GEN_8812; // @[rob.scala 411:{25,25}]
  wire  _GEN_8814 = 5'h19 == com_idx ? rob_uop_25_is_br : _GEN_8813; // @[rob.scala 411:{25,25}]
  wire  _GEN_8815 = 5'h1a == com_idx ? rob_uop_26_is_br : _GEN_8814; // @[rob.scala 411:{25,25}]
  wire  _GEN_8816 = 5'h1b == com_idx ? rob_uop_27_is_br : _GEN_8815; // @[rob.scala 411:{25,25}]
  wire  _GEN_8817 = 5'h1c == com_idx ? rob_uop_28_is_br : _GEN_8816; // @[rob.scala 411:{25,25}]
  wire  _GEN_8818 = 5'h1d == com_idx ? rob_uop_29_is_br : _GEN_8817; // @[rob.scala 411:{25,25}]
  wire  _GEN_8819 = 5'h1e == com_idx ? rob_uop_30_is_br : _GEN_8818; // @[rob.scala 411:{25,25}]
  wire  _GEN_8822 = 5'h1 == com_idx ? rob_uop_1_iw_p2_poisoned : rob_uop_0_iw_p2_poisoned; // @[rob.scala 411:{25,25}]
  wire  _GEN_8823 = 5'h2 == com_idx ? rob_uop_2_iw_p2_poisoned : _GEN_8822; // @[rob.scala 411:{25,25}]
  wire  _GEN_8824 = 5'h3 == com_idx ? rob_uop_3_iw_p2_poisoned : _GEN_8823; // @[rob.scala 411:{25,25}]
  wire  _GEN_8825 = 5'h4 == com_idx ? rob_uop_4_iw_p2_poisoned : _GEN_8824; // @[rob.scala 411:{25,25}]
  wire  _GEN_8826 = 5'h5 == com_idx ? rob_uop_5_iw_p2_poisoned : _GEN_8825; // @[rob.scala 411:{25,25}]
  wire  _GEN_8827 = 5'h6 == com_idx ? rob_uop_6_iw_p2_poisoned : _GEN_8826; // @[rob.scala 411:{25,25}]
  wire  _GEN_8828 = 5'h7 == com_idx ? rob_uop_7_iw_p2_poisoned : _GEN_8827; // @[rob.scala 411:{25,25}]
  wire  _GEN_8829 = 5'h8 == com_idx ? rob_uop_8_iw_p2_poisoned : _GEN_8828; // @[rob.scala 411:{25,25}]
  wire  _GEN_8830 = 5'h9 == com_idx ? rob_uop_9_iw_p2_poisoned : _GEN_8829; // @[rob.scala 411:{25,25}]
  wire  _GEN_8831 = 5'ha == com_idx ? rob_uop_10_iw_p2_poisoned : _GEN_8830; // @[rob.scala 411:{25,25}]
  wire  _GEN_8832 = 5'hb == com_idx ? rob_uop_11_iw_p2_poisoned : _GEN_8831; // @[rob.scala 411:{25,25}]
  wire  _GEN_8833 = 5'hc == com_idx ? rob_uop_12_iw_p2_poisoned : _GEN_8832; // @[rob.scala 411:{25,25}]
  wire  _GEN_8834 = 5'hd == com_idx ? rob_uop_13_iw_p2_poisoned : _GEN_8833; // @[rob.scala 411:{25,25}]
  wire  _GEN_8835 = 5'he == com_idx ? rob_uop_14_iw_p2_poisoned : _GEN_8834; // @[rob.scala 411:{25,25}]
  wire  _GEN_8836 = 5'hf == com_idx ? rob_uop_15_iw_p2_poisoned : _GEN_8835; // @[rob.scala 411:{25,25}]
  wire  _GEN_8837 = 5'h10 == com_idx ? rob_uop_16_iw_p2_poisoned : _GEN_8836; // @[rob.scala 411:{25,25}]
  wire  _GEN_8838 = 5'h11 == com_idx ? rob_uop_17_iw_p2_poisoned : _GEN_8837; // @[rob.scala 411:{25,25}]
  wire  _GEN_8839 = 5'h12 == com_idx ? rob_uop_18_iw_p2_poisoned : _GEN_8838; // @[rob.scala 411:{25,25}]
  wire  _GEN_8840 = 5'h13 == com_idx ? rob_uop_19_iw_p2_poisoned : _GEN_8839; // @[rob.scala 411:{25,25}]
  wire  _GEN_8841 = 5'h14 == com_idx ? rob_uop_20_iw_p2_poisoned : _GEN_8840; // @[rob.scala 411:{25,25}]
  wire  _GEN_8842 = 5'h15 == com_idx ? rob_uop_21_iw_p2_poisoned : _GEN_8841; // @[rob.scala 411:{25,25}]
  wire  _GEN_8843 = 5'h16 == com_idx ? rob_uop_22_iw_p2_poisoned : _GEN_8842; // @[rob.scala 411:{25,25}]
  wire  _GEN_8844 = 5'h17 == com_idx ? rob_uop_23_iw_p2_poisoned : _GEN_8843; // @[rob.scala 411:{25,25}]
  wire  _GEN_8845 = 5'h18 == com_idx ? rob_uop_24_iw_p2_poisoned : _GEN_8844; // @[rob.scala 411:{25,25}]
  wire  _GEN_8846 = 5'h19 == com_idx ? rob_uop_25_iw_p2_poisoned : _GEN_8845; // @[rob.scala 411:{25,25}]
  wire  _GEN_8847 = 5'h1a == com_idx ? rob_uop_26_iw_p2_poisoned : _GEN_8846; // @[rob.scala 411:{25,25}]
  wire  _GEN_8848 = 5'h1b == com_idx ? rob_uop_27_iw_p2_poisoned : _GEN_8847; // @[rob.scala 411:{25,25}]
  wire  _GEN_8849 = 5'h1c == com_idx ? rob_uop_28_iw_p2_poisoned : _GEN_8848; // @[rob.scala 411:{25,25}]
  wire  _GEN_8850 = 5'h1d == com_idx ? rob_uop_29_iw_p2_poisoned : _GEN_8849; // @[rob.scala 411:{25,25}]
  wire  _GEN_8851 = 5'h1e == com_idx ? rob_uop_30_iw_p2_poisoned : _GEN_8850; // @[rob.scala 411:{25,25}]
  wire  _GEN_8854 = 5'h1 == com_idx ? rob_uop_1_iw_p1_poisoned : rob_uop_0_iw_p1_poisoned; // @[rob.scala 411:{25,25}]
  wire  _GEN_8855 = 5'h2 == com_idx ? rob_uop_2_iw_p1_poisoned : _GEN_8854; // @[rob.scala 411:{25,25}]
  wire  _GEN_8856 = 5'h3 == com_idx ? rob_uop_3_iw_p1_poisoned : _GEN_8855; // @[rob.scala 411:{25,25}]
  wire  _GEN_8857 = 5'h4 == com_idx ? rob_uop_4_iw_p1_poisoned : _GEN_8856; // @[rob.scala 411:{25,25}]
  wire  _GEN_8858 = 5'h5 == com_idx ? rob_uop_5_iw_p1_poisoned : _GEN_8857; // @[rob.scala 411:{25,25}]
  wire  _GEN_8859 = 5'h6 == com_idx ? rob_uop_6_iw_p1_poisoned : _GEN_8858; // @[rob.scala 411:{25,25}]
  wire  _GEN_8860 = 5'h7 == com_idx ? rob_uop_7_iw_p1_poisoned : _GEN_8859; // @[rob.scala 411:{25,25}]
  wire  _GEN_8861 = 5'h8 == com_idx ? rob_uop_8_iw_p1_poisoned : _GEN_8860; // @[rob.scala 411:{25,25}]
  wire  _GEN_8862 = 5'h9 == com_idx ? rob_uop_9_iw_p1_poisoned : _GEN_8861; // @[rob.scala 411:{25,25}]
  wire  _GEN_8863 = 5'ha == com_idx ? rob_uop_10_iw_p1_poisoned : _GEN_8862; // @[rob.scala 411:{25,25}]
  wire  _GEN_8864 = 5'hb == com_idx ? rob_uop_11_iw_p1_poisoned : _GEN_8863; // @[rob.scala 411:{25,25}]
  wire  _GEN_8865 = 5'hc == com_idx ? rob_uop_12_iw_p1_poisoned : _GEN_8864; // @[rob.scala 411:{25,25}]
  wire  _GEN_8866 = 5'hd == com_idx ? rob_uop_13_iw_p1_poisoned : _GEN_8865; // @[rob.scala 411:{25,25}]
  wire  _GEN_8867 = 5'he == com_idx ? rob_uop_14_iw_p1_poisoned : _GEN_8866; // @[rob.scala 411:{25,25}]
  wire  _GEN_8868 = 5'hf == com_idx ? rob_uop_15_iw_p1_poisoned : _GEN_8867; // @[rob.scala 411:{25,25}]
  wire  _GEN_8869 = 5'h10 == com_idx ? rob_uop_16_iw_p1_poisoned : _GEN_8868; // @[rob.scala 411:{25,25}]
  wire  _GEN_8870 = 5'h11 == com_idx ? rob_uop_17_iw_p1_poisoned : _GEN_8869; // @[rob.scala 411:{25,25}]
  wire  _GEN_8871 = 5'h12 == com_idx ? rob_uop_18_iw_p1_poisoned : _GEN_8870; // @[rob.scala 411:{25,25}]
  wire  _GEN_8872 = 5'h13 == com_idx ? rob_uop_19_iw_p1_poisoned : _GEN_8871; // @[rob.scala 411:{25,25}]
  wire  _GEN_8873 = 5'h14 == com_idx ? rob_uop_20_iw_p1_poisoned : _GEN_8872; // @[rob.scala 411:{25,25}]
  wire  _GEN_8874 = 5'h15 == com_idx ? rob_uop_21_iw_p1_poisoned : _GEN_8873; // @[rob.scala 411:{25,25}]
  wire  _GEN_8875 = 5'h16 == com_idx ? rob_uop_22_iw_p1_poisoned : _GEN_8874; // @[rob.scala 411:{25,25}]
  wire  _GEN_8876 = 5'h17 == com_idx ? rob_uop_23_iw_p1_poisoned : _GEN_8875; // @[rob.scala 411:{25,25}]
  wire  _GEN_8877 = 5'h18 == com_idx ? rob_uop_24_iw_p1_poisoned : _GEN_8876; // @[rob.scala 411:{25,25}]
  wire  _GEN_8878 = 5'h19 == com_idx ? rob_uop_25_iw_p1_poisoned : _GEN_8877; // @[rob.scala 411:{25,25}]
  wire  _GEN_8879 = 5'h1a == com_idx ? rob_uop_26_iw_p1_poisoned : _GEN_8878; // @[rob.scala 411:{25,25}]
  wire  _GEN_8880 = 5'h1b == com_idx ? rob_uop_27_iw_p1_poisoned : _GEN_8879; // @[rob.scala 411:{25,25}]
  wire  _GEN_8881 = 5'h1c == com_idx ? rob_uop_28_iw_p1_poisoned : _GEN_8880; // @[rob.scala 411:{25,25}]
  wire  _GEN_8882 = 5'h1d == com_idx ? rob_uop_29_iw_p1_poisoned : _GEN_8881; // @[rob.scala 411:{25,25}]
  wire  _GEN_8883 = 5'h1e == com_idx ? rob_uop_30_iw_p1_poisoned : _GEN_8882; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8886 = 5'h1 == com_idx ? rob_uop_1_iw_state : rob_uop_0_iw_state; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8887 = 5'h2 == com_idx ? rob_uop_2_iw_state : _GEN_8886; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8888 = 5'h3 == com_idx ? rob_uop_3_iw_state : _GEN_8887; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8889 = 5'h4 == com_idx ? rob_uop_4_iw_state : _GEN_8888; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8890 = 5'h5 == com_idx ? rob_uop_5_iw_state : _GEN_8889; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8891 = 5'h6 == com_idx ? rob_uop_6_iw_state : _GEN_8890; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8892 = 5'h7 == com_idx ? rob_uop_7_iw_state : _GEN_8891; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8893 = 5'h8 == com_idx ? rob_uop_8_iw_state : _GEN_8892; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8894 = 5'h9 == com_idx ? rob_uop_9_iw_state : _GEN_8893; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8895 = 5'ha == com_idx ? rob_uop_10_iw_state : _GEN_8894; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8896 = 5'hb == com_idx ? rob_uop_11_iw_state : _GEN_8895; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8897 = 5'hc == com_idx ? rob_uop_12_iw_state : _GEN_8896; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8898 = 5'hd == com_idx ? rob_uop_13_iw_state : _GEN_8897; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8899 = 5'he == com_idx ? rob_uop_14_iw_state : _GEN_8898; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8900 = 5'hf == com_idx ? rob_uop_15_iw_state : _GEN_8899; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8901 = 5'h10 == com_idx ? rob_uop_16_iw_state : _GEN_8900; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8902 = 5'h11 == com_idx ? rob_uop_17_iw_state : _GEN_8901; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8903 = 5'h12 == com_idx ? rob_uop_18_iw_state : _GEN_8902; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8904 = 5'h13 == com_idx ? rob_uop_19_iw_state : _GEN_8903; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8905 = 5'h14 == com_idx ? rob_uop_20_iw_state : _GEN_8904; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8906 = 5'h15 == com_idx ? rob_uop_21_iw_state : _GEN_8905; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8907 = 5'h16 == com_idx ? rob_uop_22_iw_state : _GEN_8906; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8908 = 5'h17 == com_idx ? rob_uop_23_iw_state : _GEN_8907; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8909 = 5'h18 == com_idx ? rob_uop_24_iw_state : _GEN_8908; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8910 = 5'h19 == com_idx ? rob_uop_25_iw_state : _GEN_8909; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8911 = 5'h1a == com_idx ? rob_uop_26_iw_state : _GEN_8910; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8912 = 5'h1b == com_idx ? rob_uop_27_iw_state : _GEN_8911; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8913 = 5'h1c == com_idx ? rob_uop_28_iw_state : _GEN_8912; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8914 = 5'h1d == com_idx ? rob_uop_29_iw_state : _GEN_8913; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_8915 = 5'h1e == com_idx ? rob_uop_30_iw_state : _GEN_8914; // @[rob.scala 411:{25,25}]
  wire  _GEN_8918 = 5'h1 == com_idx ? rob_uop_1_ctrl_is_std : rob_uop_0_ctrl_is_std; // @[rob.scala 411:{25,25}]
  wire  _GEN_8919 = 5'h2 == com_idx ? rob_uop_2_ctrl_is_std : _GEN_8918; // @[rob.scala 411:{25,25}]
  wire  _GEN_8920 = 5'h3 == com_idx ? rob_uop_3_ctrl_is_std : _GEN_8919; // @[rob.scala 411:{25,25}]
  wire  _GEN_8921 = 5'h4 == com_idx ? rob_uop_4_ctrl_is_std : _GEN_8920; // @[rob.scala 411:{25,25}]
  wire  _GEN_8922 = 5'h5 == com_idx ? rob_uop_5_ctrl_is_std : _GEN_8921; // @[rob.scala 411:{25,25}]
  wire  _GEN_8923 = 5'h6 == com_idx ? rob_uop_6_ctrl_is_std : _GEN_8922; // @[rob.scala 411:{25,25}]
  wire  _GEN_8924 = 5'h7 == com_idx ? rob_uop_7_ctrl_is_std : _GEN_8923; // @[rob.scala 411:{25,25}]
  wire  _GEN_8925 = 5'h8 == com_idx ? rob_uop_8_ctrl_is_std : _GEN_8924; // @[rob.scala 411:{25,25}]
  wire  _GEN_8926 = 5'h9 == com_idx ? rob_uop_9_ctrl_is_std : _GEN_8925; // @[rob.scala 411:{25,25}]
  wire  _GEN_8927 = 5'ha == com_idx ? rob_uop_10_ctrl_is_std : _GEN_8926; // @[rob.scala 411:{25,25}]
  wire  _GEN_8928 = 5'hb == com_idx ? rob_uop_11_ctrl_is_std : _GEN_8927; // @[rob.scala 411:{25,25}]
  wire  _GEN_8929 = 5'hc == com_idx ? rob_uop_12_ctrl_is_std : _GEN_8928; // @[rob.scala 411:{25,25}]
  wire  _GEN_8930 = 5'hd == com_idx ? rob_uop_13_ctrl_is_std : _GEN_8929; // @[rob.scala 411:{25,25}]
  wire  _GEN_8931 = 5'he == com_idx ? rob_uop_14_ctrl_is_std : _GEN_8930; // @[rob.scala 411:{25,25}]
  wire  _GEN_8932 = 5'hf == com_idx ? rob_uop_15_ctrl_is_std : _GEN_8931; // @[rob.scala 411:{25,25}]
  wire  _GEN_8933 = 5'h10 == com_idx ? rob_uop_16_ctrl_is_std : _GEN_8932; // @[rob.scala 411:{25,25}]
  wire  _GEN_8934 = 5'h11 == com_idx ? rob_uop_17_ctrl_is_std : _GEN_8933; // @[rob.scala 411:{25,25}]
  wire  _GEN_8935 = 5'h12 == com_idx ? rob_uop_18_ctrl_is_std : _GEN_8934; // @[rob.scala 411:{25,25}]
  wire  _GEN_8936 = 5'h13 == com_idx ? rob_uop_19_ctrl_is_std : _GEN_8935; // @[rob.scala 411:{25,25}]
  wire  _GEN_8937 = 5'h14 == com_idx ? rob_uop_20_ctrl_is_std : _GEN_8936; // @[rob.scala 411:{25,25}]
  wire  _GEN_8938 = 5'h15 == com_idx ? rob_uop_21_ctrl_is_std : _GEN_8937; // @[rob.scala 411:{25,25}]
  wire  _GEN_8939 = 5'h16 == com_idx ? rob_uop_22_ctrl_is_std : _GEN_8938; // @[rob.scala 411:{25,25}]
  wire  _GEN_8940 = 5'h17 == com_idx ? rob_uop_23_ctrl_is_std : _GEN_8939; // @[rob.scala 411:{25,25}]
  wire  _GEN_8941 = 5'h18 == com_idx ? rob_uop_24_ctrl_is_std : _GEN_8940; // @[rob.scala 411:{25,25}]
  wire  _GEN_8942 = 5'h19 == com_idx ? rob_uop_25_ctrl_is_std : _GEN_8941; // @[rob.scala 411:{25,25}]
  wire  _GEN_8943 = 5'h1a == com_idx ? rob_uop_26_ctrl_is_std : _GEN_8942; // @[rob.scala 411:{25,25}]
  wire  _GEN_8944 = 5'h1b == com_idx ? rob_uop_27_ctrl_is_std : _GEN_8943; // @[rob.scala 411:{25,25}]
  wire  _GEN_8945 = 5'h1c == com_idx ? rob_uop_28_ctrl_is_std : _GEN_8944; // @[rob.scala 411:{25,25}]
  wire  _GEN_8946 = 5'h1d == com_idx ? rob_uop_29_ctrl_is_std : _GEN_8945; // @[rob.scala 411:{25,25}]
  wire  _GEN_8947 = 5'h1e == com_idx ? rob_uop_30_ctrl_is_std : _GEN_8946; // @[rob.scala 411:{25,25}]
  wire  _GEN_8950 = 5'h1 == com_idx ? rob_uop_1_ctrl_is_sta : rob_uop_0_ctrl_is_sta; // @[rob.scala 411:{25,25}]
  wire  _GEN_8951 = 5'h2 == com_idx ? rob_uop_2_ctrl_is_sta : _GEN_8950; // @[rob.scala 411:{25,25}]
  wire  _GEN_8952 = 5'h3 == com_idx ? rob_uop_3_ctrl_is_sta : _GEN_8951; // @[rob.scala 411:{25,25}]
  wire  _GEN_8953 = 5'h4 == com_idx ? rob_uop_4_ctrl_is_sta : _GEN_8952; // @[rob.scala 411:{25,25}]
  wire  _GEN_8954 = 5'h5 == com_idx ? rob_uop_5_ctrl_is_sta : _GEN_8953; // @[rob.scala 411:{25,25}]
  wire  _GEN_8955 = 5'h6 == com_idx ? rob_uop_6_ctrl_is_sta : _GEN_8954; // @[rob.scala 411:{25,25}]
  wire  _GEN_8956 = 5'h7 == com_idx ? rob_uop_7_ctrl_is_sta : _GEN_8955; // @[rob.scala 411:{25,25}]
  wire  _GEN_8957 = 5'h8 == com_idx ? rob_uop_8_ctrl_is_sta : _GEN_8956; // @[rob.scala 411:{25,25}]
  wire  _GEN_8958 = 5'h9 == com_idx ? rob_uop_9_ctrl_is_sta : _GEN_8957; // @[rob.scala 411:{25,25}]
  wire  _GEN_8959 = 5'ha == com_idx ? rob_uop_10_ctrl_is_sta : _GEN_8958; // @[rob.scala 411:{25,25}]
  wire  _GEN_8960 = 5'hb == com_idx ? rob_uop_11_ctrl_is_sta : _GEN_8959; // @[rob.scala 411:{25,25}]
  wire  _GEN_8961 = 5'hc == com_idx ? rob_uop_12_ctrl_is_sta : _GEN_8960; // @[rob.scala 411:{25,25}]
  wire  _GEN_8962 = 5'hd == com_idx ? rob_uop_13_ctrl_is_sta : _GEN_8961; // @[rob.scala 411:{25,25}]
  wire  _GEN_8963 = 5'he == com_idx ? rob_uop_14_ctrl_is_sta : _GEN_8962; // @[rob.scala 411:{25,25}]
  wire  _GEN_8964 = 5'hf == com_idx ? rob_uop_15_ctrl_is_sta : _GEN_8963; // @[rob.scala 411:{25,25}]
  wire  _GEN_8965 = 5'h10 == com_idx ? rob_uop_16_ctrl_is_sta : _GEN_8964; // @[rob.scala 411:{25,25}]
  wire  _GEN_8966 = 5'h11 == com_idx ? rob_uop_17_ctrl_is_sta : _GEN_8965; // @[rob.scala 411:{25,25}]
  wire  _GEN_8967 = 5'h12 == com_idx ? rob_uop_18_ctrl_is_sta : _GEN_8966; // @[rob.scala 411:{25,25}]
  wire  _GEN_8968 = 5'h13 == com_idx ? rob_uop_19_ctrl_is_sta : _GEN_8967; // @[rob.scala 411:{25,25}]
  wire  _GEN_8969 = 5'h14 == com_idx ? rob_uop_20_ctrl_is_sta : _GEN_8968; // @[rob.scala 411:{25,25}]
  wire  _GEN_8970 = 5'h15 == com_idx ? rob_uop_21_ctrl_is_sta : _GEN_8969; // @[rob.scala 411:{25,25}]
  wire  _GEN_8971 = 5'h16 == com_idx ? rob_uop_22_ctrl_is_sta : _GEN_8970; // @[rob.scala 411:{25,25}]
  wire  _GEN_8972 = 5'h17 == com_idx ? rob_uop_23_ctrl_is_sta : _GEN_8971; // @[rob.scala 411:{25,25}]
  wire  _GEN_8973 = 5'h18 == com_idx ? rob_uop_24_ctrl_is_sta : _GEN_8972; // @[rob.scala 411:{25,25}]
  wire  _GEN_8974 = 5'h19 == com_idx ? rob_uop_25_ctrl_is_sta : _GEN_8973; // @[rob.scala 411:{25,25}]
  wire  _GEN_8975 = 5'h1a == com_idx ? rob_uop_26_ctrl_is_sta : _GEN_8974; // @[rob.scala 411:{25,25}]
  wire  _GEN_8976 = 5'h1b == com_idx ? rob_uop_27_ctrl_is_sta : _GEN_8975; // @[rob.scala 411:{25,25}]
  wire  _GEN_8977 = 5'h1c == com_idx ? rob_uop_28_ctrl_is_sta : _GEN_8976; // @[rob.scala 411:{25,25}]
  wire  _GEN_8978 = 5'h1d == com_idx ? rob_uop_29_ctrl_is_sta : _GEN_8977; // @[rob.scala 411:{25,25}]
  wire  _GEN_8979 = 5'h1e == com_idx ? rob_uop_30_ctrl_is_sta : _GEN_8978; // @[rob.scala 411:{25,25}]
  wire  _GEN_8982 = 5'h1 == com_idx ? rob_uop_1_ctrl_is_load : rob_uop_0_ctrl_is_load; // @[rob.scala 411:{25,25}]
  wire  _GEN_8983 = 5'h2 == com_idx ? rob_uop_2_ctrl_is_load : _GEN_8982; // @[rob.scala 411:{25,25}]
  wire  _GEN_8984 = 5'h3 == com_idx ? rob_uop_3_ctrl_is_load : _GEN_8983; // @[rob.scala 411:{25,25}]
  wire  _GEN_8985 = 5'h4 == com_idx ? rob_uop_4_ctrl_is_load : _GEN_8984; // @[rob.scala 411:{25,25}]
  wire  _GEN_8986 = 5'h5 == com_idx ? rob_uop_5_ctrl_is_load : _GEN_8985; // @[rob.scala 411:{25,25}]
  wire  _GEN_8987 = 5'h6 == com_idx ? rob_uop_6_ctrl_is_load : _GEN_8986; // @[rob.scala 411:{25,25}]
  wire  _GEN_8988 = 5'h7 == com_idx ? rob_uop_7_ctrl_is_load : _GEN_8987; // @[rob.scala 411:{25,25}]
  wire  _GEN_8989 = 5'h8 == com_idx ? rob_uop_8_ctrl_is_load : _GEN_8988; // @[rob.scala 411:{25,25}]
  wire  _GEN_8990 = 5'h9 == com_idx ? rob_uop_9_ctrl_is_load : _GEN_8989; // @[rob.scala 411:{25,25}]
  wire  _GEN_8991 = 5'ha == com_idx ? rob_uop_10_ctrl_is_load : _GEN_8990; // @[rob.scala 411:{25,25}]
  wire  _GEN_8992 = 5'hb == com_idx ? rob_uop_11_ctrl_is_load : _GEN_8991; // @[rob.scala 411:{25,25}]
  wire  _GEN_8993 = 5'hc == com_idx ? rob_uop_12_ctrl_is_load : _GEN_8992; // @[rob.scala 411:{25,25}]
  wire  _GEN_8994 = 5'hd == com_idx ? rob_uop_13_ctrl_is_load : _GEN_8993; // @[rob.scala 411:{25,25}]
  wire  _GEN_8995 = 5'he == com_idx ? rob_uop_14_ctrl_is_load : _GEN_8994; // @[rob.scala 411:{25,25}]
  wire  _GEN_8996 = 5'hf == com_idx ? rob_uop_15_ctrl_is_load : _GEN_8995; // @[rob.scala 411:{25,25}]
  wire  _GEN_8997 = 5'h10 == com_idx ? rob_uop_16_ctrl_is_load : _GEN_8996; // @[rob.scala 411:{25,25}]
  wire  _GEN_8998 = 5'h11 == com_idx ? rob_uop_17_ctrl_is_load : _GEN_8997; // @[rob.scala 411:{25,25}]
  wire  _GEN_8999 = 5'h12 == com_idx ? rob_uop_18_ctrl_is_load : _GEN_8998; // @[rob.scala 411:{25,25}]
  wire  _GEN_9000 = 5'h13 == com_idx ? rob_uop_19_ctrl_is_load : _GEN_8999; // @[rob.scala 411:{25,25}]
  wire  _GEN_9001 = 5'h14 == com_idx ? rob_uop_20_ctrl_is_load : _GEN_9000; // @[rob.scala 411:{25,25}]
  wire  _GEN_9002 = 5'h15 == com_idx ? rob_uop_21_ctrl_is_load : _GEN_9001; // @[rob.scala 411:{25,25}]
  wire  _GEN_9003 = 5'h16 == com_idx ? rob_uop_22_ctrl_is_load : _GEN_9002; // @[rob.scala 411:{25,25}]
  wire  _GEN_9004 = 5'h17 == com_idx ? rob_uop_23_ctrl_is_load : _GEN_9003; // @[rob.scala 411:{25,25}]
  wire  _GEN_9005 = 5'h18 == com_idx ? rob_uop_24_ctrl_is_load : _GEN_9004; // @[rob.scala 411:{25,25}]
  wire  _GEN_9006 = 5'h19 == com_idx ? rob_uop_25_ctrl_is_load : _GEN_9005; // @[rob.scala 411:{25,25}]
  wire  _GEN_9007 = 5'h1a == com_idx ? rob_uop_26_ctrl_is_load : _GEN_9006; // @[rob.scala 411:{25,25}]
  wire  _GEN_9008 = 5'h1b == com_idx ? rob_uop_27_ctrl_is_load : _GEN_9007; // @[rob.scala 411:{25,25}]
  wire  _GEN_9009 = 5'h1c == com_idx ? rob_uop_28_ctrl_is_load : _GEN_9008; // @[rob.scala 411:{25,25}]
  wire  _GEN_9010 = 5'h1d == com_idx ? rob_uop_29_ctrl_is_load : _GEN_9009; // @[rob.scala 411:{25,25}]
  wire  _GEN_9011 = 5'h1e == com_idx ? rob_uop_30_ctrl_is_load : _GEN_9010; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9014 = 5'h1 == com_idx ? rob_uop_1_ctrl_csr_cmd : rob_uop_0_ctrl_csr_cmd; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9015 = 5'h2 == com_idx ? rob_uop_2_ctrl_csr_cmd : _GEN_9014; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9016 = 5'h3 == com_idx ? rob_uop_3_ctrl_csr_cmd : _GEN_9015; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9017 = 5'h4 == com_idx ? rob_uop_4_ctrl_csr_cmd : _GEN_9016; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9018 = 5'h5 == com_idx ? rob_uop_5_ctrl_csr_cmd : _GEN_9017; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9019 = 5'h6 == com_idx ? rob_uop_6_ctrl_csr_cmd : _GEN_9018; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9020 = 5'h7 == com_idx ? rob_uop_7_ctrl_csr_cmd : _GEN_9019; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9021 = 5'h8 == com_idx ? rob_uop_8_ctrl_csr_cmd : _GEN_9020; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9022 = 5'h9 == com_idx ? rob_uop_9_ctrl_csr_cmd : _GEN_9021; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9023 = 5'ha == com_idx ? rob_uop_10_ctrl_csr_cmd : _GEN_9022; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9024 = 5'hb == com_idx ? rob_uop_11_ctrl_csr_cmd : _GEN_9023; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9025 = 5'hc == com_idx ? rob_uop_12_ctrl_csr_cmd : _GEN_9024; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9026 = 5'hd == com_idx ? rob_uop_13_ctrl_csr_cmd : _GEN_9025; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9027 = 5'he == com_idx ? rob_uop_14_ctrl_csr_cmd : _GEN_9026; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9028 = 5'hf == com_idx ? rob_uop_15_ctrl_csr_cmd : _GEN_9027; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9029 = 5'h10 == com_idx ? rob_uop_16_ctrl_csr_cmd : _GEN_9028; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9030 = 5'h11 == com_idx ? rob_uop_17_ctrl_csr_cmd : _GEN_9029; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9031 = 5'h12 == com_idx ? rob_uop_18_ctrl_csr_cmd : _GEN_9030; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9032 = 5'h13 == com_idx ? rob_uop_19_ctrl_csr_cmd : _GEN_9031; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9033 = 5'h14 == com_idx ? rob_uop_20_ctrl_csr_cmd : _GEN_9032; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9034 = 5'h15 == com_idx ? rob_uop_21_ctrl_csr_cmd : _GEN_9033; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9035 = 5'h16 == com_idx ? rob_uop_22_ctrl_csr_cmd : _GEN_9034; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9036 = 5'h17 == com_idx ? rob_uop_23_ctrl_csr_cmd : _GEN_9035; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9037 = 5'h18 == com_idx ? rob_uop_24_ctrl_csr_cmd : _GEN_9036; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9038 = 5'h19 == com_idx ? rob_uop_25_ctrl_csr_cmd : _GEN_9037; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9039 = 5'h1a == com_idx ? rob_uop_26_ctrl_csr_cmd : _GEN_9038; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9040 = 5'h1b == com_idx ? rob_uop_27_ctrl_csr_cmd : _GEN_9039; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9041 = 5'h1c == com_idx ? rob_uop_28_ctrl_csr_cmd : _GEN_9040; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9042 = 5'h1d == com_idx ? rob_uop_29_ctrl_csr_cmd : _GEN_9041; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9043 = 5'h1e == com_idx ? rob_uop_30_ctrl_csr_cmd : _GEN_9042; // @[rob.scala 411:{25,25}]
  wire  _GEN_9046 = 5'h1 == com_idx ? rob_uop_1_ctrl_fcn_dw : rob_uop_0_ctrl_fcn_dw; // @[rob.scala 411:{25,25}]
  wire  _GEN_9047 = 5'h2 == com_idx ? rob_uop_2_ctrl_fcn_dw : _GEN_9046; // @[rob.scala 411:{25,25}]
  wire  _GEN_9048 = 5'h3 == com_idx ? rob_uop_3_ctrl_fcn_dw : _GEN_9047; // @[rob.scala 411:{25,25}]
  wire  _GEN_9049 = 5'h4 == com_idx ? rob_uop_4_ctrl_fcn_dw : _GEN_9048; // @[rob.scala 411:{25,25}]
  wire  _GEN_9050 = 5'h5 == com_idx ? rob_uop_5_ctrl_fcn_dw : _GEN_9049; // @[rob.scala 411:{25,25}]
  wire  _GEN_9051 = 5'h6 == com_idx ? rob_uop_6_ctrl_fcn_dw : _GEN_9050; // @[rob.scala 411:{25,25}]
  wire  _GEN_9052 = 5'h7 == com_idx ? rob_uop_7_ctrl_fcn_dw : _GEN_9051; // @[rob.scala 411:{25,25}]
  wire  _GEN_9053 = 5'h8 == com_idx ? rob_uop_8_ctrl_fcn_dw : _GEN_9052; // @[rob.scala 411:{25,25}]
  wire  _GEN_9054 = 5'h9 == com_idx ? rob_uop_9_ctrl_fcn_dw : _GEN_9053; // @[rob.scala 411:{25,25}]
  wire  _GEN_9055 = 5'ha == com_idx ? rob_uop_10_ctrl_fcn_dw : _GEN_9054; // @[rob.scala 411:{25,25}]
  wire  _GEN_9056 = 5'hb == com_idx ? rob_uop_11_ctrl_fcn_dw : _GEN_9055; // @[rob.scala 411:{25,25}]
  wire  _GEN_9057 = 5'hc == com_idx ? rob_uop_12_ctrl_fcn_dw : _GEN_9056; // @[rob.scala 411:{25,25}]
  wire  _GEN_9058 = 5'hd == com_idx ? rob_uop_13_ctrl_fcn_dw : _GEN_9057; // @[rob.scala 411:{25,25}]
  wire  _GEN_9059 = 5'he == com_idx ? rob_uop_14_ctrl_fcn_dw : _GEN_9058; // @[rob.scala 411:{25,25}]
  wire  _GEN_9060 = 5'hf == com_idx ? rob_uop_15_ctrl_fcn_dw : _GEN_9059; // @[rob.scala 411:{25,25}]
  wire  _GEN_9061 = 5'h10 == com_idx ? rob_uop_16_ctrl_fcn_dw : _GEN_9060; // @[rob.scala 411:{25,25}]
  wire  _GEN_9062 = 5'h11 == com_idx ? rob_uop_17_ctrl_fcn_dw : _GEN_9061; // @[rob.scala 411:{25,25}]
  wire  _GEN_9063 = 5'h12 == com_idx ? rob_uop_18_ctrl_fcn_dw : _GEN_9062; // @[rob.scala 411:{25,25}]
  wire  _GEN_9064 = 5'h13 == com_idx ? rob_uop_19_ctrl_fcn_dw : _GEN_9063; // @[rob.scala 411:{25,25}]
  wire  _GEN_9065 = 5'h14 == com_idx ? rob_uop_20_ctrl_fcn_dw : _GEN_9064; // @[rob.scala 411:{25,25}]
  wire  _GEN_9066 = 5'h15 == com_idx ? rob_uop_21_ctrl_fcn_dw : _GEN_9065; // @[rob.scala 411:{25,25}]
  wire  _GEN_9067 = 5'h16 == com_idx ? rob_uop_22_ctrl_fcn_dw : _GEN_9066; // @[rob.scala 411:{25,25}]
  wire  _GEN_9068 = 5'h17 == com_idx ? rob_uop_23_ctrl_fcn_dw : _GEN_9067; // @[rob.scala 411:{25,25}]
  wire  _GEN_9069 = 5'h18 == com_idx ? rob_uop_24_ctrl_fcn_dw : _GEN_9068; // @[rob.scala 411:{25,25}]
  wire  _GEN_9070 = 5'h19 == com_idx ? rob_uop_25_ctrl_fcn_dw : _GEN_9069; // @[rob.scala 411:{25,25}]
  wire  _GEN_9071 = 5'h1a == com_idx ? rob_uop_26_ctrl_fcn_dw : _GEN_9070; // @[rob.scala 411:{25,25}]
  wire  _GEN_9072 = 5'h1b == com_idx ? rob_uop_27_ctrl_fcn_dw : _GEN_9071; // @[rob.scala 411:{25,25}]
  wire  _GEN_9073 = 5'h1c == com_idx ? rob_uop_28_ctrl_fcn_dw : _GEN_9072; // @[rob.scala 411:{25,25}]
  wire  _GEN_9074 = 5'h1d == com_idx ? rob_uop_29_ctrl_fcn_dw : _GEN_9073; // @[rob.scala 411:{25,25}]
  wire  _GEN_9075 = 5'h1e == com_idx ? rob_uop_30_ctrl_fcn_dw : _GEN_9074; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9078 = 5'h1 == com_idx ? rob_uop_1_ctrl_op_fcn : rob_uop_0_ctrl_op_fcn; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9079 = 5'h2 == com_idx ? rob_uop_2_ctrl_op_fcn : _GEN_9078; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9080 = 5'h3 == com_idx ? rob_uop_3_ctrl_op_fcn : _GEN_9079; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9081 = 5'h4 == com_idx ? rob_uop_4_ctrl_op_fcn : _GEN_9080; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9082 = 5'h5 == com_idx ? rob_uop_5_ctrl_op_fcn : _GEN_9081; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9083 = 5'h6 == com_idx ? rob_uop_6_ctrl_op_fcn : _GEN_9082; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9084 = 5'h7 == com_idx ? rob_uop_7_ctrl_op_fcn : _GEN_9083; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9085 = 5'h8 == com_idx ? rob_uop_8_ctrl_op_fcn : _GEN_9084; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9086 = 5'h9 == com_idx ? rob_uop_9_ctrl_op_fcn : _GEN_9085; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9087 = 5'ha == com_idx ? rob_uop_10_ctrl_op_fcn : _GEN_9086; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9088 = 5'hb == com_idx ? rob_uop_11_ctrl_op_fcn : _GEN_9087; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9089 = 5'hc == com_idx ? rob_uop_12_ctrl_op_fcn : _GEN_9088; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9090 = 5'hd == com_idx ? rob_uop_13_ctrl_op_fcn : _GEN_9089; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9091 = 5'he == com_idx ? rob_uop_14_ctrl_op_fcn : _GEN_9090; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9092 = 5'hf == com_idx ? rob_uop_15_ctrl_op_fcn : _GEN_9091; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9093 = 5'h10 == com_idx ? rob_uop_16_ctrl_op_fcn : _GEN_9092; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9094 = 5'h11 == com_idx ? rob_uop_17_ctrl_op_fcn : _GEN_9093; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9095 = 5'h12 == com_idx ? rob_uop_18_ctrl_op_fcn : _GEN_9094; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9096 = 5'h13 == com_idx ? rob_uop_19_ctrl_op_fcn : _GEN_9095; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9097 = 5'h14 == com_idx ? rob_uop_20_ctrl_op_fcn : _GEN_9096; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9098 = 5'h15 == com_idx ? rob_uop_21_ctrl_op_fcn : _GEN_9097; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9099 = 5'h16 == com_idx ? rob_uop_22_ctrl_op_fcn : _GEN_9098; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9100 = 5'h17 == com_idx ? rob_uop_23_ctrl_op_fcn : _GEN_9099; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9101 = 5'h18 == com_idx ? rob_uop_24_ctrl_op_fcn : _GEN_9100; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9102 = 5'h19 == com_idx ? rob_uop_25_ctrl_op_fcn : _GEN_9101; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9103 = 5'h1a == com_idx ? rob_uop_26_ctrl_op_fcn : _GEN_9102; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9104 = 5'h1b == com_idx ? rob_uop_27_ctrl_op_fcn : _GEN_9103; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9105 = 5'h1c == com_idx ? rob_uop_28_ctrl_op_fcn : _GEN_9104; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9106 = 5'h1d == com_idx ? rob_uop_29_ctrl_op_fcn : _GEN_9105; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9107 = 5'h1e == com_idx ? rob_uop_30_ctrl_op_fcn : _GEN_9106; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9110 = 5'h1 == com_idx ? rob_uop_1_ctrl_imm_sel : rob_uop_0_ctrl_imm_sel; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9111 = 5'h2 == com_idx ? rob_uop_2_ctrl_imm_sel : _GEN_9110; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9112 = 5'h3 == com_idx ? rob_uop_3_ctrl_imm_sel : _GEN_9111; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9113 = 5'h4 == com_idx ? rob_uop_4_ctrl_imm_sel : _GEN_9112; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9114 = 5'h5 == com_idx ? rob_uop_5_ctrl_imm_sel : _GEN_9113; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9115 = 5'h6 == com_idx ? rob_uop_6_ctrl_imm_sel : _GEN_9114; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9116 = 5'h7 == com_idx ? rob_uop_7_ctrl_imm_sel : _GEN_9115; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9117 = 5'h8 == com_idx ? rob_uop_8_ctrl_imm_sel : _GEN_9116; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9118 = 5'h9 == com_idx ? rob_uop_9_ctrl_imm_sel : _GEN_9117; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9119 = 5'ha == com_idx ? rob_uop_10_ctrl_imm_sel : _GEN_9118; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9120 = 5'hb == com_idx ? rob_uop_11_ctrl_imm_sel : _GEN_9119; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9121 = 5'hc == com_idx ? rob_uop_12_ctrl_imm_sel : _GEN_9120; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9122 = 5'hd == com_idx ? rob_uop_13_ctrl_imm_sel : _GEN_9121; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9123 = 5'he == com_idx ? rob_uop_14_ctrl_imm_sel : _GEN_9122; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9124 = 5'hf == com_idx ? rob_uop_15_ctrl_imm_sel : _GEN_9123; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9125 = 5'h10 == com_idx ? rob_uop_16_ctrl_imm_sel : _GEN_9124; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9126 = 5'h11 == com_idx ? rob_uop_17_ctrl_imm_sel : _GEN_9125; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9127 = 5'h12 == com_idx ? rob_uop_18_ctrl_imm_sel : _GEN_9126; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9128 = 5'h13 == com_idx ? rob_uop_19_ctrl_imm_sel : _GEN_9127; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9129 = 5'h14 == com_idx ? rob_uop_20_ctrl_imm_sel : _GEN_9128; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9130 = 5'h15 == com_idx ? rob_uop_21_ctrl_imm_sel : _GEN_9129; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9131 = 5'h16 == com_idx ? rob_uop_22_ctrl_imm_sel : _GEN_9130; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9132 = 5'h17 == com_idx ? rob_uop_23_ctrl_imm_sel : _GEN_9131; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9133 = 5'h18 == com_idx ? rob_uop_24_ctrl_imm_sel : _GEN_9132; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9134 = 5'h19 == com_idx ? rob_uop_25_ctrl_imm_sel : _GEN_9133; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9135 = 5'h1a == com_idx ? rob_uop_26_ctrl_imm_sel : _GEN_9134; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9136 = 5'h1b == com_idx ? rob_uop_27_ctrl_imm_sel : _GEN_9135; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9137 = 5'h1c == com_idx ? rob_uop_28_ctrl_imm_sel : _GEN_9136; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9138 = 5'h1d == com_idx ? rob_uop_29_ctrl_imm_sel : _GEN_9137; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9139 = 5'h1e == com_idx ? rob_uop_30_ctrl_imm_sel : _GEN_9138; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9142 = 5'h1 == com_idx ? rob_uop_1_ctrl_op2_sel : rob_uop_0_ctrl_op2_sel; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9143 = 5'h2 == com_idx ? rob_uop_2_ctrl_op2_sel : _GEN_9142; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9144 = 5'h3 == com_idx ? rob_uop_3_ctrl_op2_sel : _GEN_9143; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9145 = 5'h4 == com_idx ? rob_uop_4_ctrl_op2_sel : _GEN_9144; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9146 = 5'h5 == com_idx ? rob_uop_5_ctrl_op2_sel : _GEN_9145; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9147 = 5'h6 == com_idx ? rob_uop_6_ctrl_op2_sel : _GEN_9146; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9148 = 5'h7 == com_idx ? rob_uop_7_ctrl_op2_sel : _GEN_9147; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9149 = 5'h8 == com_idx ? rob_uop_8_ctrl_op2_sel : _GEN_9148; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9150 = 5'h9 == com_idx ? rob_uop_9_ctrl_op2_sel : _GEN_9149; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9151 = 5'ha == com_idx ? rob_uop_10_ctrl_op2_sel : _GEN_9150; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9152 = 5'hb == com_idx ? rob_uop_11_ctrl_op2_sel : _GEN_9151; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9153 = 5'hc == com_idx ? rob_uop_12_ctrl_op2_sel : _GEN_9152; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9154 = 5'hd == com_idx ? rob_uop_13_ctrl_op2_sel : _GEN_9153; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9155 = 5'he == com_idx ? rob_uop_14_ctrl_op2_sel : _GEN_9154; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9156 = 5'hf == com_idx ? rob_uop_15_ctrl_op2_sel : _GEN_9155; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9157 = 5'h10 == com_idx ? rob_uop_16_ctrl_op2_sel : _GEN_9156; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9158 = 5'h11 == com_idx ? rob_uop_17_ctrl_op2_sel : _GEN_9157; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9159 = 5'h12 == com_idx ? rob_uop_18_ctrl_op2_sel : _GEN_9158; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9160 = 5'h13 == com_idx ? rob_uop_19_ctrl_op2_sel : _GEN_9159; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9161 = 5'h14 == com_idx ? rob_uop_20_ctrl_op2_sel : _GEN_9160; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9162 = 5'h15 == com_idx ? rob_uop_21_ctrl_op2_sel : _GEN_9161; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9163 = 5'h16 == com_idx ? rob_uop_22_ctrl_op2_sel : _GEN_9162; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9164 = 5'h17 == com_idx ? rob_uop_23_ctrl_op2_sel : _GEN_9163; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9165 = 5'h18 == com_idx ? rob_uop_24_ctrl_op2_sel : _GEN_9164; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9166 = 5'h19 == com_idx ? rob_uop_25_ctrl_op2_sel : _GEN_9165; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9167 = 5'h1a == com_idx ? rob_uop_26_ctrl_op2_sel : _GEN_9166; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9168 = 5'h1b == com_idx ? rob_uop_27_ctrl_op2_sel : _GEN_9167; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9169 = 5'h1c == com_idx ? rob_uop_28_ctrl_op2_sel : _GEN_9168; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9170 = 5'h1d == com_idx ? rob_uop_29_ctrl_op2_sel : _GEN_9169; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9171 = 5'h1e == com_idx ? rob_uop_30_ctrl_op2_sel : _GEN_9170; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9174 = 5'h1 == com_idx ? rob_uop_1_ctrl_op1_sel : rob_uop_0_ctrl_op1_sel; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9175 = 5'h2 == com_idx ? rob_uop_2_ctrl_op1_sel : _GEN_9174; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9176 = 5'h3 == com_idx ? rob_uop_3_ctrl_op1_sel : _GEN_9175; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9177 = 5'h4 == com_idx ? rob_uop_4_ctrl_op1_sel : _GEN_9176; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9178 = 5'h5 == com_idx ? rob_uop_5_ctrl_op1_sel : _GEN_9177; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9179 = 5'h6 == com_idx ? rob_uop_6_ctrl_op1_sel : _GEN_9178; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9180 = 5'h7 == com_idx ? rob_uop_7_ctrl_op1_sel : _GEN_9179; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9181 = 5'h8 == com_idx ? rob_uop_8_ctrl_op1_sel : _GEN_9180; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9182 = 5'h9 == com_idx ? rob_uop_9_ctrl_op1_sel : _GEN_9181; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9183 = 5'ha == com_idx ? rob_uop_10_ctrl_op1_sel : _GEN_9182; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9184 = 5'hb == com_idx ? rob_uop_11_ctrl_op1_sel : _GEN_9183; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9185 = 5'hc == com_idx ? rob_uop_12_ctrl_op1_sel : _GEN_9184; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9186 = 5'hd == com_idx ? rob_uop_13_ctrl_op1_sel : _GEN_9185; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9187 = 5'he == com_idx ? rob_uop_14_ctrl_op1_sel : _GEN_9186; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9188 = 5'hf == com_idx ? rob_uop_15_ctrl_op1_sel : _GEN_9187; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9189 = 5'h10 == com_idx ? rob_uop_16_ctrl_op1_sel : _GEN_9188; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9190 = 5'h11 == com_idx ? rob_uop_17_ctrl_op1_sel : _GEN_9189; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9191 = 5'h12 == com_idx ? rob_uop_18_ctrl_op1_sel : _GEN_9190; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9192 = 5'h13 == com_idx ? rob_uop_19_ctrl_op1_sel : _GEN_9191; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9193 = 5'h14 == com_idx ? rob_uop_20_ctrl_op1_sel : _GEN_9192; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9194 = 5'h15 == com_idx ? rob_uop_21_ctrl_op1_sel : _GEN_9193; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9195 = 5'h16 == com_idx ? rob_uop_22_ctrl_op1_sel : _GEN_9194; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9196 = 5'h17 == com_idx ? rob_uop_23_ctrl_op1_sel : _GEN_9195; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9197 = 5'h18 == com_idx ? rob_uop_24_ctrl_op1_sel : _GEN_9196; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9198 = 5'h19 == com_idx ? rob_uop_25_ctrl_op1_sel : _GEN_9197; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9199 = 5'h1a == com_idx ? rob_uop_26_ctrl_op1_sel : _GEN_9198; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9200 = 5'h1b == com_idx ? rob_uop_27_ctrl_op1_sel : _GEN_9199; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9201 = 5'h1c == com_idx ? rob_uop_28_ctrl_op1_sel : _GEN_9200; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9202 = 5'h1d == com_idx ? rob_uop_29_ctrl_op1_sel : _GEN_9201; // @[rob.scala 411:{25,25}]
  wire [1:0] _GEN_9203 = 5'h1e == com_idx ? rob_uop_30_ctrl_op1_sel : _GEN_9202; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9206 = 5'h1 == com_idx ? rob_uop_1_ctrl_br_type : rob_uop_0_ctrl_br_type; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9207 = 5'h2 == com_idx ? rob_uop_2_ctrl_br_type : _GEN_9206; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9208 = 5'h3 == com_idx ? rob_uop_3_ctrl_br_type : _GEN_9207; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9209 = 5'h4 == com_idx ? rob_uop_4_ctrl_br_type : _GEN_9208; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9210 = 5'h5 == com_idx ? rob_uop_5_ctrl_br_type : _GEN_9209; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9211 = 5'h6 == com_idx ? rob_uop_6_ctrl_br_type : _GEN_9210; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9212 = 5'h7 == com_idx ? rob_uop_7_ctrl_br_type : _GEN_9211; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9213 = 5'h8 == com_idx ? rob_uop_8_ctrl_br_type : _GEN_9212; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9214 = 5'h9 == com_idx ? rob_uop_9_ctrl_br_type : _GEN_9213; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9215 = 5'ha == com_idx ? rob_uop_10_ctrl_br_type : _GEN_9214; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9216 = 5'hb == com_idx ? rob_uop_11_ctrl_br_type : _GEN_9215; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9217 = 5'hc == com_idx ? rob_uop_12_ctrl_br_type : _GEN_9216; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9218 = 5'hd == com_idx ? rob_uop_13_ctrl_br_type : _GEN_9217; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9219 = 5'he == com_idx ? rob_uop_14_ctrl_br_type : _GEN_9218; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9220 = 5'hf == com_idx ? rob_uop_15_ctrl_br_type : _GEN_9219; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9221 = 5'h10 == com_idx ? rob_uop_16_ctrl_br_type : _GEN_9220; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9222 = 5'h11 == com_idx ? rob_uop_17_ctrl_br_type : _GEN_9221; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9223 = 5'h12 == com_idx ? rob_uop_18_ctrl_br_type : _GEN_9222; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9224 = 5'h13 == com_idx ? rob_uop_19_ctrl_br_type : _GEN_9223; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9225 = 5'h14 == com_idx ? rob_uop_20_ctrl_br_type : _GEN_9224; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9226 = 5'h15 == com_idx ? rob_uop_21_ctrl_br_type : _GEN_9225; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9227 = 5'h16 == com_idx ? rob_uop_22_ctrl_br_type : _GEN_9226; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9228 = 5'h17 == com_idx ? rob_uop_23_ctrl_br_type : _GEN_9227; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9229 = 5'h18 == com_idx ? rob_uop_24_ctrl_br_type : _GEN_9228; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9230 = 5'h19 == com_idx ? rob_uop_25_ctrl_br_type : _GEN_9229; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9231 = 5'h1a == com_idx ? rob_uop_26_ctrl_br_type : _GEN_9230; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9232 = 5'h1b == com_idx ? rob_uop_27_ctrl_br_type : _GEN_9231; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9233 = 5'h1c == com_idx ? rob_uop_28_ctrl_br_type : _GEN_9232; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9234 = 5'h1d == com_idx ? rob_uop_29_ctrl_br_type : _GEN_9233; // @[rob.scala 411:{25,25}]
  wire [3:0] _GEN_9235 = 5'h1e == com_idx ? rob_uop_30_ctrl_br_type : _GEN_9234; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9238 = 5'h1 == com_idx ? rob_uop_1_fu_code : rob_uop_0_fu_code; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9239 = 5'h2 == com_idx ? rob_uop_2_fu_code : _GEN_9238; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9240 = 5'h3 == com_idx ? rob_uop_3_fu_code : _GEN_9239; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9241 = 5'h4 == com_idx ? rob_uop_4_fu_code : _GEN_9240; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9242 = 5'h5 == com_idx ? rob_uop_5_fu_code : _GEN_9241; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9243 = 5'h6 == com_idx ? rob_uop_6_fu_code : _GEN_9242; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9244 = 5'h7 == com_idx ? rob_uop_7_fu_code : _GEN_9243; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9245 = 5'h8 == com_idx ? rob_uop_8_fu_code : _GEN_9244; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9246 = 5'h9 == com_idx ? rob_uop_9_fu_code : _GEN_9245; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9247 = 5'ha == com_idx ? rob_uop_10_fu_code : _GEN_9246; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9248 = 5'hb == com_idx ? rob_uop_11_fu_code : _GEN_9247; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9249 = 5'hc == com_idx ? rob_uop_12_fu_code : _GEN_9248; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9250 = 5'hd == com_idx ? rob_uop_13_fu_code : _GEN_9249; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9251 = 5'he == com_idx ? rob_uop_14_fu_code : _GEN_9250; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9252 = 5'hf == com_idx ? rob_uop_15_fu_code : _GEN_9251; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9253 = 5'h10 == com_idx ? rob_uop_16_fu_code : _GEN_9252; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9254 = 5'h11 == com_idx ? rob_uop_17_fu_code : _GEN_9253; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9255 = 5'h12 == com_idx ? rob_uop_18_fu_code : _GEN_9254; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9256 = 5'h13 == com_idx ? rob_uop_19_fu_code : _GEN_9255; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9257 = 5'h14 == com_idx ? rob_uop_20_fu_code : _GEN_9256; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9258 = 5'h15 == com_idx ? rob_uop_21_fu_code : _GEN_9257; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9259 = 5'h16 == com_idx ? rob_uop_22_fu_code : _GEN_9258; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9260 = 5'h17 == com_idx ? rob_uop_23_fu_code : _GEN_9259; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9261 = 5'h18 == com_idx ? rob_uop_24_fu_code : _GEN_9260; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9262 = 5'h19 == com_idx ? rob_uop_25_fu_code : _GEN_9261; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9263 = 5'h1a == com_idx ? rob_uop_26_fu_code : _GEN_9262; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9264 = 5'h1b == com_idx ? rob_uop_27_fu_code : _GEN_9263; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9265 = 5'h1c == com_idx ? rob_uop_28_fu_code : _GEN_9264; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9266 = 5'h1d == com_idx ? rob_uop_29_fu_code : _GEN_9265; // @[rob.scala 411:{25,25}]
  wire [9:0] _GEN_9267 = 5'h1e == com_idx ? rob_uop_30_fu_code : _GEN_9266; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9270 = 5'h1 == com_idx ? rob_uop_1_iq_type : rob_uop_0_iq_type; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9271 = 5'h2 == com_idx ? rob_uop_2_iq_type : _GEN_9270; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9272 = 5'h3 == com_idx ? rob_uop_3_iq_type : _GEN_9271; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9273 = 5'h4 == com_idx ? rob_uop_4_iq_type : _GEN_9272; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9274 = 5'h5 == com_idx ? rob_uop_5_iq_type : _GEN_9273; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9275 = 5'h6 == com_idx ? rob_uop_6_iq_type : _GEN_9274; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9276 = 5'h7 == com_idx ? rob_uop_7_iq_type : _GEN_9275; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9277 = 5'h8 == com_idx ? rob_uop_8_iq_type : _GEN_9276; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9278 = 5'h9 == com_idx ? rob_uop_9_iq_type : _GEN_9277; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9279 = 5'ha == com_idx ? rob_uop_10_iq_type : _GEN_9278; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9280 = 5'hb == com_idx ? rob_uop_11_iq_type : _GEN_9279; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9281 = 5'hc == com_idx ? rob_uop_12_iq_type : _GEN_9280; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9282 = 5'hd == com_idx ? rob_uop_13_iq_type : _GEN_9281; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9283 = 5'he == com_idx ? rob_uop_14_iq_type : _GEN_9282; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9284 = 5'hf == com_idx ? rob_uop_15_iq_type : _GEN_9283; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9285 = 5'h10 == com_idx ? rob_uop_16_iq_type : _GEN_9284; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9286 = 5'h11 == com_idx ? rob_uop_17_iq_type : _GEN_9285; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9287 = 5'h12 == com_idx ? rob_uop_18_iq_type : _GEN_9286; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9288 = 5'h13 == com_idx ? rob_uop_19_iq_type : _GEN_9287; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9289 = 5'h14 == com_idx ? rob_uop_20_iq_type : _GEN_9288; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9290 = 5'h15 == com_idx ? rob_uop_21_iq_type : _GEN_9289; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9291 = 5'h16 == com_idx ? rob_uop_22_iq_type : _GEN_9290; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9292 = 5'h17 == com_idx ? rob_uop_23_iq_type : _GEN_9291; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9293 = 5'h18 == com_idx ? rob_uop_24_iq_type : _GEN_9292; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9294 = 5'h19 == com_idx ? rob_uop_25_iq_type : _GEN_9293; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9295 = 5'h1a == com_idx ? rob_uop_26_iq_type : _GEN_9294; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9296 = 5'h1b == com_idx ? rob_uop_27_iq_type : _GEN_9295; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9297 = 5'h1c == com_idx ? rob_uop_28_iq_type : _GEN_9296; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9298 = 5'h1d == com_idx ? rob_uop_29_iq_type : _GEN_9297; // @[rob.scala 411:{25,25}]
  wire [2:0] _GEN_9299 = 5'h1e == com_idx ? rob_uop_30_iq_type : _GEN_9298; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9302 = 5'h1 == com_idx ? rob_uop_1_debug_pc : rob_uop_0_debug_pc; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9303 = 5'h2 == com_idx ? rob_uop_2_debug_pc : _GEN_9302; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9304 = 5'h3 == com_idx ? rob_uop_3_debug_pc : _GEN_9303; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9305 = 5'h4 == com_idx ? rob_uop_4_debug_pc : _GEN_9304; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9306 = 5'h5 == com_idx ? rob_uop_5_debug_pc : _GEN_9305; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9307 = 5'h6 == com_idx ? rob_uop_6_debug_pc : _GEN_9306; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9308 = 5'h7 == com_idx ? rob_uop_7_debug_pc : _GEN_9307; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9309 = 5'h8 == com_idx ? rob_uop_8_debug_pc : _GEN_9308; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9310 = 5'h9 == com_idx ? rob_uop_9_debug_pc : _GEN_9309; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9311 = 5'ha == com_idx ? rob_uop_10_debug_pc : _GEN_9310; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9312 = 5'hb == com_idx ? rob_uop_11_debug_pc : _GEN_9311; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9313 = 5'hc == com_idx ? rob_uop_12_debug_pc : _GEN_9312; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9314 = 5'hd == com_idx ? rob_uop_13_debug_pc : _GEN_9313; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9315 = 5'he == com_idx ? rob_uop_14_debug_pc : _GEN_9314; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9316 = 5'hf == com_idx ? rob_uop_15_debug_pc : _GEN_9315; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9317 = 5'h10 == com_idx ? rob_uop_16_debug_pc : _GEN_9316; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9318 = 5'h11 == com_idx ? rob_uop_17_debug_pc : _GEN_9317; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9319 = 5'h12 == com_idx ? rob_uop_18_debug_pc : _GEN_9318; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9320 = 5'h13 == com_idx ? rob_uop_19_debug_pc : _GEN_9319; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9321 = 5'h14 == com_idx ? rob_uop_20_debug_pc : _GEN_9320; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9322 = 5'h15 == com_idx ? rob_uop_21_debug_pc : _GEN_9321; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9323 = 5'h16 == com_idx ? rob_uop_22_debug_pc : _GEN_9322; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9324 = 5'h17 == com_idx ? rob_uop_23_debug_pc : _GEN_9323; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9325 = 5'h18 == com_idx ? rob_uop_24_debug_pc : _GEN_9324; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9326 = 5'h19 == com_idx ? rob_uop_25_debug_pc : _GEN_9325; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9327 = 5'h1a == com_idx ? rob_uop_26_debug_pc : _GEN_9326; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9328 = 5'h1b == com_idx ? rob_uop_27_debug_pc : _GEN_9327; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9329 = 5'h1c == com_idx ? rob_uop_28_debug_pc : _GEN_9328; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9330 = 5'h1d == com_idx ? rob_uop_29_debug_pc : _GEN_9329; // @[rob.scala 411:{25,25}]
  wire [39:0] _GEN_9331 = 5'h1e == com_idx ? rob_uop_30_debug_pc : _GEN_9330; // @[rob.scala 411:{25,25}]
  wire  _GEN_9334 = 5'h1 == com_idx ? rob_uop_1_is_rvc : rob_uop_0_is_rvc; // @[rob.scala 411:{25,25}]
  wire  _GEN_9335 = 5'h2 == com_idx ? rob_uop_2_is_rvc : _GEN_9334; // @[rob.scala 411:{25,25}]
  wire  _GEN_9336 = 5'h3 == com_idx ? rob_uop_3_is_rvc : _GEN_9335; // @[rob.scala 411:{25,25}]
  wire  _GEN_9337 = 5'h4 == com_idx ? rob_uop_4_is_rvc : _GEN_9336; // @[rob.scala 411:{25,25}]
  wire  _GEN_9338 = 5'h5 == com_idx ? rob_uop_5_is_rvc : _GEN_9337; // @[rob.scala 411:{25,25}]
  wire  _GEN_9339 = 5'h6 == com_idx ? rob_uop_6_is_rvc : _GEN_9338; // @[rob.scala 411:{25,25}]
  wire  _GEN_9340 = 5'h7 == com_idx ? rob_uop_7_is_rvc : _GEN_9339; // @[rob.scala 411:{25,25}]
  wire  _GEN_9341 = 5'h8 == com_idx ? rob_uop_8_is_rvc : _GEN_9340; // @[rob.scala 411:{25,25}]
  wire  _GEN_9342 = 5'h9 == com_idx ? rob_uop_9_is_rvc : _GEN_9341; // @[rob.scala 411:{25,25}]
  wire  _GEN_9343 = 5'ha == com_idx ? rob_uop_10_is_rvc : _GEN_9342; // @[rob.scala 411:{25,25}]
  wire  _GEN_9344 = 5'hb == com_idx ? rob_uop_11_is_rvc : _GEN_9343; // @[rob.scala 411:{25,25}]
  wire  _GEN_9345 = 5'hc == com_idx ? rob_uop_12_is_rvc : _GEN_9344; // @[rob.scala 411:{25,25}]
  wire  _GEN_9346 = 5'hd == com_idx ? rob_uop_13_is_rvc : _GEN_9345; // @[rob.scala 411:{25,25}]
  wire  _GEN_9347 = 5'he == com_idx ? rob_uop_14_is_rvc : _GEN_9346; // @[rob.scala 411:{25,25}]
  wire  _GEN_9348 = 5'hf == com_idx ? rob_uop_15_is_rvc : _GEN_9347; // @[rob.scala 411:{25,25}]
  wire  _GEN_9349 = 5'h10 == com_idx ? rob_uop_16_is_rvc : _GEN_9348; // @[rob.scala 411:{25,25}]
  wire  _GEN_9350 = 5'h11 == com_idx ? rob_uop_17_is_rvc : _GEN_9349; // @[rob.scala 411:{25,25}]
  wire  _GEN_9351 = 5'h12 == com_idx ? rob_uop_18_is_rvc : _GEN_9350; // @[rob.scala 411:{25,25}]
  wire  _GEN_9352 = 5'h13 == com_idx ? rob_uop_19_is_rvc : _GEN_9351; // @[rob.scala 411:{25,25}]
  wire  _GEN_9353 = 5'h14 == com_idx ? rob_uop_20_is_rvc : _GEN_9352; // @[rob.scala 411:{25,25}]
  wire  _GEN_9354 = 5'h15 == com_idx ? rob_uop_21_is_rvc : _GEN_9353; // @[rob.scala 411:{25,25}]
  wire  _GEN_9355 = 5'h16 == com_idx ? rob_uop_22_is_rvc : _GEN_9354; // @[rob.scala 411:{25,25}]
  wire  _GEN_9356 = 5'h17 == com_idx ? rob_uop_23_is_rvc : _GEN_9355; // @[rob.scala 411:{25,25}]
  wire  _GEN_9357 = 5'h18 == com_idx ? rob_uop_24_is_rvc : _GEN_9356; // @[rob.scala 411:{25,25}]
  wire  _GEN_9358 = 5'h19 == com_idx ? rob_uop_25_is_rvc : _GEN_9357; // @[rob.scala 411:{25,25}]
  wire  _GEN_9359 = 5'h1a == com_idx ? rob_uop_26_is_rvc : _GEN_9358; // @[rob.scala 411:{25,25}]
  wire  _GEN_9360 = 5'h1b == com_idx ? rob_uop_27_is_rvc : _GEN_9359; // @[rob.scala 411:{25,25}]
  wire  _GEN_9361 = 5'h1c == com_idx ? rob_uop_28_is_rvc : _GEN_9360; // @[rob.scala 411:{25,25}]
  wire  _GEN_9362 = 5'h1d == com_idx ? rob_uop_29_is_rvc : _GEN_9361; // @[rob.scala 411:{25,25}]
  wire  _GEN_9363 = 5'h1e == com_idx ? rob_uop_30_is_rvc : _GEN_9362; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9366 = 5'h1 == com_idx ? rob_uop_1_debug_inst : rob_uop_0_debug_inst; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9367 = 5'h2 == com_idx ? rob_uop_2_debug_inst : _GEN_9366; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9368 = 5'h3 == com_idx ? rob_uop_3_debug_inst : _GEN_9367; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9369 = 5'h4 == com_idx ? rob_uop_4_debug_inst : _GEN_9368; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9370 = 5'h5 == com_idx ? rob_uop_5_debug_inst : _GEN_9369; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9371 = 5'h6 == com_idx ? rob_uop_6_debug_inst : _GEN_9370; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9372 = 5'h7 == com_idx ? rob_uop_7_debug_inst : _GEN_9371; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9373 = 5'h8 == com_idx ? rob_uop_8_debug_inst : _GEN_9372; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9374 = 5'h9 == com_idx ? rob_uop_9_debug_inst : _GEN_9373; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9375 = 5'ha == com_idx ? rob_uop_10_debug_inst : _GEN_9374; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9376 = 5'hb == com_idx ? rob_uop_11_debug_inst : _GEN_9375; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9377 = 5'hc == com_idx ? rob_uop_12_debug_inst : _GEN_9376; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9378 = 5'hd == com_idx ? rob_uop_13_debug_inst : _GEN_9377; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9379 = 5'he == com_idx ? rob_uop_14_debug_inst : _GEN_9378; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9380 = 5'hf == com_idx ? rob_uop_15_debug_inst : _GEN_9379; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9381 = 5'h10 == com_idx ? rob_uop_16_debug_inst : _GEN_9380; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9382 = 5'h11 == com_idx ? rob_uop_17_debug_inst : _GEN_9381; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9383 = 5'h12 == com_idx ? rob_uop_18_debug_inst : _GEN_9382; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9384 = 5'h13 == com_idx ? rob_uop_19_debug_inst : _GEN_9383; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9385 = 5'h14 == com_idx ? rob_uop_20_debug_inst : _GEN_9384; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9386 = 5'h15 == com_idx ? rob_uop_21_debug_inst : _GEN_9385; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9387 = 5'h16 == com_idx ? rob_uop_22_debug_inst : _GEN_9386; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9388 = 5'h17 == com_idx ? rob_uop_23_debug_inst : _GEN_9387; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9389 = 5'h18 == com_idx ? rob_uop_24_debug_inst : _GEN_9388; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9390 = 5'h19 == com_idx ? rob_uop_25_debug_inst : _GEN_9389; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9391 = 5'h1a == com_idx ? rob_uop_26_debug_inst : _GEN_9390; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9392 = 5'h1b == com_idx ? rob_uop_27_debug_inst : _GEN_9391; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9393 = 5'h1c == com_idx ? rob_uop_28_debug_inst : _GEN_9392; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9394 = 5'h1d == com_idx ? rob_uop_29_debug_inst : _GEN_9393; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9395 = 5'h1e == com_idx ? rob_uop_30_debug_inst : _GEN_9394; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9398 = 5'h1 == com_idx ? rob_uop_1_inst : rob_uop_0_inst; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9399 = 5'h2 == com_idx ? rob_uop_2_inst : _GEN_9398; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9400 = 5'h3 == com_idx ? rob_uop_3_inst : _GEN_9399; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9401 = 5'h4 == com_idx ? rob_uop_4_inst : _GEN_9400; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9402 = 5'h5 == com_idx ? rob_uop_5_inst : _GEN_9401; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9403 = 5'h6 == com_idx ? rob_uop_6_inst : _GEN_9402; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9404 = 5'h7 == com_idx ? rob_uop_7_inst : _GEN_9403; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9405 = 5'h8 == com_idx ? rob_uop_8_inst : _GEN_9404; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9406 = 5'h9 == com_idx ? rob_uop_9_inst : _GEN_9405; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9407 = 5'ha == com_idx ? rob_uop_10_inst : _GEN_9406; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9408 = 5'hb == com_idx ? rob_uop_11_inst : _GEN_9407; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9409 = 5'hc == com_idx ? rob_uop_12_inst : _GEN_9408; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9410 = 5'hd == com_idx ? rob_uop_13_inst : _GEN_9409; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9411 = 5'he == com_idx ? rob_uop_14_inst : _GEN_9410; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9412 = 5'hf == com_idx ? rob_uop_15_inst : _GEN_9411; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9413 = 5'h10 == com_idx ? rob_uop_16_inst : _GEN_9412; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9414 = 5'h11 == com_idx ? rob_uop_17_inst : _GEN_9413; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9415 = 5'h12 == com_idx ? rob_uop_18_inst : _GEN_9414; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9416 = 5'h13 == com_idx ? rob_uop_19_inst : _GEN_9415; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9417 = 5'h14 == com_idx ? rob_uop_20_inst : _GEN_9416; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9418 = 5'h15 == com_idx ? rob_uop_21_inst : _GEN_9417; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9419 = 5'h16 == com_idx ? rob_uop_22_inst : _GEN_9418; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9420 = 5'h17 == com_idx ? rob_uop_23_inst : _GEN_9419; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9421 = 5'h18 == com_idx ? rob_uop_24_inst : _GEN_9420; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9422 = 5'h19 == com_idx ? rob_uop_25_inst : _GEN_9421; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9423 = 5'h1a == com_idx ? rob_uop_26_inst : _GEN_9422; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9424 = 5'h1b == com_idx ? rob_uop_27_inst : _GEN_9423; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9425 = 5'h1c == com_idx ? rob_uop_28_inst : _GEN_9424; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9426 = 5'h1d == com_idx ? rob_uop_29_inst : _GEN_9425; // @[rob.scala 411:{25,25}]
  wire [31:0] _GEN_9427 = 5'h1e == com_idx ? rob_uop_30_inst : _GEN_9426; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9430 = 5'h1 == com_idx ? rob_uop_1_uopc : rob_uop_0_uopc; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9431 = 5'h2 == com_idx ? rob_uop_2_uopc : _GEN_9430; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9432 = 5'h3 == com_idx ? rob_uop_3_uopc : _GEN_9431; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9433 = 5'h4 == com_idx ? rob_uop_4_uopc : _GEN_9432; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9434 = 5'h5 == com_idx ? rob_uop_5_uopc : _GEN_9433; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9435 = 5'h6 == com_idx ? rob_uop_6_uopc : _GEN_9434; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9436 = 5'h7 == com_idx ? rob_uop_7_uopc : _GEN_9435; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9437 = 5'h8 == com_idx ? rob_uop_8_uopc : _GEN_9436; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9438 = 5'h9 == com_idx ? rob_uop_9_uopc : _GEN_9437; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9439 = 5'ha == com_idx ? rob_uop_10_uopc : _GEN_9438; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9440 = 5'hb == com_idx ? rob_uop_11_uopc : _GEN_9439; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9441 = 5'hc == com_idx ? rob_uop_12_uopc : _GEN_9440; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9442 = 5'hd == com_idx ? rob_uop_13_uopc : _GEN_9441; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9443 = 5'he == com_idx ? rob_uop_14_uopc : _GEN_9442; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9444 = 5'hf == com_idx ? rob_uop_15_uopc : _GEN_9443; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9445 = 5'h10 == com_idx ? rob_uop_16_uopc : _GEN_9444; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9446 = 5'h11 == com_idx ? rob_uop_17_uopc : _GEN_9445; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9447 = 5'h12 == com_idx ? rob_uop_18_uopc : _GEN_9446; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9448 = 5'h13 == com_idx ? rob_uop_19_uopc : _GEN_9447; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9449 = 5'h14 == com_idx ? rob_uop_20_uopc : _GEN_9448; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9450 = 5'h15 == com_idx ? rob_uop_21_uopc : _GEN_9449; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9451 = 5'h16 == com_idx ? rob_uop_22_uopc : _GEN_9450; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9452 = 5'h17 == com_idx ? rob_uop_23_uopc : _GEN_9451; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9453 = 5'h18 == com_idx ? rob_uop_24_uopc : _GEN_9452; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9454 = 5'h19 == com_idx ? rob_uop_25_uopc : _GEN_9453; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9455 = 5'h1a == com_idx ? rob_uop_26_uopc : _GEN_9454; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9456 = 5'h1b == com_idx ? rob_uop_27_uopc : _GEN_9455; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9457 = 5'h1c == com_idx ? rob_uop_28_uopc : _GEN_9456; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9458 = 5'h1d == com_idx ? rob_uop_29_uopc : _GEN_9457; // @[rob.scala 411:{25,25}]
  wire [6:0] _GEN_9459 = 5'h1e == com_idx ? rob_uop_30_uopc : _GEN_9458; // @[rob.scala 411:{25,25}]
  wire  _T_78 = io_brupdate_b2_uop_rob_idx == com_idx; // @[rob.scala 418:45]
  wire  _T_79 = io_brupdate_b2_mispredict & _T_78; // @[rob.scala 417:57]
  wire  _T_597 = rob_tail == rob_head; // @[rob.scala 787:26]
  wire  full = rob_tail == rob_head & maybe_full; // @[rob.scala 787:39]
  wire  _T_81 = ~full; // @[rob.scala 425:47]
  wire  rbk_row = _T & ~full; // @[rob.scala 425:44]
  wire  _GEN_9464 = 5'h1 == com_idx ? rob_val_1 : rob_val_0; // @[rob.scala 427:{40,40}]
  wire  _GEN_9465 = 5'h2 == com_idx ? rob_val_2 : _GEN_9464; // @[rob.scala 427:{40,40}]
  wire  _GEN_9466 = 5'h3 == com_idx ? rob_val_3 : _GEN_9465; // @[rob.scala 427:{40,40}]
  wire  _GEN_9467 = 5'h4 == com_idx ? rob_val_4 : _GEN_9466; // @[rob.scala 427:{40,40}]
  wire  _GEN_9468 = 5'h5 == com_idx ? rob_val_5 : _GEN_9467; // @[rob.scala 427:{40,40}]
  wire  _GEN_9469 = 5'h6 == com_idx ? rob_val_6 : _GEN_9468; // @[rob.scala 427:{40,40}]
  wire  _GEN_9470 = 5'h7 == com_idx ? rob_val_7 : _GEN_9469; // @[rob.scala 427:{40,40}]
  wire  _GEN_9471 = 5'h8 == com_idx ? rob_val_8 : _GEN_9470; // @[rob.scala 427:{40,40}]
  wire  _GEN_9472 = 5'h9 == com_idx ? rob_val_9 : _GEN_9471; // @[rob.scala 427:{40,40}]
  wire  _GEN_9473 = 5'ha == com_idx ? rob_val_10 : _GEN_9472; // @[rob.scala 427:{40,40}]
  wire  _GEN_9474 = 5'hb == com_idx ? rob_val_11 : _GEN_9473; // @[rob.scala 427:{40,40}]
  wire  _GEN_9475 = 5'hc == com_idx ? rob_val_12 : _GEN_9474; // @[rob.scala 427:{40,40}]
  wire  _GEN_9476 = 5'hd == com_idx ? rob_val_13 : _GEN_9475; // @[rob.scala 427:{40,40}]
  wire  _GEN_9477 = 5'he == com_idx ? rob_val_14 : _GEN_9476; // @[rob.scala 427:{40,40}]
  wire  _GEN_9478 = 5'hf == com_idx ? rob_val_15 : _GEN_9477; // @[rob.scala 427:{40,40}]
  wire  _GEN_9479 = 5'h10 == com_idx ? rob_val_16 : _GEN_9478; // @[rob.scala 427:{40,40}]
  wire  _GEN_9480 = 5'h11 == com_idx ? rob_val_17 : _GEN_9479; // @[rob.scala 427:{40,40}]
  wire  _GEN_9481 = 5'h12 == com_idx ? rob_val_18 : _GEN_9480; // @[rob.scala 427:{40,40}]
  wire  _GEN_9482 = 5'h13 == com_idx ? rob_val_19 : _GEN_9481; // @[rob.scala 427:{40,40}]
  wire  _GEN_9483 = 5'h14 == com_idx ? rob_val_20 : _GEN_9482; // @[rob.scala 427:{40,40}]
  wire  _GEN_9484 = 5'h15 == com_idx ? rob_val_21 : _GEN_9483; // @[rob.scala 427:{40,40}]
  wire  _GEN_9485 = 5'h16 == com_idx ? rob_val_22 : _GEN_9484; // @[rob.scala 427:{40,40}]
  wire  _GEN_9486 = 5'h17 == com_idx ? rob_val_23 : _GEN_9485; // @[rob.scala 427:{40,40}]
  wire  _GEN_9487 = 5'h18 == com_idx ? rob_val_24 : _GEN_9486; // @[rob.scala 427:{40,40}]
  wire  _GEN_9488 = 5'h19 == com_idx ? rob_val_25 : _GEN_9487; // @[rob.scala 427:{40,40}]
  wire  _GEN_9489 = 5'h1a == com_idx ? rob_val_26 : _GEN_9488; // @[rob.scala 427:{40,40}]
  wire  _GEN_9490 = 5'h1b == com_idx ? rob_val_27 : _GEN_9489; // @[rob.scala 427:{40,40}]
  wire  _GEN_9491 = 5'h1c == com_idx ? rob_val_28 : _GEN_9490; // @[rob.scala 427:{40,40}]
  wire  _GEN_9492 = 5'h1d == com_idx ? rob_val_29 : _GEN_9491; // @[rob.scala 427:{40,40}]
  wire  _GEN_9493 = 5'h1e == com_idx ? rob_val_30 : _GEN_9492; // @[rob.scala 427:{40,40}]
  wire  _GEN_9494 = 5'h1f == com_idx ? rob_val_31 : _GEN_9493; // @[rob.scala 427:{40,40}]
  wire  _GEN_9495 = 5'h0 == com_idx ? 1'h0 : _GEN_2790; // @[rob.scala 434:{30,30}]
  wire  _GEN_9496 = 5'h1 == com_idx ? 1'h0 : _GEN_2791; // @[rob.scala 434:{30,30}]
  wire  _GEN_9497 = 5'h2 == com_idx ? 1'h0 : _GEN_2792; // @[rob.scala 434:{30,30}]
  wire  _GEN_9498 = 5'h3 == com_idx ? 1'h0 : _GEN_2793; // @[rob.scala 434:{30,30}]
  wire  _GEN_9499 = 5'h4 == com_idx ? 1'h0 : _GEN_2794; // @[rob.scala 434:{30,30}]
  wire  _GEN_9500 = 5'h5 == com_idx ? 1'h0 : _GEN_2795; // @[rob.scala 434:{30,30}]
  wire  _GEN_9501 = 5'h6 == com_idx ? 1'h0 : _GEN_2796; // @[rob.scala 434:{30,30}]
  wire  _GEN_9502 = 5'h7 == com_idx ? 1'h0 : _GEN_2797; // @[rob.scala 434:{30,30}]
  wire  _GEN_9503 = 5'h8 == com_idx ? 1'h0 : _GEN_2798; // @[rob.scala 434:{30,30}]
  wire  _GEN_9504 = 5'h9 == com_idx ? 1'h0 : _GEN_2799; // @[rob.scala 434:{30,30}]
  wire  _GEN_9505 = 5'ha == com_idx ? 1'h0 : _GEN_2800; // @[rob.scala 434:{30,30}]
  wire  _GEN_9506 = 5'hb == com_idx ? 1'h0 : _GEN_2801; // @[rob.scala 434:{30,30}]
  wire  _GEN_9507 = 5'hc == com_idx ? 1'h0 : _GEN_2802; // @[rob.scala 434:{30,30}]
  wire  _GEN_9508 = 5'hd == com_idx ? 1'h0 : _GEN_2803; // @[rob.scala 434:{30,30}]
  wire  _GEN_9509 = 5'he == com_idx ? 1'h0 : _GEN_2804; // @[rob.scala 434:{30,30}]
  wire  _GEN_9510 = 5'hf == com_idx ? 1'h0 : _GEN_2805; // @[rob.scala 434:{30,30}]
  wire  _GEN_9511 = 5'h10 == com_idx ? 1'h0 : _GEN_2806; // @[rob.scala 434:{30,30}]
  wire  _GEN_9512 = 5'h11 == com_idx ? 1'h0 : _GEN_2807; // @[rob.scala 434:{30,30}]
  wire  _GEN_9513 = 5'h12 == com_idx ? 1'h0 : _GEN_2808; // @[rob.scala 434:{30,30}]
  wire  _GEN_9514 = 5'h13 == com_idx ? 1'h0 : _GEN_2809; // @[rob.scala 434:{30,30}]
  wire  _GEN_9515 = 5'h14 == com_idx ? 1'h0 : _GEN_2810; // @[rob.scala 434:{30,30}]
  wire  _GEN_9516 = 5'h15 == com_idx ? 1'h0 : _GEN_2811; // @[rob.scala 434:{30,30}]
  wire  _GEN_9517 = 5'h16 == com_idx ? 1'h0 : _GEN_2812; // @[rob.scala 434:{30,30}]
  wire  _GEN_9518 = 5'h17 == com_idx ? 1'h0 : _GEN_2813; // @[rob.scala 434:{30,30}]
  wire  _GEN_9519 = 5'h18 == com_idx ? 1'h0 : _GEN_2814; // @[rob.scala 434:{30,30}]
  wire  _GEN_9520 = 5'h19 == com_idx ? 1'h0 : _GEN_2815; // @[rob.scala 434:{30,30}]
  wire  _GEN_9521 = 5'h1a == com_idx ? 1'h0 : _GEN_2816; // @[rob.scala 434:{30,30}]
  wire  _GEN_9522 = 5'h1b == com_idx ? 1'h0 : _GEN_2817; // @[rob.scala 434:{30,30}]
  wire  _GEN_9523 = 5'h1c == com_idx ? 1'h0 : _GEN_2818; // @[rob.scala 434:{30,30}]
  wire  _GEN_9524 = 5'h1d == com_idx ? 1'h0 : _GEN_2819; // @[rob.scala 434:{30,30}]
  wire  _GEN_9525 = 5'h1e == com_idx ? 1'h0 : _GEN_2820; // @[rob.scala 434:{30,30}]
  wire  _GEN_9526 = 5'h1f == com_idx ? 1'h0 : _GEN_2821; // @[rob.scala 434:{30,30}]
  wire  _GEN_9559 = rbk_row ? _GEN_9495 : _GEN_2790; // @[rob.scala 433:20]
  wire  _GEN_9560 = rbk_row ? _GEN_9496 : _GEN_2791; // @[rob.scala 433:20]
  wire  _GEN_9561 = rbk_row ? _GEN_9497 : _GEN_2792; // @[rob.scala 433:20]
  wire  _GEN_9562 = rbk_row ? _GEN_9498 : _GEN_2793; // @[rob.scala 433:20]
  wire  _GEN_9563 = rbk_row ? _GEN_9499 : _GEN_2794; // @[rob.scala 433:20]
  wire  _GEN_9564 = rbk_row ? _GEN_9500 : _GEN_2795; // @[rob.scala 433:20]
  wire  _GEN_9565 = rbk_row ? _GEN_9501 : _GEN_2796; // @[rob.scala 433:20]
  wire  _GEN_9566 = rbk_row ? _GEN_9502 : _GEN_2797; // @[rob.scala 433:20]
  wire  _GEN_9567 = rbk_row ? _GEN_9503 : _GEN_2798; // @[rob.scala 433:20]
  wire  _GEN_9568 = rbk_row ? _GEN_9504 : _GEN_2799; // @[rob.scala 433:20]
  wire  _GEN_9569 = rbk_row ? _GEN_9505 : _GEN_2800; // @[rob.scala 433:20]
  wire  _GEN_9570 = rbk_row ? _GEN_9506 : _GEN_2801; // @[rob.scala 433:20]
  wire  _GEN_9571 = rbk_row ? _GEN_9507 : _GEN_2802; // @[rob.scala 433:20]
  wire  _GEN_9572 = rbk_row ? _GEN_9508 : _GEN_2803; // @[rob.scala 433:20]
  wire  _GEN_9573 = rbk_row ? _GEN_9509 : _GEN_2804; // @[rob.scala 433:20]
  wire  _GEN_9574 = rbk_row ? _GEN_9510 : _GEN_2805; // @[rob.scala 433:20]
  wire  _GEN_9575 = rbk_row ? _GEN_9511 : _GEN_2806; // @[rob.scala 433:20]
  wire  _GEN_9576 = rbk_row ? _GEN_9512 : _GEN_2807; // @[rob.scala 433:20]
  wire  _GEN_9577 = rbk_row ? _GEN_9513 : _GEN_2808; // @[rob.scala 433:20]
  wire  _GEN_9578 = rbk_row ? _GEN_9514 : _GEN_2809; // @[rob.scala 433:20]
  wire  _GEN_9579 = rbk_row ? _GEN_9515 : _GEN_2810; // @[rob.scala 433:20]
  wire  _GEN_9580 = rbk_row ? _GEN_9516 : _GEN_2811; // @[rob.scala 433:20]
  wire  _GEN_9581 = rbk_row ? _GEN_9517 : _GEN_2812; // @[rob.scala 433:20]
  wire  _GEN_9582 = rbk_row ? _GEN_9518 : _GEN_2813; // @[rob.scala 433:20]
  wire  _GEN_9583 = rbk_row ? _GEN_9519 : _GEN_2814; // @[rob.scala 433:20]
  wire  _GEN_9584 = rbk_row ? _GEN_9520 : _GEN_2815; // @[rob.scala 433:20]
  wire  _GEN_9585 = rbk_row ? _GEN_9521 : _GEN_2816; // @[rob.scala 433:20]
  wire  _GEN_9586 = rbk_row ? _GEN_9522 : _GEN_2817; // @[rob.scala 433:20]
  wire  _GEN_9587 = rbk_row ? _GEN_9523 : _GEN_2818; // @[rob.scala 433:20]
  wire  _GEN_9588 = rbk_row ? _GEN_9524 : _GEN_2819; // @[rob.scala 433:20]
  wire  _GEN_9589 = rbk_row ? _GEN_9525 : _GEN_2820; // @[rob.scala 433:20]
  wire  _GEN_9590 = rbk_row ? _GEN_9526 : _GEN_2821; // @[rob.scala 433:20]
  wire [7:0] _T_91 = io_brupdate_b1_mispredict_mask & rob_uop_0_br_mask; // @[util.scala 118:51]
  wire  _T_92 = _T_91 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_93 = ~io_brupdate_b1_resolve_mask; // @[util.scala 89:23]
  wire [7:0] _T_94 = rob_uop_0_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9624 = _T_92 ? 1'h0 : _GEN_9559; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9625 = _T_92 ? 32'h4033 : _GEN_5318; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_95 = io_brupdate_b1_mispredict_mask & rob_uop_1_br_mask; // @[util.scala 118:51]
  wire  _T_96 = _T_95 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_98 = rob_uop_1_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9628 = _T_96 ? 1'h0 : _GEN_9560; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9629 = _T_96 ? 32'h4033 : _GEN_5319; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_99 = io_brupdate_b1_mispredict_mask & rob_uop_2_br_mask; // @[util.scala 118:51]
  wire  _T_100 = _T_99 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_102 = rob_uop_2_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9632 = _T_100 ? 1'h0 : _GEN_9561; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9633 = _T_100 ? 32'h4033 : _GEN_5320; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_103 = io_brupdate_b1_mispredict_mask & rob_uop_3_br_mask; // @[util.scala 118:51]
  wire  _T_104 = _T_103 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_106 = rob_uop_3_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9636 = _T_104 ? 1'h0 : _GEN_9562; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9637 = _T_104 ? 32'h4033 : _GEN_5321; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_107 = io_brupdate_b1_mispredict_mask & rob_uop_4_br_mask; // @[util.scala 118:51]
  wire  _T_108 = _T_107 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_110 = rob_uop_4_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9640 = _T_108 ? 1'h0 : _GEN_9563; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9641 = _T_108 ? 32'h4033 : _GEN_5322; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_111 = io_brupdate_b1_mispredict_mask & rob_uop_5_br_mask; // @[util.scala 118:51]
  wire  _T_112 = _T_111 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_114 = rob_uop_5_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9644 = _T_112 ? 1'h0 : _GEN_9564; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9645 = _T_112 ? 32'h4033 : _GEN_5323; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_115 = io_brupdate_b1_mispredict_mask & rob_uop_6_br_mask; // @[util.scala 118:51]
  wire  _T_116 = _T_115 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_118 = rob_uop_6_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9648 = _T_116 ? 1'h0 : _GEN_9565; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9649 = _T_116 ? 32'h4033 : _GEN_5324; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_119 = io_brupdate_b1_mispredict_mask & rob_uop_7_br_mask; // @[util.scala 118:51]
  wire  _T_120 = _T_119 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_122 = rob_uop_7_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9652 = _T_120 ? 1'h0 : _GEN_9566; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9653 = _T_120 ? 32'h4033 : _GEN_5325; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_123 = io_brupdate_b1_mispredict_mask & rob_uop_8_br_mask; // @[util.scala 118:51]
  wire  _T_124 = _T_123 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_126 = rob_uop_8_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9656 = _T_124 ? 1'h0 : _GEN_9567; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9657 = _T_124 ? 32'h4033 : _GEN_5326; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_127 = io_brupdate_b1_mispredict_mask & rob_uop_9_br_mask; // @[util.scala 118:51]
  wire  _T_128 = _T_127 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_130 = rob_uop_9_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9660 = _T_128 ? 1'h0 : _GEN_9568; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9661 = _T_128 ? 32'h4033 : _GEN_5327; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_131 = io_brupdate_b1_mispredict_mask & rob_uop_10_br_mask; // @[util.scala 118:51]
  wire  _T_132 = _T_131 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_134 = rob_uop_10_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9664 = _T_132 ? 1'h0 : _GEN_9569; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9665 = _T_132 ? 32'h4033 : _GEN_5328; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_135 = io_brupdate_b1_mispredict_mask & rob_uop_11_br_mask; // @[util.scala 118:51]
  wire  _T_136 = _T_135 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_138 = rob_uop_11_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9668 = _T_136 ? 1'h0 : _GEN_9570; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9669 = _T_136 ? 32'h4033 : _GEN_5329; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_139 = io_brupdate_b1_mispredict_mask & rob_uop_12_br_mask; // @[util.scala 118:51]
  wire  _T_140 = _T_139 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_142 = rob_uop_12_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9672 = _T_140 ? 1'h0 : _GEN_9571; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9673 = _T_140 ? 32'h4033 : _GEN_5330; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_143 = io_brupdate_b1_mispredict_mask & rob_uop_13_br_mask; // @[util.scala 118:51]
  wire  _T_144 = _T_143 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_146 = rob_uop_13_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9676 = _T_144 ? 1'h0 : _GEN_9572; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9677 = _T_144 ? 32'h4033 : _GEN_5331; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_147 = io_brupdate_b1_mispredict_mask & rob_uop_14_br_mask; // @[util.scala 118:51]
  wire  _T_148 = _T_147 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_150 = rob_uop_14_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9680 = _T_148 ? 1'h0 : _GEN_9573; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9681 = _T_148 ? 32'h4033 : _GEN_5332; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_151 = io_brupdate_b1_mispredict_mask & rob_uop_15_br_mask; // @[util.scala 118:51]
  wire  _T_152 = _T_151 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_154 = rob_uop_15_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9684 = _T_152 ? 1'h0 : _GEN_9574; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9685 = _T_152 ? 32'h4033 : _GEN_5333; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_155 = io_brupdate_b1_mispredict_mask & rob_uop_16_br_mask; // @[util.scala 118:51]
  wire  _T_156 = _T_155 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_158 = rob_uop_16_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9688 = _T_156 ? 1'h0 : _GEN_9575; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9689 = _T_156 ? 32'h4033 : _GEN_5334; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_159 = io_brupdate_b1_mispredict_mask & rob_uop_17_br_mask; // @[util.scala 118:51]
  wire  _T_160 = _T_159 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_162 = rob_uop_17_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9692 = _T_160 ? 1'h0 : _GEN_9576; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9693 = _T_160 ? 32'h4033 : _GEN_5335; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_163 = io_brupdate_b1_mispredict_mask & rob_uop_18_br_mask; // @[util.scala 118:51]
  wire  _T_164 = _T_163 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_166 = rob_uop_18_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9696 = _T_164 ? 1'h0 : _GEN_9577; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9697 = _T_164 ? 32'h4033 : _GEN_5336; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_167 = io_brupdate_b1_mispredict_mask & rob_uop_19_br_mask; // @[util.scala 118:51]
  wire  _T_168 = _T_167 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_170 = rob_uop_19_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9700 = _T_168 ? 1'h0 : _GEN_9578; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9701 = _T_168 ? 32'h4033 : _GEN_5337; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_171 = io_brupdate_b1_mispredict_mask & rob_uop_20_br_mask; // @[util.scala 118:51]
  wire  _T_172 = _T_171 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_174 = rob_uop_20_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9704 = _T_172 ? 1'h0 : _GEN_9579; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9705 = _T_172 ? 32'h4033 : _GEN_5338; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_175 = io_brupdate_b1_mispredict_mask & rob_uop_21_br_mask; // @[util.scala 118:51]
  wire  _T_176 = _T_175 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_178 = rob_uop_21_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9708 = _T_176 ? 1'h0 : _GEN_9580; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9709 = _T_176 ? 32'h4033 : _GEN_5339; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_179 = io_brupdate_b1_mispredict_mask & rob_uop_22_br_mask; // @[util.scala 118:51]
  wire  _T_180 = _T_179 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_182 = rob_uop_22_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9712 = _T_180 ? 1'h0 : _GEN_9581; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9713 = _T_180 ? 32'h4033 : _GEN_5340; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_183 = io_brupdate_b1_mispredict_mask & rob_uop_23_br_mask; // @[util.scala 118:51]
  wire  _T_184 = _T_183 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_186 = rob_uop_23_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9716 = _T_184 ? 1'h0 : _GEN_9582; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9717 = _T_184 ? 32'h4033 : _GEN_5341; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_187 = io_brupdate_b1_mispredict_mask & rob_uop_24_br_mask; // @[util.scala 118:51]
  wire  _T_188 = _T_187 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_190 = rob_uop_24_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9720 = _T_188 ? 1'h0 : _GEN_9583; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9721 = _T_188 ? 32'h4033 : _GEN_5342; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_191 = io_brupdate_b1_mispredict_mask & rob_uop_25_br_mask; // @[util.scala 118:51]
  wire  _T_192 = _T_191 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_194 = rob_uop_25_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9724 = _T_192 ? 1'h0 : _GEN_9584; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9725 = _T_192 ? 32'h4033 : _GEN_5343; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_195 = io_brupdate_b1_mispredict_mask & rob_uop_26_br_mask; // @[util.scala 118:51]
  wire  _T_196 = _T_195 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_198 = rob_uop_26_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9728 = _T_196 ? 1'h0 : _GEN_9585; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9729 = _T_196 ? 32'h4033 : _GEN_5344; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_199 = io_brupdate_b1_mispredict_mask & rob_uop_27_br_mask; // @[util.scala 118:51]
  wire  _T_200 = _T_199 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_202 = rob_uop_27_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9732 = _T_200 ? 1'h0 : _GEN_9586; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9733 = _T_200 ? 32'h4033 : _GEN_5345; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_203 = io_brupdate_b1_mispredict_mask & rob_uop_28_br_mask; // @[util.scala 118:51]
  wire  _T_204 = _T_203 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_206 = rob_uop_28_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9736 = _T_204 ? 1'h0 : _GEN_9587; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9737 = _T_204 ? 32'h4033 : _GEN_5346; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_207 = io_brupdate_b1_mispredict_mask & rob_uop_29_br_mask; // @[util.scala 118:51]
  wire  _T_208 = _T_207 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_210 = rob_uop_29_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9740 = _T_208 ? 1'h0 : _GEN_9588; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9741 = _T_208 ? 32'h4033 : _GEN_5347; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_211 = io_brupdate_b1_mispredict_mask & rob_uop_30_br_mask; // @[util.scala 118:51]
  wire  _T_212 = _T_211 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_214 = rob_uop_30_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9744 = _T_212 ? 1'h0 : _GEN_9589; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9745 = _T_212 ? 32'h4033 : _GEN_5348; // @[rob.scala 455:7 457:33]
  wire [7:0] _T_215 = io_brupdate_b1_mispredict_mask & rob_uop_31_br_mask; // @[util.scala 118:51]
  wire  _T_216 = _T_215 != 8'h0; // @[util.scala 118:59]
  wire [7:0] _T_218 = rob_uop_31_br_mask & _T_93; // @[util.scala 89:21]
  wire  _GEN_9748 = _T_216 ? 1'h0 : _GEN_9590; // @[rob.scala 455:7 456:20]
  wire [31:0] _GEN_9749 = _T_216 ? 32'h4033 : _GEN_5349; // @[rob.scala 455:7 457:33]
  wire  _GEN_9976 = 5'h1 == rob_head ? rob_uop_1_uses_ldq : rob_uop_0_uses_ldq; // @[rob.scala 485:{26,26}]
  wire  _GEN_9977 = 5'h2 == rob_head ? rob_uop_2_uses_ldq : _GEN_9976; // @[rob.scala 485:{26,26}]
  wire  _GEN_9978 = 5'h3 == rob_head ? rob_uop_3_uses_ldq : _GEN_9977; // @[rob.scala 485:{26,26}]
  wire  _GEN_9979 = 5'h4 == rob_head ? rob_uop_4_uses_ldq : _GEN_9978; // @[rob.scala 485:{26,26}]
  wire  _GEN_9980 = 5'h5 == rob_head ? rob_uop_5_uses_ldq : _GEN_9979; // @[rob.scala 485:{26,26}]
  wire  _GEN_9981 = 5'h6 == rob_head ? rob_uop_6_uses_ldq : _GEN_9980; // @[rob.scala 485:{26,26}]
  wire  _GEN_9982 = 5'h7 == rob_head ? rob_uop_7_uses_ldq : _GEN_9981; // @[rob.scala 485:{26,26}]
  wire  _GEN_9983 = 5'h8 == rob_head ? rob_uop_8_uses_ldq : _GEN_9982; // @[rob.scala 485:{26,26}]
  wire  _GEN_9984 = 5'h9 == rob_head ? rob_uop_9_uses_ldq : _GEN_9983; // @[rob.scala 485:{26,26}]
  wire  _GEN_9985 = 5'ha == rob_head ? rob_uop_10_uses_ldq : _GEN_9984; // @[rob.scala 485:{26,26}]
  wire  _GEN_9986 = 5'hb == rob_head ? rob_uop_11_uses_ldq : _GEN_9985; // @[rob.scala 485:{26,26}]
  wire  _GEN_9987 = 5'hc == rob_head ? rob_uop_12_uses_ldq : _GEN_9986; // @[rob.scala 485:{26,26}]
  wire  _GEN_9988 = 5'hd == rob_head ? rob_uop_13_uses_ldq : _GEN_9987; // @[rob.scala 485:{26,26}]
  wire  _GEN_9989 = 5'he == rob_head ? rob_uop_14_uses_ldq : _GEN_9988; // @[rob.scala 485:{26,26}]
  wire  _GEN_9990 = 5'hf == rob_head ? rob_uop_15_uses_ldq : _GEN_9989; // @[rob.scala 485:{26,26}]
  wire  _GEN_9991 = 5'h10 == rob_head ? rob_uop_16_uses_ldq : _GEN_9990; // @[rob.scala 485:{26,26}]
  wire  _GEN_9992 = 5'h11 == rob_head ? rob_uop_17_uses_ldq : _GEN_9991; // @[rob.scala 485:{26,26}]
  wire  _GEN_9993 = 5'h12 == rob_head ? rob_uop_18_uses_ldq : _GEN_9992; // @[rob.scala 485:{26,26}]
  wire  _GEN_9994 = 5'h13 == rob_head ? rob_uop_19_uses_ldq : _GEN_9993; // @[rob.scala 485:{26,26}]
  wire  _GEN_9995 = 5'h14 == rob_head ? rob_uop_20_uses_ldq : _GEN_9994; // @[rob.scala 485:{26,26}]
  wire  _GEN_9996 = 5'h15 == rob_head ? rob_uop_21_uses_ldq : _GEN_9995; // @[rob.scala 485:{26,26}]
  wire  _GEN_9997 = 5'h16 == rob_head ? rob_uop_22_uses_ldq : _GEN_9996; // @[rob.scala 485:{26,26}]
  wire  _GEN_9998 = 5'h17 == rob_head ? rob_uop_23_uses_ldq : _GEN_9997; // @[rob.scala 485:{26,26}]
  wire  _GEN_9999 = 5'h18 == rob_head ? rob_uop_24_uses_ldq : _GEN_9998; // @[rob.scala 485:{26,26}]
  wire  _GEN_10000 = 5'h19 == rob_head ? rob_uop_25_uses_ldq : _GEN_9999; // @[rob.scala 485:{26,26}]
  wire  _GEN_10001 = 5'h1a == rob_head ? rob_uop_26_uses_ldq : _GEN_10000; // @[rob.scala 485:{26,26}]
  wire  _GEN_10002 = 5'h1b == rob_head ? rob_uop_27_uses_ldq : _GEN_10001; // @[rob.scala 485:{26,26}]
  wire  _GEN_10003 = 5'h1c == rob_head ? rob_uop_28_uses_ldq : _GEN_10002; // @[rob.scala 485:{26,26}]
  wire  _GEN_10004 = 5'h1d == rob_head ? rob_uop_29_uses_ldq : _GEN_10003; // @[rob.scala 485:{26,26}]
  wire  _GEN_10005 = 5'h1e == rob_head ? rob_uop_30_uses_ldq : _GEN_10004; // @[rob.scala 485:{26,26}]
  wire  rob_head_uses_ldq_0 = 5'h1f == rob_head ? rob_uop_31_uses_ldq : _GEN_10005; // @[rob.scala 485:{26,26}]
  wire  _GEN_10008 = 5'h1 == rob_pnr ? rob_unsafe_1 : rob_unsafe_0; // @[rob.scala 493:{67,67}]
  wire  _GEN_10009 = 5'h2 == rob_pnr ? rob_unsafe_2 : _GEN_10008; // @[rob.scala 493:{67,67}]
  wire  _GEN_10010 = 5'h3 == rob_pnr ? rob_unsafe_3 : _GEN_10009; // @[rob.scala 493:{67,67}]
  wire  _GEN_10011 = 5'h4 == rob_pnr ? rob_unsafe_4 : _GEN_10010; // @[rob.scala 493:{67,67}]
  wire  _GEN_10012 = 5'h5 == rob_pnr ? rob_unsafe_5 : _GEN_10011; // @[rob.scala 493:{67,67}]
  wire  _GEN_10013 = 5'h6 == rob_pnr ? rob_unsafe_6 : _GEN_10012; // @[rob.scala 493:{67,67}]
  wire  _GEN_10014 = 5'h7 == rob_pnr ? rob_unsafe_7 : _GEN_10013; // @[rob.scala 493:{67,67}]
  wire  _GEN_10015 = 5'h8 == rob_pnr ? rob_unsafe_8 : _GEN_10014; // @[rob.scala 493:{67,67}]
  wire  _GEN_10016 = 5'h9 == rob_pnr ? rob_unsafe_9 : _GEN_10015; // @[rob.scala 493:{67,67}]
  wire  _GEN_10017 = 5'ha == rob_pnr ? rob_unsafe_10 : _GEN_10016; // @[rob.scala 493:{67,67}]
  wire  _GEN_10018 = 5'hb == rob_pnr ? rob_unsafe_11 : _GEN_10017; // @[rob.scala 493:{67,67}]
  wire  _GEN_10019 = 5'hc == rob_pnr ? rob_unsafe_12 : _GEN_10018; // @[rob.scala 493:{67,67}]
  wire  _GEN_10020 = 5'hd == rob_pnr ? rob_unsafe_13 : _GEN_10019; // @[rob.scala 493:{67,67}]
  wire  _GEN_10021 = 5'he == rob_pnr ? rob_unsafe_14 : _GEN_10020; // @[rob.scala 493:{67,67}]
  wire  _GEN_10022 = 5'hf == rob_pnr ? rob_unsafe_15 : _GEN_10021; // @[rob.scala 493:{67,67}]
  wire  _GEN_10023 = 5'h10 == rob_pnr ? rob_unsafe_16 : _GEN_10022; // @[rob.scala 493:{67,67}]
  wire  _GEN_10024 = 5'h11 == rob_pnr ? rob_unsafe_17 : _GEN_10023; // @[rob.scala 493:{67,67}]
  wire  _GEN_10025 = 5'h12 == rob_pnr ? rob_unsafe_18 : _GEN_10024; // @[rob.scala 493:{67,67}]
  wire  _GEN_10026 = 5'h13 == rob_pnr ? rob_unsafe_19 : _GEN_10025; // @[rob.scala 493:{67,67}]
  wire  _GEN_10027 = 5'h14 == rob_pnr ? rob_unsafe_20 : _GEN_10026; // @[rob.scala 493:{67,67}]
  wire  _GEN_10028 = 5'h15 == rob_pnr ? rob_unsafe_21 : _GEN_10027; // @[rob.scala 493:{67,67}]
  wire  _GEN_10029 = 5'h16 == rob_pnr ? rob_unsafe_22 : _GEN_10028; // @[rob.scala 493:{67,67}]
  wire  _GEN_10030 = 5'h17 == rob_pnr ? rob_unsafe_23 : _GEN_10029; // @[rob.scala 493:{67,67}]
  wire  _GEN_10031 = 5'h18 == rob_pnr ? rob_unsafe_24 : _GEN_10030; // @[rob.scala 493:{67,67}]
  wire  _GEN_10032 = 5'h19 == rob_pnr ? rob_unsafe_25 : _GEN_10031; // @[rob.scala 493:{67,67}]
  wire  _GEN_10033 = 5'h1a == rob_pnr ? rob_unsafe_26 : _GEN_10032; // @[rob.scala 493:{67,67}]
  wire  _GEN_10034 = 5'h1b == rob_pnr ? rob_unsafe_27 : _GEN_10033; // @[rob.scala 493:{67,67}]
  wire  _GEN_10035 = 5'h1c == rob_pnr ? rob_unsafe_28 : _GEN_10034; // @[rob.scala 493:{67,67}]
  wire  _GEN_10036 = 5'h1d == rob_pnr ? rob_unsafe_29 : _GEN_10035; // @[rob.scala 493:{67,67}]
  wire  _GEN_10037 = 5'h1e == rob_pnr ? rob_unsafe_30 : _GEN_10036; // @[rob.scala 493:{67,67}]
  wire  _GEN_10038 = 5'h1f == rob_pnr ? rob_unsafe_31 : _GEN_10037; // @[rob.scala 493:{67,67}]
  wire  _GEN_10040 = 5'h1 == rob_pnr ? rob_exception_1 : rob_exception_0; // @[rob.scala 493:{67,67}]
  wire  _GEN_10041 = 5'h2 == rob_pnr ? rob_exception_2 : _GEN_10040; // @[rob.scala 493:{67,67}]
  wire  _GEN_10042 = 5'h3 == rob_pnr ? rob_exception_3 : _GEN_10041; // @[rob.scala 493:{67,67}]
  wire  _GEN_10043 = 5'h4 == rob_pnr ? rob_exception_4 : _GEN_10042; // @[rob.scala 493:{67,67}]
  wire  _GEN_10044 = 5'h5 == rob_pnr ? rob_exception_5 : _GEN_10043; // @[rob.scala 493:{67,67}]
  wire  _GEN_10045 = 5'h6 == rob_pnr ? rob_exception_6 : _GEN_10044; // @[rob.scala 493:{67,67}]
  wire  _GEN_10046 = 5'h7 == rob_pnr ? rob_exception_7 : _GEN_10045; // @[rob.scala 493:{67,67}]
  wire  _GEN_10047 = 5'h8 == rob_pnr ? rob_exception_8 : _GEN_10046; // @[rob.scala 493:{67,67}]
  wire  _GEN_10048 = 5'h9 == rob_pnr ? rob_exception_9 : _GEN_10047; // @[rob.scala 493:{67,67}]
  wire  _GEN_10049 = 5'ha == rob_pnr ? rob_exception_10 : _GEN_10048; // @[rob.scala 493:{67,67}]
  wire  _GEN_10050 = 5'hb == rob_pnr ? rob_exception_11 : _GEN_10049; // @[rob.scala 493:{67,67}]
  wire  _GEN_10051 = 5'hc == rob_pnr ? rob_exception_12 : _GEN_10050; // @[rob.scala 493:{67,67}]
  wire  _GEN_10052 = 5'hd == rob_pnr ? rob_exception_13 : _GEN_10051; // @[rob.scala 493:{67,67}]
  wire  _GEN_10053 = 5'he == rob_pnr ? rob_exception_14 : _GEN_10052; // @[rob.scala 493:{67,67}]
  wire  _GEN_10054 = 5'hf == rob_pnr ? rob_exception_15 : _GEN_10053; // @[rob.scala 493:{67,67}]
  wire  _GEN_10055 = 5'h10 == rob_pnr ? rob_exception_16 : _GEN_10054; // @[rob.scala 493:{67,67}]
  wire  _GEN_10056 = 5'h11 == rob_pnr ? rob_exception_17 : _GEN_10055; // @[rob.scala 493:{67,67}]
  wire  _GEN_10057 = 5'h12 == rob_pnr ? rob_exception_18 : _GEN_10056; // @[rob.scala 493:{67,67}]
  wire  _GEN_10058 = 5'h13 == rob_pnr ? rob_exception_19 : _GEN_10057; // @[rob.scala 493:{67,67}]
  wire  _GEN_10059 = 5'h14 == rob_pnr ? rob_exception_20 : _GEN_10058; // @[rob.scala 493:{67,67}]
  wire  _GEN_10060 = 5'h15 == rob_pnr ? rob_exception_21 : _GEN_10059; // @[rob.scala 493:{67,67}]
  wire  _GEN_10061 = 5'h16 == rob_pnr ? rob_exception_22 : _GEN_10060; // @[rob.scala 493:{67,67}]
  wire  _GEN_10062 = 5'h17 == rob_pnr ? rob_exception_23 : _GEN_10061; // @[rob.scala 493:{67,67}]
  wire  _GEN_10063 = 5'h18 == rob_pnr ? rob_exception_24 : _GEN_10062; // @[rob.scala 493:{67,67}]
  wire  _GEN_10064 = 5'h19 == rob_pnr ? rob_exception_25 : _GEN_10063; // @[rob.scala 493:{67,67}]
  wire  _GEN_10065 = 5'h1a == rob_pnr ? rob_exception_26 : _GEN_10064; // @[rob.scala 493:{67,67}]
  wire  _GEN_10066 = 5'h1b == rob_pnr ? rob_exception_27 : _GEN_10065; // @[rob.scala 493:{67,67}]
  wire  _GEN_10067 = 5'h1c == rob_pnr ? rob_exception_28 : _GEN_10066; // @[rob.scala 493:{67,67}]
  wire  _GEN_10068 = 5'h1d == rob_pnr ? rob_exception_29 : _GEN_10067; // @[rob.scala 493:{67,67}]
  wire  _GEN_10069 = 5'h1e == rob_pnr ? rob_exception_30 : _GEN_10068; // @[rob.scala 493:{67,67}]
  wire  _GEN_10070 = 5'h1f == rob_pnr ? rob_exception_31 : _GEN_10069; // @[rob.scala 493:{67,67}]
  wire  _GEN_10072 = 5'h1 == rob_pnr ? rob_val_1 : rob_val_0; // @[rob.scala 493:{43,43}]
  wire  _GEN_10073 = 5'h2 == rob_pnr ? rob_val_2 : _GEN_10072; // @[rob.scala 493:{43,43}]
  wire  _GEN_10074 = 5'h3 == rob_pnr ? rob_val_3 : _GEN_10073; // @[rob.scala 493:{43,43}]
  wire  _GEN_10075 = 5'h4 == rob_pnr ? rob_val_4 : _GEN_10074; // @[rob.scala 493:{43,43}]
  wire  _GEN_10076 = 5'h5 == rob_pnr ? rob_val_5 : _GEN_10075; // @[rob.scala 493:{43,43}]
  wire  _GEN_10077 = 5'h6 == rob_pnr ? rob_val_6 : _GEN_10076; // @[rob.scala 493:{43,43}]
  wire  _GEN_10078 = 5'h7 == rob_pnr ? rob_val_7 : _GEN_10077; // @[rob.scala 493:{43,43}]
  wire  _GEN_10079 = 5'h8 == rob_pnr ? rob_val_8 : _GEN_10078; // @[rob.scala 493:{43,43}]
  wire  _GEN_10080 = 5'h9 == rob_pnr ? rob_val_9 : _GEN_10079; // @[rob.scala 493:{43,43}]
  wire  _GEN_10081 = 5'ha == rob_pnr ? rob_val_10 : _GEN_10080; // @[rob.scala 493:{43,43}]
  wire  _GEN_10082 = 5'hb == rob_pnr ? rob_val_11 : _GEN_10081; // @[rob.scala 493:{43,43}]
  wire  _GEN_10083 = 5'hc == rob_pnr ? rob_val_12 : _GEN_10082; // @[rob.scala 493:{43,43}]
  wire  _GEN_10084 = 5'hd == rob_pnr ? rob_val_13 : _GEN_10083; // @[rob.scala 493:{43,43}]
  wire  _GEN_10085 = 5'he == rob_pnr ? rob_val_14 : _GEN_10084; // @[rob.scala 493:{43,43}]
  wire  _GEN_10086 = 5'hf == rob_pnr ? rob_val_15 : _GEN_10085; // @[rob.scala 493:{43,43}]
  wire  _GEN_10087 = 5'h10 == rob_pnr ? rob_val_16 : _GEN_10086; // @[rob.scala 493:{43,43}]
  wire  _GEN_10088 = 5'h11 == rob_pnr ? rob_val_17 : _GEN_10087; // @[rob.scala 493:{43,43}]
  wire  _GEN_10089 = 5'h12 == rob_pnr ? rob_val_18 : _GEN_10088; // @[rob.scala 493:{43,43}]
  wire  _GEN_10090 = 5'h13 == rob_pnr ? rob_val_19 : _GEN_10089; // @[rob.scala 493:{43,43}]
  wire  _GEN_10091 = 5'h14 == rob_pnr ? rob_val_20 : _GEN_10090; // @[rob.scala 493:{43,43}]
  wire  _GEN_10092 = 5'h15 == rob_pnr ? rob_val_21 : _GEN_10091; // @[rob.scala 493:{43,43}]
  wire  _GEN_10093 = 5'h16 == rob_pnr ? rob_val_22 : _GEN_10092; // @[rob.scala 493:{43,43}]
  wire  _GEN_10094 = 5'h17 == rob_pnr ? rob_val_23 : _GEN_10093; // @[rob.scala 493:{43,43}]
  wire  _GEN_10095 = 5'h18 == rob_pnr ? rob_val_24 : _GEN_10094; // @[rob.scala 493:{43,43}]
  wire  _GEN_10096 = 5'h19 == rob_pnr ? rob_val_25 : _GEN_10095; // @[rob.scala 493:{43,43}]
  wire  _GEN_10097 = 5'h1a == rob_pnr ? rob_val_26 : _GEN_10096; // @[rob.scala 493:{43,43}]
  wire  _GEN_10098 = 5'h1b == rob_pnr ? rob_val_27 : _GEN_10097; // @[rob.scala 493:{43,43}]
  wire  _GEN_10099 = 5'h1c == rob_pnr ? rob_val_28 : _GEN_10098; // @[rob.scala 493:{43,43}]
  wire  _GEN_10100 = 5'h1d == rob_pnr ? rob_val_29 : _GEN_10099; // @[rob.scala 493:{43,43}]
  wire  _GEN_10101 = 5'h1e == rob_pnr ? rob_val_30 : _GEN_10100; // @[rob.scala 493:{43,43}]
  wire  _GEN_10102 = 5'h1f == rob_pnr ? rob_val_31 : _GEN_10101; // @[rob.scala 493:{43,43}]
  wire  rob_pnr_unsafe_0 = _GEN_10102 & (_GEN_10038 | _GEN_10070); // @[rob.scala 493:43]
  wire  _GEN_10237 = 5'h1 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_1 : rob_val_0; // @[rob.scala 515:{16,16}]
  wire  _GEN_10238 = 5'h2 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_2 : _GEN_10237; // @[rob.scala 515:{16,16}]
  wire  _GEN_10239 = 5'h3 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_3 : _GEN_10238; // @[rob.scala 515:{16,16}]
  wire  _GEN_10240 = 5'h4 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_4 : _GEN_10239; // @[rob.scala 515:{16,16}]
  wire  _GEN_10241 = 5'h5 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_5 : _GEN_10240; // @[rob.scala 515:{16,16}]
  wire  _GEN_10242 = 5'h6 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_6 : _GEN_10241; // @[rob.scala 515:{16,16}]
  wire  _GEN_10243 = 5'h7 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_7 : _GEN_10242; // @[rob.scala 515:{16,16}]
  wire  _GEN_10244 = 5'h8 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_8 : _GEN_10243; // @[rob.scala 515:{16,16}]
  wire  _GEN_10245 = 5'h9 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_9 : _GEN_10244; // @[rob.scala 515:{16,16}]
  wire  _GEN_10246 = 5'ha == io_wb_resps_0_bits_uop_rob_idx ? rob_val_10 : _GEN_10245; // @[rob.scala 515:{16,16}]
  wire  _GEN_10247 = 5'hb == io_wb_resps_0_bits_uop_rob_idx ? rob_val_11 : _GEN_10246; // @[rob.scala 515:{16,16}]
  wire  _GEN_10248 = 5'hc == io_wb_resps_0_bits_uop_rob_idx ? rob_val_12 : _GEN_10247; // @[rob.scala 515:{16,16}]
  wire  _GEN_10249 = 5'hd == io_wb_resps_0_bits_uop_rob_idx ? rob_val_13 : _GEN_10248; // @[rob.scala 515:{16,16}]
  wire  _GEN_10250 = 5'he == io_wb_resps_0_bits_uop_rob_idx ? rob_val_14 : _GEN_10249; // @[rob.scala 515:{16,16}]
  wire  _GEN_10251 = 5'hf == io_wb_resps_0_bits_uop_rob_idx ? rob_val_15 : _GEN_10250; // @[rob.scala 515:{16,16}]
  wire  _GEN_10252 = 5'h10 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_16 : _GEN_10251; // @[rob.scala 515:{16,16}]
  wire  _GEN_10253 = 5'h11 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_17 : _GEN_10252; // @[rob.scala 515:{16,16}]
  wire  _GEN_10254 = 5'h12 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_18 : _GEN_10253; // @[rob.scala 515:{16,16}]
  wire  _GEN_10255 = 5'h13 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_19 : _GEN_10254; // @[rob.scala 515:{16,16}]
  wire  _GEN_10256 = 5'h14 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_20 : _GEN_10255; // @[rob.scala 515:{16,16}]
  wire  _GEN_10257 = 5'h15 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_21 : _GEN_10256; // @[rob.scala 515:{16,16}]
  wire  _GEN_10258 = 5'h16 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_22 : _GEN_10257; // @[rob.scala 515:{16,16}]
  wire  _GEN_10259 = 5'h17 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_23 : _GEN_10258; // @[rob.scala 515:{16,16}]
  wire  _GEN_10260 = 5'h18 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_24 : _GEN_10259; // @[rob.scala 515:{16,16}]
  wire  _GEN_10261 = 5'h19 == io_wb_resps_0_bits_uop_rob_idx ? rob_val_25 : _GEN_10260; // @[rob.scala 515:{16,16}]
  wire  _GEN_10262 = 5'h1a == io_wb_resps_0_bits_uop_rob_idx ? rob_val_26 : _GEN_10261; // @[rob.scala 515:{16,16}]
  wire  _GEN_10263 = 5'h1b == io_wb_resps_0_bits_uop_rob_idx ? rob_val_27 : _GEN_10262; // @[rob.scala 515:{16,16}]
  wire  _GEN_10264 = 5'h1c == io_wb_resps_0_bits_uop_rob_idx ? rob_val_28 : _GEN_10263; // @[rob.scala 515:{16,16}]
  wire  _GEN_10265 = 5'h1d == io_wb_resps_0_bits_uop_rob_idx ? rob_val_29 : _GEN_10264; // @[rob.scala 515:{16,16}]
  wire  _GEN_10266 = 5'h1e == io_wb_resps_0_bits_uop_rob_idx ? rob_val_30 : _GEN_10265; // @[rob.scala 515:{16,16}]
  wire  _GEN_10267 = 5'h1f == io_wb_resps_0_bits_uop_rob_idx ? rob_val_31 : _GEN_10266; // @[rob.scala 515:{16,16}]
  wire  _T_293 = ~_GEN_10267; // @[rob.scala 515:16]
  wire  _GEN_10269 = 5'h1 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_1 : rob_bsy_0; // @[rob.scala 518:{16,16}]
  wire  _GEN_10270 = 5'h2 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_2 : _GEN_10269; // @[rob.scala 518:{16,16}]
  wire  _GEN_10271 = 5'h3 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_3 : _GEN_10270; // @[rob.scala 518:{16,16}]
  wire  _GEN_10272 = 5'h4 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_4 : _GEN_10271; // @[rob.scala 518:{16,16}]
  wire  _GEN_10273 = 5'h5 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_5 : _GEN_10272; // @[rob.scala 518:{16,16}]
  wire  _GEN_10274 = 5'h6 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_6 : _GEN_10273; // @[rob.scala 518:{16,16}]
  wire  _GEN_10275 = 5'h7 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_7 : _GEN_10274; // @[rob.scala 518:{16,16}]
  wire  _GEN_10276 = 5'h8 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_8 : _GEN_10275; // @[rob.scala 518:{16,16}]
  wire  _GEN_10277 = 5'h9 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_9 : _GEN_10276; // @[rob.scala 518:{16,16}]
  wire  _GEN_10278 = 5'ha == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_10 : _GEN_10277; // @[rob.scala 518:{16,16}]
  wire  _GEN_10279 = 5'hb == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_11 : _GEN_10278; // @[rob.scala 518:{16,16}]
  wire  _GEN_10280 = 5'hc == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_12 : _GEN_10279; // @[rob.scala 518:{16,16}]
  wire  _GEN_10281 = 5'hd == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_13 : _GEN_10280; // @[rob.scala 518:{16,16}]
  wire  _GEN_10282 = 5'he == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_14 : _GEN_10281; // @[rob.scala 518:{16,16}]
  wire  _GEN_10283 = 5'hf == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_15 : _GEN_10282; // @[rob.scala 518:{16,16}]
  wire  _GEN_10284 = 5'h10 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_16 : _GEN_10283; // @[rob.scala 518:{16,16}]
  wire  _GEN_10285 = 5'h11 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_17 : _GEN_10284; // @[rob.scala 518:{16,16}]
  wire  _GEN_10286 = 5'h12 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_18 : _GEN_10285; // @[rob.scala 518:{16,16}]
  wire  _GEN_10287 = 5'h13 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_19 : _GEN_10286; // @[rob.scala 518:{16,16}]
  wire  _GEN_10288 = 5'h14 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_20 : _GEN_10287; // @[rob.scala 518:{16,16}]
  wire  _GEN_10289 = 5'h15 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_21 : _GEN_10288; // @[rob.scala 518:{16,16}]
  wire  _GEN_10290 = 5'h16 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_22 : _GEN_10289; // @[rob.scala 518:{16,16}]
  wire  _GEN_10291 = 5'h17 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_23 : _GEN_10290; // @[rob.scala 518:{16,16}]
  wire  _GEN_10292 = 5'h18 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_24 : _GEN_10291; // @[rob.scala 518:{16,16}]
  wire  _GEN_10293 = 5'h19 == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_25 : _GEN_10292; // @[rob.scala 518:{16,16}]
  wire  _GEN_10294 = 5'h1a == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_26 : _GEN_10293; // @[rob.scala 518:{16,16}]
  wire  _GEN_10295 = 5'h1b == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_27 : _GEN_10294; // @[rob.scala 518:{16,16}]
  wire  _GEN_10296 = 5'h1c == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_28 : _GEN_10295; // @[rob.scala 518:{16,16}]
  wire  _GEN_10297 = 5'h1d == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_29 : _GEN_10296; // @[rob.scala 518:{16,16}]
  wire  _GEN_10298 = 5'h1e == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_30 : _GEN_10297; // @[rob.scala 518:{16,16}]
  wire  _GEN_10299 = 5'h1f == io_wb_resps_0_bits_uop_rob_idx ? rob_bsy_31 : _GEN_10298; // @[rob.scala 518:{16,16}]
  wire  _T_301 = ~_GEN_10299; // @[rob.scala 518:16]
  wire  _GEN_10301 = 5'h1 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_1_ldst_val : rob_uop_0_ldst_val; // @[rob.scala 520:{72,72}]
  wire  _GEN_10302 = 5'h2 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_2_ldst_val : _GEN_10301; // @[rob.scala 520:{72,72}]
  wire  _GEN_10303 = 5'h3 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_3_ldst_val : _GEN_10302; // @[rob.scala 520:{72,72}]
  wire  _GEN_10304 = 5'h4 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_4_ldst_val : _GEN_10303; // @[rob.scala 520:{72,72}]
  wire  _GEN_10305 = 5'h5 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_5_ldst_val : _GEN_10304; // @[rob.scala 520:{72,72}]
  wire  _GEN_10306 = 5'h6 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_6_ldst_val : _GEN_10305; // @[rob.scala 520:{72,72}]
  wire  _GEN_10307 = 5'h7 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_7_ldst_val : _GEN_10306; // @[rob.scala 520:{72,72}]
  wire  _GEN_10308 = 5'h8 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_8_ldst_val : _GEN_10307; // @[rob.scala 520:{72,72}]
  wire  _GEN_10309 = 5'h9 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_9_ldst_val : _GEN_10308; // @[rob.scala 520:{72,72}]
  wire  _GEN_10310 = 5'ha == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_10_ldst_val : _GEN_10309; // @[rob.scala 520:{72,72}]
  wire  _GEN_10311 = 5'hb == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_11_ldst_val : _GEN_10310; // @[rob.scala 520:{72,72}]
  wire  _GEN_10312 = 5'hc == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_12_ldst_val : _GEN_10311; // @[rob.scala 520:{72,72}]
  wire  _GEN_10313 = 5'hd == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_13_ldst_val : _GEN_10312; // @[rob.scala 520:{72,72}]
  wire  _GEN_10314 = 5'he == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_14_ldst_val : _GEN_10313; // @[rob.scala 520:{72,72}]
  wire  _GEN_10315 = 5'hf == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_15_ldst_val : _GEN_10314; // @[rob.scala 520:{72,72}]
  wire  _GEN_10316 = 5'h10 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_16_ldst_val : _GEN_10315; // @[rob.scala 520:{72,72}]
  wire  _GEN_10317 = 5'h11 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_17_ldst_val : _GEN_10316; // @[rob.scala 520:{72,72}]
  wire  _GEN_10318 = 5'h12 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_18_ldst_val : _GEN_10317; // @[rob.scala 520:{72,72}]
  wire  _GEN_10319 = 5'h13 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_19_ldst_val : _GEN_10318; // @[rob.scala 520:{72,72}]
  wire  _GEN_10320 = 5'h14 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_20_ldst_val : _GEN_10319; // @[rob.scala 520:{72,72}]
  wire  _GEN_10321 = 5'h15 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_21_ldst_val : _GEN_10320; // @[rob.scala 520:{72,72}]
  wire  _GEN_10322 = 5'h16 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_22_ldst_val : _GEN_10321; // @[rob.scala 520:{72,72}]
  wire  _GEN_10323 = 5'h17 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_23_ldst_val : _GEN_10322; // @[rob.scala 520:{72,72}]
  wire  _GEN_10324 = 5'h18 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_24_ldst_val : _GEN_10323; // @[rob.scala 520:{72,72}]
  wire  _GEN_10325 = 5'h19 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_25_ldst_val : _GEN_10324; // @[rob.scala 520:{72,72}]
  wire  _GEN_10326 = 5'h1a == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_26_ldst_val : _GEN_10325; // @[rob.scala 520:{72,72}]
  wire  _GEN_10327 = 5'h1b == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_27_ldst_val : _GEN_10326; // @[rob.scala 520:{72,72}]
  wire  _GEN_10328 = 5'h1c == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_28_ldst_val : _GEN_10327; // @[rob.scala 520:{72,72}]
  wire  _GEN_10329 = 5'h1d == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_29_ldst_val : _GEN_10328; // @[rob.scala 520:{72,72}]
  wire  _GEN_10330 = 5'h1e == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_30_ldst_val : _GEN_10329; // @[rob.scala 520:{72,72}]
  wire  _GEN_10331 = 5'h1f == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_31_ldst_val : _GEN_10330; // @[rob.scala 520:{72,72}]
  wire  _T_309 = io_wb_resps_0_valid & _GEN_10331; // @[rob.scala 520:72]
  wire [5:0] _GEN_10333 = 5'h1 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_1_pdst : rob_uop_0_pdst; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10334 = 5'h2 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_2_pdst : _GEN_10333; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10335 = 5'h3 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_3_pdst : _GEN_10334; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10336 = 5'h4 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_4_pdst : _GEN_10335; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10337 = 5'h5 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_5_pdst : _GEN_10336; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10338 = 5'h6 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_6_pdst : _GEN_10337; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10339 = 5'h7 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_7_pdst : _GEN_10338; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10340 = 5'h8 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_8_pdst : _GEN_10339; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10341 = 5'h9 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_9_pdst : _GEN_10340; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10342 = 5'ha == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_10_pdst : _GEN_10341; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10343 = 5'hb == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_11_pdst : _GEN_10342; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10344 = 5'hc == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_12_pdst : _GEN_10343; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10345 = 5'hd == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_13_pdst : _GEN_10344; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10346 = 5'he == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_14_pdst : _GEN_10345; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10347 = 5'hf == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_15_pdst : _GEN_10346; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10348 = 5'h10 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_16_pdst : _GEN_10347; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10349 = 5'h11 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_17_pdst : _GEN_10348; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10350 = 5'h12 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_18_pdst : _GEN_10349; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10351 = 5'h13 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_19_pdst : _GEN_10350; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10352 = 5'h14 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_20_pdst : _GEN_10351; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10353 = 5'h15 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_21_pdst : _GEN_10352; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10354 = 5'h16 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_22_pdst : _GEN_10353; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10355 = 5'h17 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_23_pdst : _GEN_10354; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10356 = 5'h18 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_24_pdst : _GEN_10355; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10357 = 5'h19 == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_25_pdst : _GEN_10356; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10358 = 5'h1a == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_26_pdst : _GEN_10357; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10359 = 5'h1b == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_27_pdst : _GEN_10358; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10360 = 5'h1c == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_28_pdst : _GEN_10359; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10361 = 5'h1d == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_29_pdst : _GEN_10360; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10362 = 5'h1e == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_30_pdst : _GEN_10361; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10363 = 5'h1f == io_wb_resps_0_bits_uop_rob_idx ? rob_uop_31_pdst : _GEN_10362; // @[rob.scala 521:{51,51}]
  wire  _T_311 = _T_309 & _GEN_10363 != io_wb_resps_0_bits_uop_pdst; // @[rob.scala 521:34]
  wire  _GEN_10370 = 5'h1 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_1 : rob_val_0; // @[rob.scala 515:{16,16}]
  wire  _GEN_10371 = 5'h2 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_2 : _GEN_10370; // @[rob.scala 515:{16,16}]
  wire  _GEN_10372 = 5'h3 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_3 : _GEN_10371; // @[rob.scala 515:{16,16}]
  wire  _GEN_10373 = 5'h4 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_4 : _GEN_10372; // @[rob.scala 515:{16,16}]
  wire  _GEN_10374 = 5'h5 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_5 : _GEN_10373; // @[rob.scala 515:{16,16}]
  wire  _GEN_10375 = 5'h6 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_6 : _GEN_10374; // @[rob.scala 515:{16,16}]
  wire  _GEN_10376 = 5'h7 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_7 : _GEN_10375; // @[rob.scala 515:{16,16}]
  wire  _GEN_10377 = 5'h8 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_8 : _GEN_10376; // @[rob.scala 515:{16,16}]
  wire  _GEN_10378 = 5'h9 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_9 : _GEN_10377; // @[rob.scala 515:{16,16}]
  wire  _GEN_10379 = 5'ha == io_wb_resps_1_bits_uop_rob_idx ? rob_val_10 : _GEN_10378; // @[rob.scala 515:{16,16}]
  wire  _GEN_10380 = 5'hb == io_wb_resps_1_bits_uop_rob_idx ? rob_val_11 : _GEN_10379; // @[rob.scala 515:{16,16}]
  wire  _GEN_10381 = 5'hc == io_wb_resps_1_bits_uop_rob_idx ? rob_val_12 : _GEN_10380; // @[rob.scala 515:{16,16}]
  wire  _GEN_10382 = 5'hd == io_wb_resps_1_bits_uop_rob_idx ? rob_val_13 : _GEN_10381; // @[rob.scala 515:{16,16}]
  wire  _GEN_10383 = 5'he == io_wb_resps_1_bits_uop_rob_idx ? rob_val_14 : _GEN_10382; // @[rob.scala 515:{16,16}]
  wire  _GEN_10384 = 5'hf == io_wb_resps_1_bits_uop_rob_idx ? rob_val_15 : _GEN_10383; // @[rob.scala 515:{16,16}]
  wire  _GEN_10385 = 5'h10 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_16 : _GEN_10384; // @[rob.scala 515:{16,16}]
  wire  _GEN_10386 = 5'h11 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_17 : _GEN_10385; // @[rob.scala 515:{16,16}]
  wire  _GEN_10387 = 5'h12 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_18 : _GEN_10386; // @[rob.scala 515:{16,16}]
  wire  _GEN_10388 = 5'h13 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_19 : _GEN_10387; // @[rob.scala 515:{16,16}]
  wire  _GEN_10389 = 5'h14 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_20 : _GEN_10388; // @[rob.scala 515:{16,16}]
  wire  _GEN_10390 = 5'h15 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_21 : _GEN_10389; // @[rob.scala 515:{16,16}]
  wire  _GEN_10391 = 5'h16 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_22 : _GEN_10390; // @[rob.scala 515:{16,16}]
  wire  _GEN_10392 = 5'h17 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_23 : _GEN_10391; // @[rob.scala 515:{16,16}]
  wire  _GEN_10393 = 5'h18 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_24 : _GEN_10392; // @[rob.scala 515:{16,16}]
  wire  _GEN_10394 = 5'h19 == io_wb_resps_1_bits_uop_rob_idx ? rob_val_25 : _GEN_10393; // @[rob.scala 515:{16,16}]
  wire  _GEN_10395 = 5'h1a == io_wb_resps_1_bits_uop_rob_idx ? rob_val_26 : _GEN_10394; // @[rob.scala 515:{16,16}]
  wire  _GEN_10396 = 5'h1b == io_wb_resps_1_bits_uop_rob_idx ? rob_val_27 : _GEN_10395; // @[rob.scala 515:{16,16}]
  wire  _GEN_10397 = 5'h1c == io_wb_resps_1_bits_uop_rob_idx ? rob_val_28 : _GEN_10396; // @[rob.scala 515:{16,16}]
  wire  _GEN_10398 = 5'h1d == io_wb_resps_1_bits_uop_rob_idx ? rob_val_29 : _GEN_10397; // @[rob.scala 515:{16,16}]
  wire  _GEN_10399 = 5'h1e == io_wb_resps_1_bits_uop_rob_idx ? rob_val_30 : _GEN_10398; // @[rob.scala 515:{16,16}]
  wire  _GEN_10400 = 5'h1f == io_wb_resps_1_bits_uop_rob_idx ? rob_val_31 : _GEN_10399; // @[rob.scala 515:{16,16}]
  wire  _T_321 = ~_GEN_10400; // @[rob.scala 515:16]
  wire  _GEN_10402 = 5'h1 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_1 : rob_bsy_0; // @[rob.scala 518:{16,16}]
  wire  _GEN_10403 = 5'h2 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_2 : _GEN_10402; // @[rob.scala 518:{16,16}]
  wire  _GEN_10404 = 5'h3 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_3 : _GEN_10403; // @[rob.scala 518:{16,16}]
  wire  _GEN_10405 = 5'h4 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_4 : _GEN_10404; // @[rob.scala 518:{16,16}]
  wire  _GEN_10406 = 5'h5 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_5 : _GEN_10405; // @[rob.scala 518:{16,16}]
  wire  _GEN_10407 = 5'h6 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_6 : _GEN_10406; // @[rob.scala 518:{16,16}]
  wire  _GEN_10408 = 5'h7 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_7 : _GEN_10407; // @[rob.scala 518:{16,16}]
  wire  _GEN_10409 = 5'h8 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_8 : _GEN_10408; // @[rob.scala 518:{16,16}]
  wire  _GEN_10410 = 5'h9 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_9 : _GEN_10409; // @[rob.scala 518:{16,16}]
  wire  _GEN_10411 = 5'ha == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_10 : _GEN_10410; // @[rob.scala 518:{16,16}]
  wire  _GEN_10412 = 5'hb == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_11 : _GEN_10411; // @[rob.scala 518:{16,16}]
  wire  _GEN_10413 = 5'hc == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_12 : _GEN_10412; // @[rob.scala 518:{16,16}]
  wire  _GEN_10414 = 5'hd == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_13 : _GEN_10413; // @[rob.scala 518:{16,16}]
  wire  _GEN_10415 = 5'he == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_14 : _GEN_10414; // @[rob.scala 518:{16,16}]
  wire  _GEN_10416 = 5'hf == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_15 : _GEN_10415; // @[rob.scala 518:{16,16}]
  wire  _GEN_10417 = 5'h10 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_16 : _GEN_10416; // @[rob.scala 518:{16,16}]
  wire  _GEN_10418 = 5'h11 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_17 : _GEN_10417; // @[rob.scala 518:{16,16}]
  wire  _GEN_10419 = 5'h12 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_18 : _GEN_10418; // @[rob.scala 518:{16,16}]
  wire  _GEN_10420 = 5'h13 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_19 : _GEN_10419; // @[rob.scala 518:{16,16}]
  wire  _GEN_10421 = 5'h14 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_20 : _GEN_10420; // @[rob.scala 518:{16,16}]
  wire  _GEN_10422 = 5'h15 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_21 : _GEN_10421; // @[rob.scala 518:{16,16}]
  wire  _GEN_10423 = 5'h16 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_22 : _GEN_10422; // @[rob.scala 518:{16,16}]
  wire  _GEN_10424 = 5'h17 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_23 : _GEN_10423; // @[rob.scala 518:{16,16}]
  wire  _GEN_10425 = 5'h18 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_24 : _GEN_10424; // @[rob.scala 518:{16,16}]
  wire  _GEN_10426 = 5'h19 == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_25 : _GEN_10425; // @[rob.scala 518:{16,16}]
  wire  _GEN_10427 = 5'h1a == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_26 : _GEN_10426; // @[rob.scala 518:{16,16}]
  wire  _GEN_10428 = 5'h1b == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_27 : _GEN_10427; // @[rob.scala 518:{16,16}]
  wire  _GEN_10429 = 5'h1c == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_28 : _GEN_10428; // @[rob.scala 518:{16,16}]
  wire  _GEN_10430 = 5'h1d == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_29 : _GEN_10429; // @[rob.scala 518:{16,16}]
  wire  _GEN_10431 = 5'h1e == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_30 : _GEN_10430; // @[rob.scala 518:{16,16}]
  wire  _GEN_10432 = 5'h1f == io_wb_resps_1_bits_uop_rob_idx ? rob_bsy_31 : _GEN_10431; // @[rob.scala 518:{16,16}]
  wire  _T_329 = ~_GEN_10432; // @[rob.scala 518:16]
  wire  _GEN_10434 = 5'h1 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_1_ldst_val : rob_uop_0_ldst_val; // @[rob.scala 520:{72,72}]
  wire  _GEN_10435 = 5'h2 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_2_ldst_val : _GEN_10434; // @[rob.scala 520:{72,72}]
  wire  _GEN_10436 = 5'h3 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_3_ldst_val : _GEN_10435; // @[rob.scala 520:{72,72}]
  wire  _GEN_10437 = 5'h4 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_4_ldst_val : _GEN_10436; // @[rob.scala 520:{72,72}]
  wire  _GEN_10438 = 5'h5 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_5_ldst_val : _GEN_10437; // @[rob.scala 520:{72,72}]
  wire  _GEN_10439 = 5'h6 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_6_ldst_val : _GEN_10438; // @[rob.scala 520:{72,72}]
  wire  _GEN_10440 = 5'h7 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_7_ldst_val : _GEN_10439; // @[rob.scala 520:{72,72}]
  wire  _GEN_10441 = 5'h8 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_8_ldst_val : _GEN_10440; // @[rob.scala 520:{72,72}]
  wire  _GEN_10442 = 5'h9 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_9_ldst_val : _GEN_10441; // @[rob.scala 520:{72,72}]
  wire  _GEN_10443 = 5'ha == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_10_ldst_val : _GEN_10442; // @[rob.scala 520:{72,72}]
  wire  _GEN_10444 = 5'hb == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_11_ldst_val : _GEN_10443; // @[rob.scala 520:{72,72}]
  wire  _GEN_10445 = 5'hc == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_12_ldst_val : _GEN_10444; // @[rob.scala 520:{72,72}]
  wire  _GEN_10446 = 5'hd == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_13_ldst_val : _GEN_10445; // @[rob.scala 520:{72,72}]
  wire  _GEN_10447 = 5'he == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_14_ldst_val : _GEN_10446; // @[rob.scala 520:{72,72}]
  wire  _GEN_10448 = 5'hf == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_15_ldst_val : _GEN_10447; // @[rob.scala 520:{72,72}]
  wire  _GEN_10449 = 5'h10 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_16_ldst_val : _GEN_10448; // @[rob.scala 520:{72,72}]
  wire  _GEN_10450 = 5'h11 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_17_ldst_val : _GEN_10449; // @[rob.scala 520:{72,72}]
  wire  _GEN_10451 = 5'h12 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_18_ldst_val : _GEN_10450; // @[rob.scala 520:{72,72}]
  wire  _GEN_10452 = 5'h13 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_19_ldst_val : _GEN_10451; // @[rob.scala 520:{72,72}]
  wire  _GEN_10453 = 5'h14 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_20_ldst_val : _GEN_10452; // @[rob.scala 520:{72,72}]
  wire  _GEN_10454 = 5'h15 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_21_ldst_val : _GEN_10453; // @[rob.scala 520:{72,72}]
  wire  _GEN_10455 = 5'h16 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_22_ldst_val : _GEN_10454; // @[rob.scala 520:{72,72}]
  wire  _GEN_10456 = 5'h17 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_23_ldst_val : _GEN_10455; // @[rob.scala 520:{72,72}]
  wire  _GEN_10457 = 5'h18 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_24_ldst_val : _GEN_10456; // @[rob.scala 520:{72,72}]
  wire  _GEN_10458 = 5'h19 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_25_ldst_val : _GEN_10457; // @[rob.scala 520:{72,72}]
  wire  _GEN_10459 = 5'h1a == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_26_ldst_val : _GEN_10458; // @[rob.scala 520:{72,72}]
  wire  _GEN_10460 = 5'h1b == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_27_ldst_val : _GEN_10459; // @[rob.scala 520:{72,72}]
  wire  _GEN_10461 = 5'h1c == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_28_ldst_val : _GEN_10460; // @[rob.scala 520:{72,72}]
  wire  _GEN_10462 = 5'h1d == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_29_ldst_val : _GEN_10461; // @[rob.scala 520:{72,72}]
  wire  _GEN_10463 = 5'h1e == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_30_ldst_val : _GEN_10462; // @[rob.scala 520:{72,72}]
  wire  _GEN_10464 = 5'h1f == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_31_ldst_val : _GEN_10463; // @[rob.scala 520:{72,72}]
  wire  _T_337 = io_wb_resps_1_valid & _GEN_10464; // @[rob.scala 520:72]
  wire [5:0] _GEN_10466 = 5'h1 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_1_pdst : rob_uop_0_pdst; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10467 = 5'h2 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_2_pdst : _GEN_10466; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10468 = 5'h3 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_3_pdst : _GEN_10467; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10469 = 5'h4 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_4_pdst : _GEN_10468; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10470 = 5'h5 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_5_pdst : _GEN_10469; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10471 = 5'h6 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_6_pdst : _GEN_10470; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10472 = 5'h7 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_7_pdst : _GEN_10471; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10473 = 5'h8 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_8_pdst : _GEN_10472; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10474 = 5'h9 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_9_pdst : _GEN_10473; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10475 = 5'ha == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_10_pdst : _GEN_10474; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10476 = 5'hb == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_11_pdst : _GEN_10475; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10477 = 5'hc == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_12_pdst : _GEN_10476; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10478 = 5'hd == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_13_pdst : _GEN_10477; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10479 = 5'he == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_14_pdst : _GEN_10478; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10480 = 5'hf == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_15_pdst : _GEN_10479; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10481 = 5'h10 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_16_pdst : _GEN_10480; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10482 = 5'h11 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_17_pdst : _GEN_10481; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10483 = 5'h12 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_18_pdst : _GEN_10482; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10484 = 5'h13 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_19_pdst : _GEN_10483; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10485 = 5'h14 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_20_pdst : _GEN_10484; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10486 = 5'h15 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_21_pdst : _GEN_10485; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10487 = 5'h16 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_22_pdst : _GEN_10486; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10488 = 5'h17 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_23_pdst : _GEN_10487; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10489 = 5'h18 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_24_pdst : _GEN_10488; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10490 = 5'h19 == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_25_pdst : _GEN_10489; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10491 = 5'h1a == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_26_pdst : _GEN_10490; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10492 = 5'h1b == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_27_pdst : _GEN_10491; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10493 = 5'h1c == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_28_pdst : _GEN_10492; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10494 = 5'h1d == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_29_pdst : _GEN_10493; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10495 = 5'h1e == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_30_pdst : _GEN_10494; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10496 = 5'h1f == io_wb_resps_1_bits_uop_rob_idx ? rob_uop_31_pdst : _GEN_10495; // @[rob.scala 521:{51,51}]
  wire  _T_339 = _T_337 & _GEN_10496 != io_wb_resps_1_bits_uop_pdst; // @[rob.scala 521:34]
  wire  _GEN_10503 = 5'h1 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_1 : rob_val_0; // @[rob.scala 515:{16,16}]
  wire  _GEN_10504 = 5'h2 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_2 : _GEN_10503; // @[rob.scala 515:{16,16}]
  wire  _GEN_10505 = 5'h3 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_3 : _GEN_10504; // @[rob.scala 515:{16,16}]
  wire  _GEN_10506 = 5'h4 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_4 : _GEN_10505; // @[rob.scala 515:{16,16}]
  wire  _GEN_10507 = 5'h5 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_5 : _GEN_10506; // @[rob.scala 515:{16,16}]
  wire  _GEN_10508 = 5'h6 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_6 : _GEN_10507; // @[rob.scala 515:{16,16}]
  wire  _GEN_10509 = 5'h7 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_7 : _GEN_10508; // @[rob.scala 515:{16,16}]
  wire  _GEN_10510 = 5'h8 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_8 : _GEN_10509; // @[rob.scala 515:{16,16}]
  wire  _GEN_10511 = 5'h9 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_9 : _GEN_10510; // @[rob.scala 515:{16,16}]
  wire  _GEN_10512 = 5'ha == io_wb_resps_2_bits_uop_rob_idx ? rob_val_10 : _GEN_10511; // @[rob.scala 515:{16,16}]
  wire  _GEN_10513 = 5'hb == io_wb_resps_2_bits_uop_rob_idx ? rob_val_11 : _GEN_10512; // @[rob.scala 515:{16,16}]
  wire  _GEN_10514 = 5'hc == io_wb_resps_2_bits_uop_rob_idx ? rob_val_12 : _GEN_10513; // @[rob.scala 515:{16,16}]
  wire  _GEN_10515 = 5'hd == io_wb_resps_2_bits_uop_rob_idx ? rob_val_13 : _GEN_10514; // @[rob.scala 515:{16,16}]
  wire  _GEN_10516 = 5'he == io_wb_resps_2_bits_uop_rob_idx ? rob_val_14 : _GEN_10515; // @[rob.scala 515:{16,16}]
  wire  _GEN_10517 = 5'hf == io_wb_resps_2_bits_uop_rob_idx ? rob_val_15 : _GEN_10516; // @[rob.scala 515:{16,16}]
  wire  _GEN_10518 = 5'h10 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_16 : _GEN_10517; // @[rob.scala 515:{16,16}]
  wire  _GEN_10519 = 5'h11 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_17 : _GEN_10518; // @[rob.scala 515:{16,16}]
  wire  _GEN_10520 = 5'h12 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_18 : _GEN_10519; // @[rob.scala 515:{16,16}]
  wire  _GEN_10521 = 5'h13 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_19 : _GEN_10520; // @[rob.scala 515:{16,16}]
  wire  _GEN_10522 = 5'h14 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_20 : _GEN_10521; // @[rob.scala 515:{16,16}]
  wire  _GEN_10523 = 5'h15 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_21 : _GEN_10522; // @[rob.scala 515:{16,16}]
  wire  _GEN_10524 = 5'h16 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_22 : _GEN_10523; // @[rob.scala 515:{16,16}]
  wire  _GEN_10525 = 5'h17 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_23 : _GEN_10524; // @[rob.scala 515:{16,16}]
  wire  _GEN_10526 = 5'h18 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_24 : _GEN_10525; // @[rob.scala 515:{16,16}]
  wire  _GEN_10527 = 5'h19 == io_wb_resps_2_bits_uop_rob_idx ? rob_val_25 : _GEN_10526; // @[rob.scala 515:{16,16}]
  wire  _GEN_10528 = 5'h1a == io_wb_resps_2_bits_uop_rob_idx ? rob_val_26 : _GEN_10527; // @[rob.scala 515:{16,16}]
  wire  _GEN_10529 = 5'h1b == io_wb_resps_2_bits_uop_rob_idx ? rob_val_27 : _GEN_10528; // @[rob.scala 515:{16,16}]
  wire  _GEN_10530 = 5'h1c == io_wb_resps_2_bits_uop_rob_idx ? rob_val_28 : _GEN_10529; // @[rob.scala 515:{16,16}]
  wire  _GEN_10531 = 5'h1d == io_wb_resps_2_bits_uop_rob_idx ? rob_val_29 : _GEN_10530; // @[rob.scala 515:{16,16}]
  wire  _GEN_10532 = 5'h1e == io_wb_resps_2_bits_uop_rob_idx ? rob_val_30 : _GEN_10531; // @[rob.scala 515:{16,16}]
  wire  _GEN_10533 = 5'h1f == io_wb_resps_2_bits_uop_rob_idx ? rob_val_31 : _GEN_10532; // @[rob.scala 515:{16,16}]
  wire  _T_349 = ~_GEN_10533; // @[rob.scala 515:16]
  wire  _GEN_10535 = 5'h1 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_1 : rob_bsy_0; // @[rob.scala 518:{16,16}]
  wire  _GEN_10536 = 5'h2 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_2 : _GEN_10535; // @[rob.scala 518:{16,16}]
  wire  _GEN_10537 = 5'h3 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_3 : _GEN_10536; // @[rob.scala 518:{16,16}]
  wire  _GEN_10538 = 5'h4 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_4 : _GEN_10537; // @[rob.scala 518:{16,16}]
  wire  _GEN_10539 = 5'h5 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_5 : _GEN_10538; // @[rob.scala 518:{16,16}]
  wire  _GEN_10540 = 5'h6 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_6 : _GEN_10539; // @[rob.scala 518:{16,16}]
  wire  _GEN_10541 = 5'h7 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_7 : _GEN_10540; // @[rob.scala 518:{16,16}]
  wire  _GEN_10542 = 5'h8 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_8 : _GEN_10541; // @[rob.scala 518:{16,16}]
  wire  _GEN_10543 = 5'h9 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_9 : _GEN_10542; // @[rob.scala 518:{16,16}]
  wire  _GEN_10544 = 5'ha == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_10 : _GEN_10543; // @[rob.scala 518:{16,16}]
  wire  _GEN_10545 = 5'hb == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_11 : _GEN_10544; // @[rob.scala 518:{16,16}]
  wire  _GEN_10546 = 5'hc == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_12 : _GEN_10545; // @[rob.scala 518:{16,16}]
  wire  _GEN_10547 = 5'hd == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_13 : _GEN_10546; // @[rob.scala 518:{16,16}]
  wire  _GEN_10548 = 5'he == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_14 : _GEN_10547; // @[rob.scala 518:{16,16}]
  wire  _GEN_10549 = 5'hf == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_15 : _GEN_10548; // @[rob.scala 518:{16,16}]
  wire  _GEN_10550 = 5'h10 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_16 : _GEN_10549; // @[rob.scala 518:{16,16}]
  wire  _GEN_10551 = 5'h11 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_17 : _GEN_10550; // @[rob.scala 518:{16,16}]
  wire  _GEN_10552 = 5'h12 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_18 : _GEN_10551; // @[rob.scala 518:{16,16}]
  wire  _GEN_10553 = 5'h13 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_19 : _GEN_10552; // @[rob.scala 518:{16,16}]
  wire  _GEN_10554 = 5'h14 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_20 : _GEN_10553; // @[rob.scala 518:{16,16}]
  wire  _GEN_10555 = 5'h15 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_21 : _GEN_10554; // @[rob.scala 518:{16,16}]
  wire  _GEN_10556 = 5'h16 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_22 : _GEN_10555; // @[rob.scala 518:{16,16}]
  wire  _GEN_10557 = 5'h17 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_23 : _GEN_10556; // @[rob.scala 518:{16,16}]
  wire  _GEN_10558 = 5'h18 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_24 : _GEN_10557; // @[rob.scala 518:{16,16}]
  wire  _GEN_10559 = 5'h19 == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_25 : _GEN_10558; // @[rob.scala 518:{16,16}]
  wire  _GEN_10560 = 5'h1a == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_26 : _GEN_10559; // @[rob.scala 518:{16,16}]
  wire  _GEN_10561 = 5'h1b == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_27 : _GEN_10560; // @[rob.scala 518:{16,16}]
  wire  _GEN_10562 = 5'h1c == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_28 : _GEN_10561; // @[rob.scala 518:{16,16}]
  wire  _GEN_10563 = 5'h1d == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_29 : _GEN_10562; // @[rob.scala 518:{16,16}]
  wire  _GEN_10564 = 5'h1e == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_30 : _GEN_10563; // @[rob.scala 518:{16,16}]
  wire  _GEN_10565 = 5'h1f == io_wb_resps_2_bits_uop_rob_idx ? rob_bsy_31 : _GEN_10564; // @[rob.scala 518:{16,16}]
  wire  _T_357 = ~_GEN_10565; // @[rob.scala 518:16]
  wire  _GEN_10567 = 5'h1 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_1_ldst_val : rob_uop_0_ldst_val; // @[rob.scala 520:{72,72}]
  wire  _GEN_10568 = 5'h2 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_2_ldst_val : _GEN_10567; // @[rob.scala 520:{72,72}]
  wire  _GEN_10569 = 5'h3 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_3_ldst_val : _GEN_10568; // @[rob.scala 520:{72,72}]
  wire  _GEN_10570 = 5'h4 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_4_ldst_val : _GEN_10569; // @[rob.scala 520:{72,72}]
  wire  _GEN_10571 = 5'h5 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_5_ldst_val : _GEN_10570; // @[rob.scala 520:{72,72}]
  wire  _GEN_10572 = 5'h6 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_6_ldst_val : _GEN_10571; // @[rob.scala 520:{72,72}]
  wire  _GEN_10573 = 5'h7 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_7_ldst_val : _GEN_10572; // @[rob.scala 520:{72,72}]
  wire  _GEN_10574 = 5'h8 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_8_ldst_val : _GEN_10573; // @[rob.scala 520:{72,72}]
  wire  _GEN_10575 = 5'h9 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_9_ldst_val : _GEN_10574; // @[rob.scala 520:{72,72}]
  wire  _GEN_10576 = 5'ha == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_10_ldst_val : _GEN_10575; // @[rob.scala 520:{72,72}]
  wire  _GEN_10577 = 5'hb == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_11_ldst_val : _GEN_10576; // @[rob.scala 520:{72,72}]
  wire  _GEN_10578 = 5'hc == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_12_ldst_val : _GEN_10577; // @[rob.scala 520:{72,72}]
  wire  _GEN_10579 = 5'hd == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_13_ldst_val : _GEN_10578; // @[rob.scala 520:{72,72}]
  wire  _GEN_10580 = 5'he == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_14_ldst_val : _GEN_10579; // @[rob.scala 520:{72,72}]
  wire  _GEN_10581 = 5'hf == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_15_ldst_val : _GEN_10580; // @[rob.scala 520:{72,72}]
  wire  _GEN_10582 = 5'h10 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_16_ldst_val : _GEN_10581; // @[rob.scala 520:{72,72}]
  wire  _GEN_10583 = 5'h11 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_17_ldst_val : _GEN_10582; // @[rob.scala 520:{72,72}]
  wire  _GEN_10584 = 5'h12 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_18_ldst_val : _GEN_10583; // @[rob.scala 520:{72,72}]
  wire  _GEN_10585 = 5'h13 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_19_ldst_val : _GEN_10584; // @[rob.scala 520:{72,72}]
  wire  _GEN_10586 = 5'h14 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_20_ldst_val : _GEN_10585; // @[rob.scala 520:{72,72}]
  wire  _GEN_10587 = 5'h15 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_21_ldst_val : _GEN_10586; // @[rob.scala 520:{72,72}]
  wire  _GEN_10588 = 5'h16 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_22_ldst_val : _GEN_10587; // @[rob.scala 520:{72,72}]
  wire  _GEN_10589 = 5'h17 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_23_ldst_val : _GEN_10588; // @[rob.scala 520:{72,72}]
  wire  _GEN_10590 = 5'h18 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_24_ldst_val : _GEN_10589; // @[rob.scala 520:{72,72}]
  wire  _GEN_10591 = 5'h19 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_25_ldst_val : _GEN_10590; // @[rob.scala 520:{72,72}]
  wire  _GEN_10592 = 5'h1a == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_26_ldst_val : _GEN_10591; // @[rob.scala 520:{72,72}]
  wire  _GEN_10593 = 5'h1b == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_27_ldst_val : _GEN_10592; // @[rob.scala 520:{72,72}]
  wire  _GEN_10594 = 5'h1c == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_28_ldst_val : _GEN_10593; // @[rob.scala 520:{72,72}]
  wire  _GEN_10595 = 5'h1d == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_29_ldst_val : _GEN_10594; // @[rob.scala 520:{72,72}]
  wire  _GEN_10596 = 5'h1e == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_30_ldst_val : _GEN_10595; // @[rob.scala 520:{72,72}]
  wire  _GEN_10597 = 5'h1f == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_31_ldst_val : _GEN_10596; // @[rob.scala 520:{72,72}]
  wire  _T_365 = io_wb_resps_2_valid & _GEN_10597; // @[rob.scala 520:72]
  wire [5:0] _GEN_10599 = 5'h1 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_1_pdst : rob_uop_0_pdst; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10600 = 5'h2 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_2_pdst : _GEN_10599; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10601 = 5'h3 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_3_pdst : _GEN_10600; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10602 = 5'h4 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_4_pdst : _GEN_10601; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10603 = 5'h5 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_5_pdst : _GEN_10602; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10604 = 5'h6 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_6_pdst : _GEN_10603; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10605 = 5'h7 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_7_pdst : _GEN_10604; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10606 = 5'h8 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_8_pdst : _GEN_10605; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10607 = 5'h9 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_9_pdst : _GEN_10606; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10608 = 5'ha == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_10_pdst : _GEN_10607; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10609 = 5'hb == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_11_pdst : _GEN_10608; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10610 = 5'hc == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_12_pdst : _GEN_10609; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10611 = 5'hd == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_13_pdst : _GEN_10610; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10612 = 5'he == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_14_pdst : _GEN_10611; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10613 = 5'hf == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_15_pdst : _GEN_10612; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10614 = 5'h10 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_16_pdst : _GEN_10613; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10615 = 5'h11 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_17_pdst : _GEN_10614; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10616 = 5'h12 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_18_pdst : _GEN_10615; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10617 = 5'h13 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_19_pdst : _GEN_10616; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10618 = 5'h14 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_20_pdst : _GEN_10617; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10619 = 5'h15 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_21_pdst : _GEN_10618; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10620 = 5'h16 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_22_pdst : _GEN_10619; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10621 = 5'h17 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_23_pdst : _GEN_10620; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10622 = 5'h18 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_24_pdst : _GEN_10621; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10623 = 5'h19 == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_25_pdst : _GEN_10622; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10624 = 5'h1a == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_26_pdst : _GEN_10623; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10625 = 5'h1b == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_27_pdst : _GEN_10624; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10626 = 5'h1c == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_28_pdst : _GEN_10625; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10627 = 5'h1d == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_29_pdst : _GEN_10626; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10628 = 5'h1e == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_30_pdst : _GEN_10627; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10629 = 5'h1f == io_wb_resps_2_bits_uop_rob_idx ? rob_uop_31_pdst : _GEN_10628; // @[rob.scala 521:{51,51}]
  wire  _T_367 = _T_365 & _GEN_10629 != io_wb_resps_2_bits_uop_pdst; // @[rob.scala 521:34]
  wire  _GEN_10636 = 5'h1 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_1 : rob_val_0; // @[rob.scala 515:{16,16}]
  wire  _GEN_10637 = 5'h2 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_2 : _GEN_10636; // @[rob.scala 515:{16,16}]
  wire  _GEN_10638 = 5'h3 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_3 : _GEN_10637; // @[rob.scala 515:{16,16}]
  wire  _GEN_10639 = 5'h4 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_4 : _GEN_10638; // @[rob.scala 515:{16,16}]
  wire  _GEN_10640 = 5'h5 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_5 : _GEN_10639; // @[rob.scala 515:{16,16}]
  wire  _GEN_10641 = 5'h6 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_6 : _GEN_10640; // @[rob.scala 515:{16,16}]
  wire  _GEN_10642 = 5'h7 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_7 : _GEN_10641; // @[rob.scala 515:{16,16}]
  wire  _GEN_10643 = 5'h8 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_8 : _GEN_10642; // @[rob.scala 515:{16,16}]
  wire  _GEN_10644 = 5'h9 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_9 : _GEN_10643; // @[rob.scala 515:{16,16}]
  wire  _GEN_10645 = 5'ha == io_wb_resps_3_bits_uop_rob_idx ? rob_val_10 : _GEN_10644; // @[rob.scala 515:{16,16}]
  wire  _GEN_10646 = 5'hb == io_wb_resps_3_bits_uop_rob_idx ? rob_val_11 : _GEN_10645; // @[rob.scala 515:{16,16}]
  wire  _GEN_10647 = 5'hc == io_wb_resps_3_bits_uop_rob_idx ? rob_val_12 : _GEN_10646; // @[rob.scala 515:{16,16}]
  wire  _GEN_10648 = 5'hd == io_wb_resps_3_bits_uop_rob_idx ? rob_val_13 : _GEN_10647; // @[rob.scala 515:{16,16}]
  wire  _GEN_10649 = 5'he == io_wb_resps_3_bits_uop_rob_idx ? rob_val_14 : _GEN_10648; // @[rob.scala 515:{16,16}]
  wire  _GEN_10650 = 5'hf == io_wb_resps_3_bits_uop_rob_idx ? rob_val_15 : _GEN_10649; // @[rob.scala 515:{16,16}]
  wire  _GEN_10651 = 5'h10 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_16 : _GEN_10650; // @[rob.scala 515:{16,16}]
  wire  _GEN_10652 = 5'h11 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_17 : _GEN_10651; // @[rob.scala 515:{16,16}]
  wire  _GEN_10653 = 5'h12 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_18 : _GEN_10652; // @[rob.scala 515:{16,16}]
  wire  _GEN_10654 = 5'h13 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_19 : _GEN_10653; // @[rob.scala 515:{16,16}]
  wire  _GEN_10655 = 5'h14 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_20 : _GEN_10654; // @[rob.scala 515:{16,16}]
  wire  _GEN_10656 = 5'h15 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_21 : _GEN_10655; // @[rob.scala 515:{16,16}]
  wire  _GEN_10657 = 5'h16 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_22 : _GEN_10656; // @[rob.scala 515:{16,16}]
  wire  _GEN_10658 = 5'h17 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_23 : _GEN_10657; // @[rob.scala 515:{16,16}]
  wire  _GEN_10659 = 5'h18 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_24 : _GEN_10658; // @[rob.scala 515:{16,16}]
  wire  _GEN_10660 = 5'h19 == io_wb_resps_3_bits_uop_rob_idx ? rob_val_25 : _GEN_10659; // @[rob.scala 515:{16,16}]
  wire  _GEN_10661 = 5'h1a == io_wb_resps_3_bits_uop_rob_idx ? rob_val_26 : _GEN_10660; // @[rob.scala 515:{16,16}]
  wire  _GEN_10662 = 5'h1b == io_wb_resps_3_bits_uop_rob_idx ? rob_val_27 : _GEN_10661; // @[rob.scala 515:{16,16}]
  wire  _GEN_10663 = 5'h1c == io_wb_resps_3_bits_uop_rob_idx ? rob_val_28 : _GEN_10662; // @[rob.scala 515:{16,16}]
  wire  _GEN_10664 = 5'h1d == io_wb_resps_3_bits_uop_rob_idx ? rob_val_29 : _GEN_10663; // @[rob.scala 515:{16,16}]
  wire  _GEN_10665 = 5'h1e == io_wb_resps_3_bits_uop_rob_idx ? rob_val_30 : _GEN_10664; // @[rob.scala 515:{16,16}]
  wire  _GEN_10666 = 5'h1f == io_wb_resps_3_bits_uop_rob_idx ? rob_val_31 : _GEN_10665; // @[rob.scala 515:{16,16}]
  wire  _T_377 = ~_GEN_10666; // @[rob.scala 515:16]
  wire  _GEN_10668 = 5'h1 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_1 : rob_bsy_0; // @[rob.scala 518:{16,16}]
  wire  _GEN_10669 = 5'h2 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_2 : _GEN_10668; // @[rob.scala 518:{16,16}]
  wire  _GEN_10670 = 5'h3 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_3 : _GEN_10669; // @[rob.scala 518:{16,16}]
  wire  _GEN_10671 = 5'h4 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_4 : _GEN_10670; // @[rob.scala 518:{16,16}]
  wire  _GEN_10672 = 5'h5 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_5 : _GEN_10671; // @[rob.scala 518:{16,16}]
  wire  _GEN_10673 = 5'h6 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_6 : _GEN_10672; // @[rob.scala 518:{16,16}]
  wire  _GEN_10674 = 5'h7 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_7 : _GEN_10673; // @[rob.scala 518:{16,16}]
  wire  _GEN_10675 = 5'h8 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_8 : _GEN_10674; // @[rob.scala 518:{16,16}]
  wire  _GEN_10676 = 5'h9 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_9 : _GEN_10675; // @[rob.scala 518:{16,16}]
  wire  _GEN_10677 = 5'ha == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_10 : _GEN_10676; // @[rob.scala 518:{16,16}]
  wire  _GEN_10678 = 5'hb == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_11 : _GEN_10677; // @[rob.scala 518:{16,16}]
  wire  _GEN_10679 = 5'hc == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_12 : _GEN_10678; // @[rob.scala 518:{16,16}]
  wire  _GEN_10680 = 5'hd == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_13 : _GEN_10679; // @[rob.scala 518:{16,16}]
  wire  _GEN_10681 = 5'he == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_14 : _GEN_10680; // @[rob.scala 518:{16,16}]
  wire  _GEN_10682 = 5'hf == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_15 : _GEN_10681; // @[rob.scala 518:{16,16}]
  wire  _GEN_10683 = 5'h10 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_16 : _GEN_10682; // @[rob.scala 518:{16,16}]
  wire  _GEN_10684 = 5'h11 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_17 : _GEN_10683; // @[rob.scala 518:{16,16}]
  wire  _GEN_10685 = 5'h12 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_18 : _GEN_10684; // @[rob.scala 518:{16,16}]
  wire  _GEN_10686 = 5'h13 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_19 : _GEN_10685; // @[rob.scala 518:{16,16}]
  wire  _GEN_10687 = 5'h14 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_20 : _GEN_10686; // @[rob.scala 518:{16,16}]
  wire  _GEN_10688 = 5'h15 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_21 : _GEN_10687; // @[rob.scala 518:{16,16}]
  wire  _GEN_10689 = 5'h16 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_22 : _GEN_10688; // @[rob.scala 518:{16,16}]
  wire  _GEN_10690 = 5'h17 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_23 : _GEN_10689; // @[rob.scala 518:{16,16}]
  wire  _GEN_10691 = 5'h18 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_24 : _GEN_10690; // @[rob.scala 518:{16,16}]
  wire  _GEN_10692 = 5'h19 == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_25 : _GEN_10691; // @[rob.scala 518:{16,16}]
  wire  _GEN_10693 = 5'h1a == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_26 : _GEN_10692; // @[rob.scala 518:{16,16}]
  wire  _GEN_10694 = 5'h1b == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_27 : _GEN_10693; // @[rob.scala 518:{16,16}]
  wire  _GEN_10695 = 5'h1c == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_28 : _GEN_10694; // @[rob.scala 518:{16,16}]
  wire  _GEN_10696 = 5'h1d == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_29 : _GEN_10695; // @[rob.scala 518:{16,16}]
  wire  _GEN_10697 = 5'h1e == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_30 : _GEN_10696; // @[rob.scala 518:{16,16}]
  wire  _GEN_10698 = 5'h1f == io_wb_resps_3_bits_uop_rob_idx ? rob_bsy_31 : _GEN_10697; // @[rob.scala 518:{16,16}]
  wire  _T_385 = ~_GEN_10698; // @[rob.scala 518:16]
  wire  _GEN_10700 = 5'h1 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_1_ldst_val : rob_uop_0_ldst_val; // @[rob.scala 520:{72,72}]
  wire  _GEN_10701 = 5'h2 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_2_ldst_val : _GEN_10700; // @[rob.scala 520:{72,72}]
  wire  _GEN_10702 = 5'h3 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_3_ldst_val : _GEN_10701; // @[rob.scala 520:{72,72}]
  wire  _GEN_10703 = 5'h4 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_4_ldst_val : _GEN_10702; // @[rob.scala 520:{72,72}]
  wire  _GEN_10704 = 5'h5 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_5_ldst_val : _GEN_10703; // @[rob.scala 520:{72,72}]
  wire  _GEN_10705 = 5'h6 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_6_ldst_val : _GEN_10704; // @[rob.scala 520:{72,72}]
  wire  _GEN_10706 = 5'h7 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_7_ldst_val : _GEN_10705; // @[rob.scala 520:{72,72}]
  wire  _GEN_10707 = 5'h8 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_8_ldst_val : _GEN_10706; // @[rob.scala 520:{72,72}]
  wire  _GEN_10708 = 5'h9 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_9_ldst_val : _GEN_10707; // @[rob.scala 520:{72,72}]
  wire  _GEN_10709 = 5'ha == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_10_ldst_val : _GEN_10708; // @[rob.scala 520:{72,72}]
  wire  _GEN_10710 = 5'hb == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_11_ldst_val : _GEN_10709; // @[rob.scala 520:{72,72}]
  wire  _GEN_10711 = 5'hc == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_12_ldst_val : _GEN_10710; // @[rob.scala 520:{72,72}]
  wire  _GEN_10712 = 5'hd == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_13_ldst_val : _GEN_10711; // @[rob.scala 520:{72,72}]
  wire  _GEN_10713 = 5'he == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_14_ldst_val : _GEN_10712; // @[rob.scala 520:{72,72}]
  wire  _GEN_10714 = 5'hf == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_15_ldst_val : _GEN_10713; // @[rob.scala 520:{72,72}]
  wire  _GEN_10715 = 5'h10 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_16_ldst_val : _GEN_10714; // @[rob.scala 520:{72,72}]
  wire  _GEN_10716 = 5'h11 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_17_ldst_val : _GEN_10715; // @[rob.scala 520:{72,72}]
  wire  _GEN_10717 = 5'h12 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_18_ldst_val : _GEN_10716; // @[rob.scala 520:{72,72}]
  wire  _GEN_10718 = 5'h13 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_19_ldst_val : _GEN_10717; // @[rob.scala 520:{72,72}]
  wire  _GEN_10719 = 5'h14 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_20_ldst_val : _GEN_10718; // @[rob.scala 520:{72,72}]
  wire  _GEN_10720 = 5'h15 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_21_ldst_val : _GEN_10719; // @[rob.scala 520:{72,72}]
  wire  _GEN_10721 = 5'h16 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_22_ldst_val : _GEN_10720; // @[rob.scala 520:{72,72}]
  wire  _GEN_10722 = 5'h17 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_23_ldst_val : _GEN_10721; // @[rob.scala 520:{72,72}]
  wire  _GEN_10723 = 5'h18 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_24_ldst_val : _GEN_10722; // @[rob.scala 520:{72,72}]
  wire  _GEN_10724 = 5'h19 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_25_ldst_val : _GEN_10723; // @[rob.scala 520:{72,72}]
  wire  _GEN_10725 = 5'h1a == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_26_ldst_val : _GEN_10724; // @[rob.scala 520:{72,72}]
  wire  _GEN_10726 = 5'h1b == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_27_ldst_val : _GEN_10725; // @[rob.scala 520:{72,72}]
  wire  _GEN_10727 = 5'h1c == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_28_ldst_val : _GEN_10726; // @[rob.scala 520:{72,72}]
  wire  _GEN_10728 = 5'h1d == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_29_ldst_val : _GEN_10727; // @[rob.scala 520:{72,72}]
  wire  _GEN_10729 = 5'h1e == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_30_ldst_val : _GEN_10728; // @[rob.scala 520:{72,72}]
  wire  _GEN_10730 = 5'h1f == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_31_ldst_val : _GEN_10729; // @[rob.scala 520:{72,72}]
  wire  _T_393 = io_wb_resps_3_valid & _GEN_10730; // @[rob.scala 520:72]
  wire [5:0] _GEN_10732 = 5'h1 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_1_pdst : rob_uop_0_pdst; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10733 = 5'h2 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_2_pdst : _GEN_10732; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10734 = 5'h3 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_3_pdst : _GEN_10733; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10735 = 5'h4 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_4_pdst : _GEN_10734; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10736 = 5'h5 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_5_pdst : _GEN_10735; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10737 = 5'h6 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_6_pdst : _GEN_10736; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10738 = 5'h7 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_7_pdst : _GEN_10737; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10739 = 5'h8 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_8_pdst : _GEN_10738; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10740 = 5'h9 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_9_pdst : _GEN_10739; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10741 = 5'ha == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_10_pdst : _GEN_10740; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10742 = 5'hb == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_11_pdst : _GEN_10741; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10743 = 5'hc == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_12_pdst : _GEN_10742; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10744 = 5'hd == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_13_pdst : _GEN_10743; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10745 = 5'he == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_14_pdst : _GEN_10744; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10746 = 5'hf == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_15_pdst : _GEN_10745; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10747 = 5'h10 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_16_pdst : _GEN_10746; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10748 = 5'h11 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_17_pdst : _GEN_10747; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10749 = 5'h12 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_18_pdst : _GEN_10748; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10750 = 5'h13 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_19_pdst : _GEN_10749; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10751 = 5'h14 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_20_pdst : _GEN_10750; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10752 = 5'h15 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_21_pdst : _GEN_10751; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10753 = 5'h16 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_22_pdst : _GEN_10752; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10754 = 5'h17 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_23_pdst : _GEN_10753; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10755 = 5'h18 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_24_pdst : _GEN_10754; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10756 = 5'h19 == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_25_pdst : _GEN_10755; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10757 = 5'h1a == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_26_pdst : _GEN_10756; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10758 = 5'h1b == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_27_pdst : _GEN_10757; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10759 = 5'h1c == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_28_pdst : _GEN_10758; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10760 = 5'h1d == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_29_pdst : _GEN_10759; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10761 = 5'h1e == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_30_pdst : _GEN_10760; // @[rob.scala 521:{51,51}]
  wire [5:0] _GEN_10762 = 5'h1f == io_wb_resps_3_bits_uop_rob_idx ? rob_uop_31_pdst : _GEN_10761; // @[rob.scala 521:{51,51}]
  wire  _T_395 = _T_393 & _GEN_10762 != io_wb_resps_3_bits_uop_pdst; // @[rob.scala 521:34]
  reg  _T_406; // @[rob.scala 540:131]
  wire  will_throw_exception = can_throw_exception_0 & _T_415; // @[rob.scala 545:52]
  wire  is_mini_exception = io_com_xcpt_bits_cause == 64'h10; // @[rob.scala 556:50]
  wire  _T_421 = will_throw_exception & ~is_mini_exception; // @[rob.scala 557:41]
  wire [23:0] _T_424 = r_xcpt_badvaddr[39] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  wire  insn_sys_pc2epc = rob_head_vals_0 & io_commit_uops_0_is_sys_pc2epc; // @[rob.scala 562:31]
  wire  refetch_inst = will_throw_exception | insn_sys_pc2epc; // @[rob.scala 564:39]
  wire  flush_commit_mask_0 = io_commit_valids_0 & io_commit_uops_0_flush_on_commit; // @[rob.scala 571:75]
  wire  flush_val = will_throw_exception | flush_commit_mask_0; // @[rob.scala 573:36]
  wire  _T_434 = flush_commit_mask_0 & io_commit_uops_0_uopc == 7'h6a; // @[rob.scala 588:62]
  wire [2:0] _T_436 = refetch_inst ? 3'h2 : 3'h4; // @[rob.scala 175:10]
  wire [2:0] _T_437 = _T_421 ? 3'h1 : _T_436; // @[rob.scala 174:10]
  wire [2:0] _T_438 = _T_434 ? 3'h3 : _T_437; // @[rob.scala 173:10]
  wire  _T_440 = io_commit_valids_0 & io_commit_uops_0_fp_val; // @[rob.scala 601:27]
  wire  _T_441 = ~io_commit_uops_0_uses_stq; // @[rob.scala 603:7]
  wire  fflags_val_0 = _T_440 & _T_441; // @[rob.scala 602:32]
  wire [4:0] rob_head_fflags_0 = rob_fflags__T_221_data; // @[rob.scala 252:33 483:26]
  wire  _T_444 = ~io_commit_uops_0_fp_val; // @[rob.scala 608:14]
  wire  _T_445 = io_commit_valids_0 & _T_444; // @[rob.scala 607:35]
  wire  _T_446 = rob_head_fflags_0 != 5'h0; // @[rob.scala 609:33]
  wire  _T_447 = _T_445 & _T_446; // @[rob.scala 608:40]
  wire  _T_453 = io_commit_uops_0_uses_ldq | io_commit_uops_0_uses_stq; // @[rob.scala 613:42]
  wire  _T_454 = _T_440 & _T_453; // @[rob.scala 612:39]
  wire  _T_456 = _T_454 & _T_446; // @[rob.scala 613:73]
  wire  enq_xcpts_0 = io_enq_valids_0 & io_enq_uops_0_exception; // @[rob.scala 628:38]
  wire  _T_466 = ~r_xcpt_val; // @[rob.scala 635:13]
  wire  _T_471 = io_lxcpt_bits_uop_rob_idx < r_xcpt_uop_rob_idx ^ io_lxcpt_bits_uop_rob_idx < rob_head ^
    r_xcpt_uop_rob_idx < rob_head; // @[util.scala 363:72]
  wire  _GEN_10763 = ~r_xcpt_val | _T_471 | r_xcpt_val; // @[rob.scala 258:33 635:93 636:33]
  wire [7:0] _GEN_10818 = ~r_xcpt_val | _T_471 ? io_lxcpt_bits_uop_br_mask : r_xcpt_uop_br_mask; // @[rob.scala 625:17 635:93 637:33]
  wire [39:0] _T_475 = ~io_xcpt_fetch_pc; // @[util.scala 237:7]
  wire [39:0] _T_476 = _T_475 | 40'h3f; // @[util.scala 237:11]
  wire [39:0] _T_477 = ~_T_476; // @[util.scala 237:5]
  wire [39:0] _GEN_11185 = {{34'd0}, io_enq_uops_0_pc_lob}; // @[rob.scala 647:76]
  wire [39:0] _T_478 = _T_477 | _GEN_11185; // @[rob.scala 647:76]
  wire  _GEN_10844 = _T_466 & enq_xcpts_0 | r_xcpt_val; // @[rob.scala 641:56 645:23 258:33]
  wire [7:0] _GEN_10899 = _T_466 & enq_xcpts_0 ? io_enq_uops_0_br_mask : r_xcpt_uop_br_mask; // @[rob.scala 625:17 641:56 646:23]
  wire [7:0] _GEN_10980 = io_lxcpt_valid ? _GEN_10818 : _GEN_10899; // @[rob.scala 632:27]
  wire [7:0] next_xcpt_uop_br_mask = ~(io_flush_valid | will_throw_exception) & rob_state != 2'h2 ? _GEN_10980 :
    r_xcpt_uop_br_mask; // @[rob.scala 625:17 631:76]
  wire [7:0] _T_481 = io_brupdate_b1_mispredict_mask & next_xcpt_uop_br_mask; // @[util.scala 118:51]
  wire  _T_482 = _T_481 != 8'h0; // @[util.scala 118:59]
  wire  _T_599 = rob_head == rob_tail; // @[rob.scala 788:27]
  wire  empty = rob_head == rob_tail & ~rob_head_vals_0; // @[rob.scala 788:41]
  reg  r_partial_row; // @[rob.scala 677:30]
  wire  _T_503 = ~(will_commit_0 ^ rob_head_vals_0); // @[rob.scala 685:50]
  wire  _T_504 = io_commit_valids_0 & _T_503; // @[rob.scala 684:39]
  wire  _T_507 = ~maybe_full; // @[rob.scala 686:49]
  wire  _T_509 = ~(r_partial_row & _T_599 & ~maybe_full); // @[rob.scala 686:5]
  wire  finished_committing_row = _T_504 & _T_509; // @[rob.scala 685:59]
  wire [4:0] _T_511 = rob_head + 5'h1; // @[util.scala 203:14]
  reg  pnr_maybe_at_tail; // @[rob.scala 714:36]
  wire  _T_515 = rob_state == 2'h1; // @[rob.scala 716:33]
  wire  safe_to_inc = rob_state == 2'h1 | rob_state == 2'h3; // @[rob.scala 716:46]
  wire  do_inc_row = ~rob_pnr_unsafe_0 & (rob_pnr != rob_tail | full & ~pnr_maybe_at_tail); // @[rob.scala 717:52]
  wire [4:0] _T_526 = rob_pnr + 5'h1; // @[util.scala 203:14]
  wire  rob_deq = _T & (rob_tail != rob_head | maybe_full) | finished_committing_row; // @[rob.scala 750:76 754:13]
  wire  _T_542 = ~rob_deq; // @[rob.scala 736:26]
  wire  _T_549 = rob_pnr < rob_head ^ rob_pnr < rob_tail ^ rob_head < rob_tail; // @[util.scala 363:72]
  wire  _T_560 = rob_tail < rob_pnr ^ rob_tail < rob_head ^ rob_pnr < rob_head; // @[util.scala 363:72]
  wire [4:0] _T_571 = rob_tail - 5'h1; // @[util.scala 220:14]
  wire [4:0] _T_579 = io_brupdate_b2_uop_rob_idx + 5'h1; // @[util.scala 203:14]
  wire  _T_583 = io_enq_valids_0 & ~io_enq_partial_stall; // @[rob.scala 761:45]
  wire [4:0] _T_585 = rob_tail + 5'h1; // @[util.scala 203:14]
  wire [4:0] _GEN_11100 = io_enq_valids_0 & ~io_enq_partial_stall ? _T_585 : rob_tail; // @[rob.scala 761:71 762:18 228:29]
  wire  _GEN_11105 = io_brupdate_b2_mispredict ? 1'h0 : _T_583; // @[rob.scala 758:43]
  wire  _GEN_11108 = _T & _T_597 & _T_507 ? 1'h0 : _GEN_11105; // @[rob.scala 755:84]
  wire  rob_enq = _T & (rob_tail != rob_head | maybe_full) ? 1'h0 : _GEN_11108; // @[rob.scala 750:76]
  wire  _T_607 = 2'h0 == rob_state; // @[Conditional.scala 37:30]
  wire  _T_608 = 2'h1 == rob_state; // @[Conditional.scala 37:30]
  reg  _T_609; // @[rob.scala 808:30]
  reg  _T_610; // @[rob.scala 808:22]
  wire [1:0] _GEN_11113 = io_enq_valids_0 & io_enq_uops_0_is_unique ? 2'h3 : rob_state; // @[rob.scala 812:65 813:25 221:26]
  wire  _T_612 = 2'h2 == rob_state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_11115 = empty ? 2'h1 : rob_state; // @[rob.scala 819:22 820:21 221:26]
  wire  _T_613 = 2'h3 == rob_state; // @[Conditional.scala 37:30]
  reg  _T_614; // @[rob.scala 824:22]
  wire [1:0] _GEN_11116 = _T_614 ? 2'h2 : _GEN_11115; // @[rob.scala 824:42 825:21]
  wire [1:0] _GEN_11117 = _T_613 ? _GEN_11116 : rob_state; // @[Conditional.scala 39:67 rob.scala 221:26]
  wire  _T_616 = ~will_commit_0; // @[rob.scala 866:41]
  reg  _T_618; // @[rob.scala 865:40]
  assign rob_debug_inst_mem_0_rob_debug_inst_rdata_en = rob_debug_inst_mem_0_rob_debug_inst_rdata_en_pipe_0;
  assign rob_debug_inst_mem_0_rob_debug_inst_rdata_addr = rob_debug_inst_mem_0_rob_debug_inst_rdata_addr_pipe_0;
  assign rob_debug_inst_mem_0_rob_debug_inst_rdata_data =
    rob_debug_inst_mem_0[rob_debug_inst_mem_0_rob_debug_inst_rdata_addr]; // @[rob.scala 297:41]
  assign rob_debug_inst_mem_0__T_3_data = io_enq_uops_0_debug_inst;
  assign rob_debug_inst_mem_0__T_3_addr = rob_tail;
  assign rob_debug_inst_mem_0__T_3_mask = io_enq_valids_0;
  assign rob_debug_inst_mem_0__T_3_en = 1'h1;
  assign rob_fflags__T_221_en = 1'h1;
  assign rob_fflags__T_221_addr = rob_head;
  assign rob_fflags__T_221_data = rob_fflags[rob_fflags__T_221_addr]; // @[rob.scala 313:28]
  assign rob_fflags__T_15_data = 5'h0;
  assign rob_fflags__T_15_addr = rob_tail;
  assign rob_fflags__T_15_mask = 1'h1;
  assign rob_fflags__T_15_en = io_enq_valids_0;
  assign rob_fflags__T_59_data = io_fflags_0_bits_flags;
  assign rob_fflags__T_59_addr = io_fflags_0_bits_uop_rob_idx;
  assign rob_fflags__T_59_mask = 1'h1;
  assign rob_fflags__T_59_en = io_fflags_0_valid;
  assign rob_fflags__T_62_data = io_fflags_1_bits_flags;
  assign rob_fflags__T_62_addr = io_fflags_1_bits_uop_rob_idx;
  assign rob_fflags__T_62_mask = 1'h1;
  assign rob_fflags__T_62_en = io_fflags_1_valid;
  assign rob_debug_wdata__T_400_en = 1'h1;
  assign rob_debug_wdata__T_400_addr = rob_head;
  assign rob_debug_wdata__T_400_data = rob_debug_wdata[rob_debug_wdata__T_400_addr]; // @[rob.scala 315:30]
  assign rob_debug_wdata__T_290_data = io_debug_wb_wdata_0;
  assign rob_debug_wdata__T_290_addr = io_wb_resps_0_bits_uop_rob_idx;
  assign rob_debug_wdata__T_290_mask = 1'h1;
  assign rob_debug_wdata__T_290_en = io_debug_wb_valids_0;
  assign rob_debug_wdata__T_318_data = io_debug_wb_wdata_1;
  assign rob_debug_wdata__T_318_addr = io_wb_resps_1_bits_uop_rob_idx;
  assign rob_debug_wdata__T_318_mask = 1'h1;
  assign rob_debug_wdata__T_318_en = io_debug_wb_valids_1;
  assign rob_debug_wdata__T_346_data = io_debug_wb_wdata_2;
  assign rob_debug_wdata__T_346_addr = io_wb_resps_2_bits_uop_rob_idx;
  assign rob_debug_wdata__T_346_mask = 1'h1;
  assign rob_debug_wdata__T_346_en = io_debug_wb_valids_2;
  assign rob_debug_wdata__T_374_data = io_debug_wb_wdata_3;
  assign rob_debug_wdata__T_374_addr = io_wb_resps_3_bits_uop_rob_idx;
  assign rob_debug_wdata__T_374_mask = 1'h1;
  assign rob_debug_wdata__T_374_en = io_debug_wb_valids_3;
  assign io_rob_tail_idx = rob_tail; // @[rob.scala 791:19]
  assign io_rob_pnr_idx = rob_pnr; // @[rob.scala 792:19]
  assign io_rob_head_idx = rob_head; // @[rob.scala 790:19]
  assign io_commit_valids_0 = can_commit_0 & ~can_throw_exception_0 & ~_T_408; // @[rob.scala 547:70]
  assign io_commit_arch_valids_0 = will_commit_0 & ~_GEN_6932; // @[rob.scala 410:48]
  assign io_commit_uops_0_uopc = 5'h1f == com_idx ? rob_uop_31_uopc : _GEN_9459; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_inst = 5'h1f == com_idx ? rob_uop_31_inst : _GEN_9427; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_debug_inst = 5'h1f == com_idx ? rob_uop_31_debug_inst : _GEN_9395; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_is_rvc = 5'h1f == com_idx ? rob_uop_31_is_rvc : _GEN_9363; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_debug_pc = 5'h1f == com_idx ? rob_uop_31_debug_pc : _GEN_9331; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_iq_type = 5'h1f == com_idx ? rob_uop_31_iq_type : _GEN_9299; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_fu_code = 5'h1f == com_idx ? rob_uop_31_fu_code : _GEN_9267; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_ctrl_br_type = 5'h1f == com_idx ? rob_uop_31_ctrl_br_type : _GEN_9235; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_ctrl_op1_sel = 5'h1f == com_idx ? rob_uop_31_ctrl_op1_sel : _GEN_9203; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_ctrl_op2_sel = 5'h1f == com_idx ? rob_uop_31_ctrl_op2_sel : _GEN_9171; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_ctrl_imm_sel = 5'h1f == com_idx ? rob_uop_31_ctrl_imm_sel : _GEN_9139; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_ctrl_op_fcn = 5'h1f == com_idx ? rob_uop_31_ctrl_op_fcn : _GEN_9107; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_ctrl_fcn_dw = 5'h1f == com_idx ? rob_uop_31_ctrl_fcn_dw : _GEN_9075; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_ctrl_csr_cmd = 5'h1f == com_idx ? rob_uop_31_ctrl_csr_cmd : _GEN_9043; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_ctrl_is_load = 5'h1f == com_idx ? rob_uop_31_ctrl_is_load : _GEN_9011; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_ctrl_is_sta = 5'h1f == com_idx ? rob_uop_31_ctrl_is_sta : _GEN_8979; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_ctrl_is_std = 5'h1f == com_idx ? rob_uop_31_ctrl_is_std : _GEN_8947; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_iw_state = 5'h1f == com_idx ? rob_uop_31_iw_state : _GEN_8915; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_iw_p1_poisoned = 5'h1f == com_idx ? rob_uop_31_iw_p1_poisoned : _GEN_8883; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_iw_p2_poisoned = 5'h1f == com_idx ? rob_uop_31_iw_p2_poisoned : _GEN_8851; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_is_br = 5'h1f == com_idx ? rob_uop_31_is_br : _GEN_8819; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_is_jalr = 5'h1f == com_idx ? rob_uop_31_is_jalr : _GEN_8787; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_is_jal = 5'h1f == com_idx ? rob_uop_31_is_jal : _GEN_8755; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_is_sfb = 5'h1f == com_idx ? rob_uop_31_is_sfb : _GEN_8723; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_br_mask = 5'h1f == com_idx ? rob_uop_31_br_mask : _GEN_8691; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_br_tag = 5'h1f == com_idx ? rob_uop_31_br_tag : _GEN_8659; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_ftq_idx = 5'h1f == com_idx ? rob_uop_31_ftq_idx : _GEN_8627; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_edge_inst = 5'h1f == com_idx ? rob_uop_31_edge_inst : _GEN_8595; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_pc_lob = 5'h1f == com_idx ? rob_uop_31_pc_lob : _GEN_8563; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_taken = _T_79 ? io_brupdate_b2_taken : _GEN_8532; // @[rob.scala 411:25 418:58 420:36]
  assign io_commit_uops_0_imm_packed = 5'h1f == com_idx ? rob_uop_31_imm_packed : _GEN_8499; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_csr_addr = 5'h1f == com_idx ? rob_uop_31_csr_addr : _GEN_8467; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_rob_idx = 5'h1f == com_idx ? rob_uop_31_rob_idx : _GEN_8435; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_ldq_idx = 5'h1f == com_idx ? rob_uop_31_ldq_idx : _GEN_8403; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_stq_idx = 5'h1f == com_idx ? rob_uop_31_stq_idx : _GEN_8371; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_rxq_idx = 5'h1f == com_idx ? rob_uop_31_rxq_idx : _GEN_8339; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_pdst = 5'h1f == com_idx ? rob_uop_31_pdst : _GEN_8307; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_prs1 = 5'h1f == com_idx ? rob_uop_31_prs1 : _GEN_8275; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_prs2 = 5'h1f == com_idx ? rob_uop_31_prs2 : _GEN_8243; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_prs3 = 5'h1f == com_idx ? rob_uop_31_prs3 : _GEN_8211; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_ppred = 5'h1f == com_idx ? rob_uop_31_ppred : _GEN_8179; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_prs1_busy = 5'h1f == com_idx ? rob_uop_31_prs1_busy : _GEN_8147; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_prs2_busy = 5'h1f == com_idx ? rob_uop_31_prs2_busy : _GEN_8115; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_prs3_busy = 5'h1f == com_idx ? rob_uop_31_prs3_busy : _GEN_8083; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_ppred_busy = 5'h1f == com_idx ? rob_uop_31_ppred_busy : _GEN_8051; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_stale_pdst = 5'h1f == com_idx ? rob_uop_31_stale_pdst : _GEN_8019; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_exception = 5'h1f == com_idx ? rob_uop_31_exception : _GEN_7987; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_exc_cause = 5'h1f == com_idx ? rob_uop_31_exc_cause : _GEN_7955; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_bypassable = 5'h1f == com_idx ? rob_uop_31_bypassable : _GEN_7923; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_mem_cmd = 5'h1f == com_idx ? rob_uop_31_mem_cmd : _GEN_7891; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_mem_size = 5'h1f == com_idx ? rob_uop_31_mem_size : _GEN_7859; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_mem_signed = 5'h1f == com_idx ? rob_uop_31_mem_signed : _GEN_7827; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_is_fence = 5'h1f == com_idx ? rob_uop_31_is_fence : _GEN_7795; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_is_fencei = 5'h1f == com_idx ? rob_uop_31_is_fencei : _GEN_7763; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_is_amo = 5'h1f == com_idx ? rob_uop_31_is_amo : _GEN_7731; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_uses_ldq = 5'h1f == com_idx ? rob_uop_31_uses_ldq : _GEN_7699; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_uses_stq = 5'h1f == com_idx ? rob_uop_31_uses_stq : _GEN_7667; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_is_sys_pc2epc = 5'h1f == com_idx ? rob_uop_31_is_sys_pc2epc : _GEN_7635; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_is_unique = 5'h1f == com_idx ? rob_uop_31_is_unique : _GEN_7603; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_flush_on_commit = 5'h1f == com_idx ? rob_uop_31_flush_on_commit : _GEN_7571; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_ldst_is_rs1 = 5'h1f == com_idx ? rob_uop_31_ldst_is_rs1 : _GEN_7539; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_ldst = 5'h1f == com_idx ? rob_uop_31_ldst : _GEN_7507; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_lrs1 = 5'h1f == com_idx ? rob_uop_31_lrs1 : _GEN_7475; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_lrs2 = 5'h1f == com_idx ? rob_uop_31_lrs2 : _GEN_7443; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_lrs3 = 5'h1f == com_idx ? rob_uop_31_lrs3 : _GEN_7411; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_ldst_val = 5'h1f == com_idx ? rob_uop_31_ldst_val : _GEN_7379; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_dst_rtype = 5'h1f == com_idx ? rob_uop_31_dst_rtype : _GEN_7347; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_lrs1_rtype = 5'h1f == com_idx ? rob_uop_31_lrs1_rtype : _GEN_7315; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_lrs2_rtype = 5'h1f == com_idx ? rob_uop_31_lrs2_rtype : _GEN_7283; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_frs3_en = 5'h1f == com_idx ? rob_uop_31_frs3_en : _GEN_7251; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_fp_val = 5'h1f == com_idx ? rob_uop_31_fp_val : _GEN_7219; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_fp_single = 5'h1f == com_idx ? rob_uop_31_fp_single : _GEN_7187; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_xcpt_pf_if = 5'h1f == com_idx ? rob_uop_31_xcpt_pf_if : _GEN_7155; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_xcpt_ae_if = 5'h1f == com_idx ? rob_uop_31_xcpt_ae_if : _GEN_7123; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_xcpt_ma_if = 5'h1f == com_idx ? rob_uop_31_xcpt_ma_if : _GEN_7091; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_bp_debug_if = 5'h1f == com_idx ? rob_uop_31_bp_debug_if : _GEN_7059; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_bp_xcpt_if = 5'h1f == com_idx ? rob_uop_31_bp_xcpt_if : _GEN_7027; // @[rob.scala 411:{25,25}]
  assign io_commit_uops_0_debug_fsrc = _T_79 ? 2'h3 : _GEN_6996; // @[rob.scala 411:25 418:58 419:36]
  assign io_commit_uops_0_debug_tsrc = 5'h1f == com_idx ? rob_uop_31_debug_tsrc : _GEN_6963; // @[rob.scala 411:{25,25}]
  assign io_commit_fflags_valid = _T_440 & _T_441; // @[rob.scala 602:32]
  assign io_commit_fflags_bits = fflags_val_0 ? rob_head_fflags_0 : 5'h0; // @[rob.scala 605:21]
  assign io_commit_debug_insts_0 = rob_debug_inst_mem_0_rob_debug_inst_rdata_data; // @[rob.scala 412:30]
  assign io_commit_rbk_valids_0 = rbk_row & _GEN_9494; // @[rob.scala 427:40]
  assign io_commit_rollback = rob_state == 2'h2; // @[rob.scala 428:38]
  assign io_commit_debug_wdata_0 = rob_debug_wdata__T_400_data; // @[rob.scala 524:30]
  assign io_com_load_is_at_rob_head = _T_618; // @[rob.scala 865:30]
  assign io_com_xcpt_valid = will_throw_exception & ~is_mini_exception; // @[rob.scala 557:41]
  assign io_com_xcpt_bits_ftq_idx = io_commit_uops_0_ftq_idx; // @[rob.scala 566:30]
  assign io_com_xcpt_bits_edge_inst = io_commit_uops_0_edge_inst; // @[rob.scala 567:30]
  assign io_com_xcpt_bits_is_rvc = io_commit_uops_0_is_rvc; // @[rob.scala 568:30]
  assign io_com_xcpt_bits_pc_lob = io_commit_uops_0_pc_lob; // @[rob.scala 569:30]
  assign io_com_xcpt_bits_cause = r_xcpt_uop_exc_cause; // @[rob.scala 558:26]
  assign io_com_xcpt_bits_badvaddr = {_T_424,r_xcpt_badvaddr}; // @[Cat.scala 29:58]
  assign io_com_xcpt_bits_flush_typ = 3'h0;
  assign io_flush_valid = will_throw_exception | flush_commit_mask_0; // @[rob.scala 573:36]
  assign io_flush_bits_ftq_idx = io_commit_uops_0_ftq_idx; // @[rob.scala 578:22]
  assign io_flush_bits_edge_inst = io_commit_uops_0_edge_inst; // @[rob.scala 578:22]
  assign io_flush_bits_is_rvc = io_commit_uops_0_is_rvc; // @[rob.scala 578:22]
  assign io_flush_bits_pc_lob = io_commit_uops_0_pc_lob; // @[rob.scala 578:22]
  assign io_flush_bits_cause = 64'h0;
  assign io_flush_bits_badvaddr = 64'h0;
  assign io_flush_bits_flush_typ = ~flush_val ? 3'h0 : _T_438; // @[rob.scala 172:10]
  assign io_empty = rob_head == rob_tail & ~rob_head_vals_0; // @[rob.scala 788:41]
  assign io_ready = _T_515 & _T_81 & _T_466; // @[rob.scala 794:56]
  assign io_flush_frontend = r_xcpt_val; // @[rob.scala 261:21]
  always @(posedge clock) begin
    if (rob_debug_inst_mem_0__T_3_en & rob_debug_inst_mem_0__T_3_mask) begin
      rob_debug_inst_mem_0[rob_debug_inst_mem_0__T_3_addr] <= rob_debug_inst_mem_0__T_3_data; // @[rob.scala 297:41]
    end
    rob_debug_inst_mem_0_rob_debug_inst_rdata_en_pipe_0 <= _T_414 & _T_415;
    if (_T_414 & _T_415) begin
      rob_debug_inst_mem_0_rob_debug_inst_rdata_addr_pipe_0 <= rob_head;
    end
    if (rob_fflags__T_15_en & rob_fflags__T_15_mask) begin
      rob_fflags[rob_fflags__T_15_addr] <= rob_fflags__T_15_data; // @[rob.scala 313:28]
    end
    if (rob_fflags__T_59_en & rob_fflags__T_59_mask) begin
      rob_fflags[rob_fflags__T_59_addr] <= rob_fflags__T_59_data; // @[rob.scala 313:28]
    end
    if (rob_fflags__T_62_en & rob_fflags__T_62_mask) begin
      rob_fflags[rob_fflags__T_62_addr] <= rob_fflags__T_62_data; // @[rob.scala 313:28]
    end
    if (rob_debug_wdata__T_290_en & rob_debug_wdata__T_290_mask) begin
      rob_debug_wdata[rob_debug_wdata__T_290_addr] <= rob_debug_wdata__T_290_data; // @[rob.scala 315:30]
    end
    if (rob_debug_wdata__T_318_en & rob_debug_wdata__T_318_mask) begin
      rob_debug_wdata[rob_debug_wdata__T_318_addr] <= rob_debug_wdata__T_318_data; // @[rob.scala 315:30]
    end
    if (rob_debug_wdata__T_346_en & rob_debug_wdata__T_346_mask) begin
      rob_debug_wdata[rob_debug_wdata__T_346_addr] <= rob_debug_wdata__T_346_data; // @[rob.scala 315:30]
    end
    if (rob_debug_wdata__T_374_en & rob_debug_wdata__T_374_mask) begin
      rob_debug_wdata[rob_debug_wdata__T_374_addr] <= rob_debug_wdata__T_374_data; // @[rob.scala 315:30]
    end
    if (reset) begin // @[rob.scala 221:26]
      rob_state <= 2'h0; // @[rob.scala 221:26]
    end else if (_T_607) begin // @[Conditional.scala 40:58]
      rob_state <= 2'h1; // @[rob.scala 804:19]
    end else if (_T_608) begin // @[Conditional.scala 39:67]
      if (_T_610) begin // @[rob.scala 808:51]
        rob_state <= 2'h2; // @[rob.scala 809:21]
      end else begin
        rob_state <= _GEN_11113;
      end
    end else if (_T_612) begin // @[Conditional.scala 39:67]
      rob_state <= _GEN_11115;
    end else begin
      rob_state <= _GEN_11117;
    end
    if (reset) begin // @[rob.scala 224:29]
      rob_head <= 5'h0; // @[rob.scala 224:29]
    end else if (finished_committing_row) begin // @[rob.scala 688:34]
      rob_head <= _T_511; // @[rob.scala 689:18]
    end
    if (reset) begin // @[rob.scala 228:29]
      rob_tail <= 5'h0; // @[rob.scala 228:29]
    end else if (_T & (rob_tail != rob_head | maybe_full)) begin // @[rob.scala 750:76]
      rob_tail <= _T_571; // @[rob.scala 752:18]
    end else if (!(_T & _T_597 & _T_507)) begin // @[rob.scala 755:84]
      if (io_brupdate_b2_mispredict) begin // @[rob.scala 758:43]
        rob_tail <= _T_579; // @[rob.scala 759:18]
      end else begin
        rob_tail <= _GEN_11100;
      end
    end
    if (reset) begin // @[rob.scala 232:29]
      rob_pnr <= 5'h0; // @[rob.scala 232:29]
    end else if (empty & io_enq_valids_0) begin // @[rob.scala 718:50]
      rob_pnr <= rob_head; // @[rob.scala 723:19]
    end else if (safe_to_inc & do_inc_row) begin // @[rob.scala 725:45]
      rob_pnr <= _T_526; // @[rob.scala 726:19]
    end
    if (reset) begin // @[rob.scala 239:29]
      maybe_full <= 1'h0; // @[rob.scala 239:29]
    end else begin
      maybe_full <= _T_542 & (rob_enq | maybe_full) | io_brupdate_b1_mispredict_mask != 8'h0; // @[rob.scala 786:14]
    end
    if (reset) begin // @[rob.scala 258:33]
      r_xcpt_val <= 1'h0; // @[rob.scala 258:33]
    end else if (io_flush_valid | _T_482) begin // @[rob.scala 654:73]
      r_xcpt_val <= 1'h0; // @[rob.scala 655:16]
    end else if (~(io_flush_valid | will_throw_exception) & rob_state != 2'h2) begin // @[rob.scala 631:76]
      if (io_lxcpt_valid) begin // @[rob.scala 632:27]
        r_xcpt_val <= _GEN_10763;
      end else begin
        r_xcpt_val <= _GEN_10844;
      end
    end
    r_xcpt_uop_br_mask <= next_xcpt_uop_br_mask & _T_93; // @[util.scala 85:25]
    if (~(io_flush_valid | will_throw_exception) & rob_state != 2'h2) begin // @[rob.scala 631:76]
      if (io_lxcpt_valid) begin // @[rob.scala 632:27]
        if (~r_xcpt_val | _T_471) begin // @[rob.scala 635:93]
          r_xcpt_uop_rob_idx <= io_lxcpt_bits_uop_rob_idx; // @[rob.scala 637:33]
        end
      end else if (_T_466 & enq_xcpts_0) begin // @[rob.scala 641:56]
        r_xcpt_uop_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 646:23]
      end
    end
    if (~(io_flush_valid | will_throw_exception) & rob_state != 2'h2) begin // @[rob.scala 631:76]
      if (io_lxcpt_valid) begin // @[rob.scala 632:27]
        if (~r_xcpt_val | _T_471) begin // @[rob.scala 635:93]
          r_xcpt_uop_exc_cause <= {{59'd0}, io_lxcpt_bits_cause}; // @[rob.scala 638:33]
        end
      end else if (_T_466 & enq_xcpts_0) begin // @[rob.scala 641:56]
        r_xcpt_uop_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 646:23]
      end
    end
    if (~(io_flush_valid | will_throw_exception) & rob_state != 2'h2) begin // @[rob.scala 631:76]
      if (io_lxcpt_valid) begin // @[rob.scala 632:27]
        if (~r_xcpt_val | _T_471) begin // @[rob.scala 635:93]
          r_xcpt_badvaddr <= io_lxcpt_bits_badvaddr; // @[rob.scala 639:33]
        end
      end else if (_T_466 & enq_xcpts_0) begin // @[rob.scala 641:56]
        r_xcpt_badvaddr <= _T_478; // @[rob.scala 647:23]
      end
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_31 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h1f == rob_head) begin // @[rob.scala 476:25]
        rob_val_31 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_31 <= _GEN_9748;
      end
    end else begin
      rob_val_31 <= _GEN_9748;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_30 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h1e == rob_head) begin // @[rob.scala 476:25]
        rob_val_30 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_30 <= _GEN_9744;
      end
    end else begin
      rob_val_30 <= _GEN_9744;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_29 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h1d == rob_head) begin // @[rob.scala 476:25]
        rob_val_29 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_29 <= _GEN_9740;
      end
    end else begin
      rob_val_29 <= _GEN_9740;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_28 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h1c == rob_head) begin // @[rob.scala 476:25]
        rob_val_28 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_28 <= _GEN_9736;
      end
    end else begin
      rob_val_28 <= _GEN_9736;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_27 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h1b == rob_head) begin // @[rob.scala 476:25]
        rob_val_27 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_27 <= _GEN_9732;
      end
    end else begin
      rob_val_27 <= _GEN_9732;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_26 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h1a == rob_head) begin // @[rob.scala 476:25]
        rob_val_26 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_26 <= _GEN_9728;
      end
    end else begin
      rob_val_26 <= _GEN_9728;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_25 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h19 == rob_head) begin // @[rob.scala 476:25]
        rob_val_25 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_25 <= _GEN_9724;
      end
    end else begin
      rob_val_25 <= _GEN_9724;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_24 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h18 == rob_head) begin // @[rob.scala 476:25]
        rob_val_24 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_24 <= _GEN_9720;
      end
    end else begin
      rob_val_24 <= _GEN_9720;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_23 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h17 == rob_head) begin // @[rob.scala 476:25]
        rob_val_23 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_23 <= _GEN_9716;
      end
    end else begin
      rob_val_23 <= _GEN_9716;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_22 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h16 == rob_head) begin // @[rob.scala 476:25]
        rob_val_22 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_22 <= _GEN_9712;
      end
    end else begin
      rob_val_22 <= _GEN_9712;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_21 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h15 == rob_head) begin // @[rob.scala 476:25]
        rob_val_21 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_21 <= _GEN_9708;
      end
    end else begin
      rob_val_21 <= _GEN_9708;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_20 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h14 == rob_head) begin // @[rob.scala 476:25]
        rob_val_20 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_20 <= _GEN_9704;
      end
    end else begin
      rob_val_20 <= _GEN_9704;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_19 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h13 == rob_head) begin // @[rob.scala 476:25]
        rob_val_19 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_19 <= _GEN_9700;
      end
    end else begin
      rob_val_19 <= _GEN_9700;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_18 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h12 == rob_head) begin // @[rob.scala 476:25]
        rob_val_18 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_18 <= _GEN_9696;
      end
    end else begin
      rob_val_18 <= _GEN_9696;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_17 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h11 == rob_head) begin // @[rob.scala 476:25]
        rob_val_17 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_17 <= _GEN_9692;
      end
    end else begin
      rob_val_17 <= _GEN_9692;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_16 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h10 == rob_head) begin // @[rob.scala 476:25]
        rob_val_16 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_16 <= _GEN_9688;
      end
    end else begin
      rob_val_16 <= _GEN_9688;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_15 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'hf == rob_head) begin // @[rob.scala 476:25]
        rob_val_15 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_15 <= _GEN_9684;
      end
    end else begin
      rob_val_15 <= _GEN_9684;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_14 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'he == rob_head) begin // @[rob.scala 476:25]
        rob_val_14 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_14 <= _GEN_9680;
      end
    end else begin
      rob_val_14 <= _GEN_9680;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_13 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'hd == rob_head) begin // @[rob.scala 476:25]
        rob_val_13 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_13 <= _GEN_9676;
      end
    end else begin
      rob_val_13 <= _GEN_9676;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_12 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'hc == rob_head) begin // @[rob.scala 476:25]
        rob_val_12 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_12 <= _GEN_9672;
      end
    end else begin
      rob_val_12 <= _GEN_9672;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_11 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'hb == rob_head) begin // @[rob.scala 476:25]
        rob_val_11 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_11 <= _GEN_9668;
      end
    end else begin
      rob_val_11 <= _GEN_9668;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_10 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'ha == rob_head) begin // @[rob.scala 476:25]
        rob_val_10 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_10 <= _GEN_9664;
      end
    end else begin
      rob_val_10 <= _GEN_9664;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_9 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h9 == rob_head) begin // @[rob.scala 476:25]
        rob_val_9 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_9 <= _GEN_9660;
      end
    end else begin
      rob_val_9 <= _GEN_9660;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_8 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h8 == rob_head) begin // @[rob.scala 476:25]
        rob_val_8 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_8 <= _GEN_9656;
      end
    end else begin
      rob_val_8 <= _GEN_9656;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_7 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h7 == rob_head) begin // @[rob.scala 476:25]
        rob_val_7 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_7 <= _GEN_9652;
      end
    end else begin
      rob_val_7 <= _GEN_9652;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_6 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h6 == rob_head) begin // @[rob.scala 476:25]
        rob_val_6 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_6 <= _GEN_9648;
      end
    end else begin
      rob_val_6 <= _GEN_9648;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_5 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h5 == rob_head) begin // @[rob.scala 476:25]
        rob_val_5 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_5 <= _GEN_9644;
      end
    end else begin
      rob_val_5 <= _GEN_9644;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_4 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h4 == rob_head) begin // @[rob.scala 476:25]
        rob_val_4 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_4 <= _GEN_9640;
      end
    end else begin
      rob_val_4 <= _GEN_9640;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_3 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h3 == rob_head) begin // @[rob.scala 476:25]
        rob_val_3 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_3 <= _GEN_9636;
      end
    end else begin
      rob_val_3 <= _GEN_9636;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_2 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h2 == rob_head) begin // @[rob.scala 476:25]
        rob_val_2 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_2 <= _GEN_9632;
      end
    end else begin
      rob_val_2 <= _GEN_9632;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_1 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h1 == rob_head) begin // @[rob.scala 476:25]
        rob_val_1 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_1 <= _GEN_9628;
      end
    end else begin
      rob_val_1 <= _GEN_9628;
    end
    if (reset) begin // @[rob.scala 307:32]
      rob_val_0 <= 1'h0; // @[rob.scala 307:32]
    end else if (will_commit_0) begin // @[rob.scala 475:27]
      if (5'h0 == rob_head) begin // @[rob.scala 476:25]
        rob_val_0 <= 1'h0; // @[rob.scala 476:25]
      end else begin
        rob_val_0 <= _GEN_9624;
      end
    end else begin
      rob_val_0 <= _GEN_9624;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h1f == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_31 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_31 <= _GEN_6410;
      end
    end else begin
      rob_bsy_31 <= _GEN_6410;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h1e == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_30 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_30 <= _GEN_6409;
      end
    end else begin
      rob_bsy_30 <= _GEN_6409;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h1d == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_29 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_29 <= _GEN_6408;
      end
    end else begin
      rob_bsy_29 <= _GEN_6408;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h1c == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_28 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_28 <= _GEN_6407;
      end
    end else begin
      rob_bsy_28 <= _GEN_6407;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h1b == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_27 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_27 <= _GEN_6406;
      end
    end else begin
      rob_bsy_27 <= _GEN_6406;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h1a == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_26 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_26 <= _GEN_6405;
      end
    end else begin
      rob_bsy_26 <= _GEN_6405;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h19 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_25 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_25 <= _GEN_6404;
      end
    end else begin
      rob_bsy_25 <= _GEN_6404;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h18 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_24 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_24 <= _GEN_6403;
      end
    end else begin
      rob_bsy_24 <= _GEN_6403;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h17 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_23 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_23 <= _GEN_6402;
      end
    end else begin
      rob_bsy_23 <= _GEN_6402;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h16 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_22 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_22 <= _GEN_6401;
      end
    end else begin
      rob_bsy_22 <= _GEN_6401;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h15 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_21 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_21 <= _GEN_6400;
      end
    end else begin
      rob_bsy_21 <= _GEN_6400;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h14 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_20 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_20 <= _GEN_6399;
      end
    end else begin
      rob_bsy_20 <= _GEN_6399;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h13 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_19 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_19 <= _GEN_6398;
      end
    end else begin
      rob_bsy_19 <= _GEN_6398;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h12 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_18 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_18 <= _GEN_6397;
      end
    end else begin
      rob_bsy_18 <= _GEN_6397;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h11 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_17 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_17 <= _GEN_6396;
      end
    end else begin
      rob_bsy_17 <= _GEN_6396;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h10 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_16 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_16 <= _GEN_6395;
      end
    end else begin
      rob_bsy_16 <= _GEN_6395;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'hf == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_15 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_15 <= _GEN_6394;
      end
    end else begin
      rob_bsy_15 <= _GEN_6394;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'he == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_14 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_14 <= _GEN_6393;
      end
    end else begin
      rob_bsy_14 <= _GEN_6393;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'hd == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_13 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_13 <= _GEN_6392;
      end
    end else begin
      rob_bsy_13 <= _GEN_6392;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'hc == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_12 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_12 <= _GEN_6391;
      end
    end else begin
      rob_bsy_12 <= _GEN_6391;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'hb == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_11 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_11 <= _GEN_6390;
      end
    end else begin
      rob_bsy_11 <= _GEN_6390;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'ha == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_10 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_10 <= _GEN_6389;
      end
    end else begin
      rob_bsy_10 <= _GEN_6389;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h9 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_9 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_9 <= _GEN_6388;
      end
    end else begin
      rob_bsy_9 <= _GEN_6388;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h8 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_8 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_8 <= _GEN_6387;
      end
    end else begin
      rob_bsy_8 <= _GEN_6387;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h7 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_7 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_7 <= _GEN_6386;
      end
    end else begin
      rob_bsy_7 <= _GEN_6386;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h6 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_6 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_6 <= _GEN_6385;
      end
    end else begin
      rob_bsy_6 <= _GEN_6385;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h5 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_5 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_5 <= _GEN_6384;
      end
    end else begin
      rob_bsy_5 <= _GEN_6384;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h4 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_4 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_4 <= _GEN_6383;
      end
    end else begin
      rob_bsy_4 <= _GEN_6383;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h3 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_3 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_3 <= _GEN_6382;
      end
    end else begin
      rob_bsy_3 <= _GEN_6382;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h2 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_2 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_2 <= _GEN_6381;
      end
    end else begin
      rob_bsy_2 <= _GEN_6381;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h1 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_1 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_1 <= _GEN_6380;
      end
    end else begin
      rob_bsy_1 <= _GEN_6380;
    end
    if (io_lsu_clr_bsy_1_valid) begin // @[rob.scala 361:75]
      if (5'h0 == io_lsu_clr_bsy_1_bits) begin // @[rob.scala 363:26]
        rob_bsy_0 <= 1'h0; // @[rob.scala 363:26]
      end else begin
        rob_bsy_0 <= _GEN_6379;
      end
    end else begin
      rob_bsy_0 <= _GEN_6379;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h1f == com_idx) begin // @[rob.scala 435:30]
        rob_exception_31 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_31 <= _GEN_6804;
      end
    end else begin
      rob_exception_31 <= _GEN_6804;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h1e == com_idx) begin // @[rob.scala 435:30]
        rob_exception_30 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_30 <= _GEN_6803;
      end
    end else begin
      rob_exception_30 <= _GEN_6803;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h1d == com_idx) begin // @[rob.scala 435:30]
        rob_exception_29 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_29 <= _GEN_6802;
      end
    end else begin
      rob_exception_29 <= _GEN_6802;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h1c == com_idx) begin // @[rob.scala 435:30]
        rob_exception_28 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_28 <= _GEN_6801;
      end
    end else begin
      rob_exception_28 <= _GEN_6801;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h1b == com_idx) begin // @[rob.scala 435:30]
        rob_exception_27 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_27 <= _GEN_6800;
      end
    end else begin
      rob_exception_27 <= _GEN_6800;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h1a == com_idx) begin // @[rob.scala 435:30]
        rob_exception_26 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_26 <= _GEN_6799;
      end
    end else begin
      rob_exception_26 <= _GEN_6799;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h19 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_25 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_25 <= _GEN_6798;
      end
    end else begin
      rob_exception_25 <= _GEN_6798;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h18 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_24 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_24 <= _GEN_6797;
      end
    end else begin
      rob_exception_24 <= _GEN_6797;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h17 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_23 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_23 <= _GEN_6796;
      end
    end else begin
      rob_exception_23 <= _GEN_6796;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h16 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_22 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_22 <= _GEN_6795;
      end
    end else begin
      rob_exception_22 <= _GEN_6795;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h15 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_21 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_21 <= _GEN_6794;
      end
    end else begin
      rob_exception_21 <= _GEN_6794;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h14 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_20 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_20 <= _GEN_6793;
      end
    end else begin
      rob_exception_20 <= _GEN_6793;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h13 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_19 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_19 <= _GEN_6792;
      end
    end else begin
      rob_exception_19 <= _GEN_6792;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h12 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_18 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_18 <= _GEN_6791;
      end
    end else begin
      rob_exception_18 <= _GEN_6791;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h11 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_17 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_17 <= _GEN_6790;
      end
    end else begin
      rob_exception_17 <= _GEN_6790;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h10 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_16 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_16 <= _GEN_6789;
      end
    end else begin
      rob_exception_16 <= _GEN_6789;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'hf == com_idx) begin // @[rob.scala 435:30]
        rob_exception_15 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_15 <= _GEN_6788;
      end
    end else begin
      rob_exception_15 <= _GEN_6788;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'he == com_idx) begin // @[rob.scala 435:30]
        rob_exception_14 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_14 <= _GEN_6787;
      end
    end else begin
      rob_exception_14 <= _GEN_6787;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'hd == com_idx) begin // @[rob.scala 435:30]
        rob_exception_13 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_13 <= _GEN_6786;
      end
    end else begin
      rob_exception_13 <= _GEN_6786;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'hc == com_idx) begin // @[rob.scala 435:30]
        rob_exception_12 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_12 <= _GEN_6785;
      end
    end else begin
      rob_exception_12 <= _GEN_6785;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'hb == com_idx) begin // @[rob.scala 435:30]
        rob_exception_11 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_11 <= _GEN_6784;
      end
    end else begin
      rob_exception_11 <= _GEN_6784;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'ha == com_idx) begin // @[rob.scala 435:30]
        rob_exception_10 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_10 <= _GEN_6783;
      end
    end else begin
      rob_exception_10 <= _GEN_6783;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h9 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_9 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_9 <= _GEN_6782;
      end
    end else begin
      rob_exception_9 <= _GEN_6782;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h8 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_8 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_8 <= _GEN_6781;
      end
    end else begin
      rob_exception_8 <= _GEN_6781;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h7 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_7 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_7 <= _GEN_6780;
      end
    end else begin
      rob_exception_7 <= _GEN_6780;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h6 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_6 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_6 <= _GEN_6779;
      end
    end else begin
      rob_exception_6 <= _GEN_6779;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h5 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_5 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_5 <= _GEN_6778;
      end
    end else begin
      rob_exception_5 <= _GEN_6778;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h4 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_4 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_4 <= _GEN_6777;
      end
    end else begin
      rob_exception_4 <= _GEN_6777;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h3 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_3 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_3 <= _GEN_6776;
      end
    end else begin
      rob_exception_3 <= _GEN_6776;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h2 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_2 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_2 <= _GEN_6775;
      end
    end else begin
      rob_exception_2 <= _GEN_6775;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h1 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_1 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_1 <= _GEN_6774;
      end
    end else begin
      rob_exception_1 <= _GEN_6774;
    end
    if (rbk_row) begin // @[rob.scala 433:20]
      if (5'h0 == com_idx) begin // @[rob.scala 435:30]
        rob_exception_0 <= 1'h0; // @[rob.scala 435:30]
      end else begin
        rob_exception_0 <= _GEN_6773;
      end
    end else begin
      rob_exception_0 <= _GEN_6773;
    end
    _T_404 <= can_throw_exception_0 & _T_415; // @[rob.scala 545:52]
    _T_407 <= _T_406; // @[rob.scala 540:123]
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h0 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_0 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_0 <= _GEN_6603;
      end
    end else begin
      rob_unsafe_0 <= _GEN_6603;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h1 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_1 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_1 <= _GEN_6604;
      end
    end else begin
      rob_unsafe_1 <= _GEN_6604;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h2 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_2 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_2 <= _GEN_6605;
      end
    end else begin
      rob_unsafe_2 <= _GEN_6605;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h3 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_3 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_3 <= _GEN_6606;
      end
    end else begin
      rob_unsafe_3 <= _GEN_6606;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h4 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_4 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_4 <= _GEN_6607;
      end
    end else begin
      rob_unsafe_4 <= _GEN_6607;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h5 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_5 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_5 <= _GEN_6608;
      end
    end else begin
      rob_unsafe_5 <= _GEN_6608;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h6 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_6 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_6 <= _GEN_6609;
      end
    end else begin
      rob_unsafe_6 <= _GEN_6609;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h7 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_7 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_7 <= _GEN_6610;
      end
    end else begin
      rob_unsafe_7 <= _GEN_6610;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h8 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_8 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_8 <= _GEN_6611;
      end
    end else begin
      rob_unsafe_8 <= _GEN_6611;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h9 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_9 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_9 <= _GEN_6612;
      end
    end else begin
      rob_unsafe_9 <= _GEN_6612;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'ha == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_10 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_10 <= _GEN_6613;
      end
    end else begin
      rob_unsafe_10 <= _GEN_6613;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'hb == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_11 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_11 <= _GEN_6614;
      end
    end else begin
      rob_unsafe_11 <= _GEN_6614;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'hc == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_12 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_12 <= _GEN_6615;
      end
    end else begin
      rob_unsafe_12 <= _GEN_6615;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'hd == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_13 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_13 <= _GEN_6616;
      end
    end else begin
      rob_unsafe_13 <= _GEN_6616;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'he == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_14 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_14 <= _GEN_6617;
      end
    end else begin
      rob_unsafe_14 <= _GEN_6617;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'hf == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_15 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_15 <= _GEN_6618;
      end
    end else begin
      rob_unsafe_15 <= _GEN_6618;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h10 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_16 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_16 <= _GEN_6619;
      end
    end else begin
      rob_unsafe_16 <= _GEN_6619;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h11 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_17 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_17 <= _GEN_6620;
      end
    end else begin
      rob_unsafe_17 <= _GEN_6620;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h12 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_18 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_18 <= _GEN_6621;
      end
    end else begin
      rob_unsafe_18 <= _GEN_6621;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h13 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_19 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_19 <= _GEN_6622;
      end
    end else begin
      rob_unsafe_19 <= _GEN_6622;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h14 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_20 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_20 <= _GEN_6623;
      end
    end else begin
      rob_unsafe_20 <= _GEN_6623;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h15 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_21 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_21 <= _GEN_6624;
      end
    end else begin
      rob_unsafe_21 <= _GEN_6624;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h16 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_22 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_22 <= _GEN_6625;
      end
    end else begin
      rob_unsafe_22 <= _GEN_6625;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h17 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_23 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_23 <= _GEN_6626;
      end
    end else begin
      rob_unsafe_23 <= _GEN_6626;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h18 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_24 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_24 <= _GEN_6627;
      end
    end else begin
      rob_unsafe_24 <= _GEN_6627;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h19 == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_25 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_25 <= _GEN_6628;
      end
    end else begin
      rob_unsafe_25 <= _GEN_6628;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h1a == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_26 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_26 <= _GEN_6629;
      end
    end else begin
      rob_unsafe_26 <= _GEN_6629;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h1b == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_27 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_27 <= _GEN_6630;
      end
    end else begin
      rob_unsafe_27 <= _GEN_6630;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h1c == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_28 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_28 <= _GEN_6631;
      end
    end else begin
      rob_unsafe_28 <= _GEN_6631;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h1d == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_29 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_29 <= _GEN_6632;
      end
    end else begin
      rob_unsafe_29 <= _GEN_6632;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h1e == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_30 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_30 <= _GEN_6633;
      end
    end else begin
      rob_unsafe_30 <= _GEN_6633;
    end
    if (io_lsu_clr_unsafe_0_valid) begin // @[rob.scala 370:59]
      if (5'h1f == io_lsu_clr_unsafe_0_bits) begin // @[rob.scala 372:26]
        rob_unsafe_31 <= 1'h0; // @[rob.scala 372:26]
      end else begin
        rob_unsafe_31 <= _GEN_6634;
      end
    end else begin
      rob_unsafe_31 <= _GEN_6634;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h0 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_0_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_0_debug_inst <= _GEN_9625;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h0 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_0_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_0_debug_inst <= _GEN_9625;
      end
    end else begin
      rob_uop_0_debug_inst <= _GEN_9625;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_92) begin // @[rob.scala 455:7]
      rob_uop_0_br_mask <= _GEN_4614;
    end else if (rob_val_0) begin // @[rob.scala 458:32]
      rob_uop_0_br_mask <= _T_94; // @[rob.scala 460:28]
    end else begin
      rob_uop_0_br_mask <= _GEN_4614;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h0 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_0_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_0_taken <= _GEN_4454;
      end
    end else begin
      rob_uop_0_taken <= _GEN_4454;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h0 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_0_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_0_debug_fsrc <= _GEN_2918;
      end
    end else begin
      rob_uop_0_debug_fsrc <= _GEN_2918;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h0 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_0_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h1 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_1_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_1_debug_inst <= _GEN_9629;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h1 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_1_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_1_debug_inst <= _GEN_9629;
      end
    end else begin
      rob_uop_1_debug_inst <= _GEN_9629;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_96) begin // @[rob.scala 455:7]
      rob_uop_1_br_mask <= _GEN_4615;
    end else if (rob_val_1) begin // @[rob.scala 458:32]
      rob_uop_1_br_mask <= _T_98; // @[rob.scala 460:28]
    end else begin
      rob_uop_1_br_mask <= _GEN_4615;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h1 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_1_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_1_taken <= _GEN_4455;
      end
    end else begin
      rob_uop_1_taken <= _GEN_4455;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h1 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_1_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_1_debug_fsrc <= _GEN_2919;
      end
    end else begin
      rob_uop_1_debug_fsrc <= _GEN_2919;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_1_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h2 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_2_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_2_debug_inst <= _GEN_9633;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h2 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_2_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_2_debug_inst <= _GEN_9633;
      end
    end else begin
      rob_uop_2_debug_inst <= _GEN_9633;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_100) begin // @[rob.scala 455:7]
      rob_uop_2_br_mask <= _GEN_4616;
    end else if (rob_val_2) begin // @[rob.scala 458:32]
      rob_uop_2_br_mask <= _T_102; // @[rob.scala 460:28]
    end else begin
      rob_uop_2_br_mask <= _GEN_4616;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h2 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_2_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_2_taken <= _GEN_4456;
      end
    end else begin
      rob_uop_2_taken <= _GEN_4456;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h2 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_2_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_2_debug_fsrc <= _GEN_2920;
      end
    end else begin
      rob_uop_2_debug_fsrc <= _GEN_2920;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h2 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_2_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h3 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_3_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_3_debug_inst <= _GEN_9637;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h3 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_3_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_3_debug_inst <= _GEN_9637;
      end
    end else begin
      rob_uop_3_debug_inst <= _GEN_9637;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_104) begin // @[rob.scala 455:7]
      rob_uop_3_br_mask <= _GEN_4617;
    end else if (rob_val_3) begin // @[rob.scala 458:32]
      rob_uop_3_br_mask <= _T_106; // @[rob.scala 460:28]
    end else begin
      rob_uop_3_br_mask <= _GEN_4617;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h3 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_3_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_3_taken <= _GEN_4457;
      end
    end else begin
      rob_uop_3_taken <= _GEN_4457;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h3 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_3_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_3_debug_fsrc <= _GEN_2921;
      end
    end else begin
      rob_uop_3_debug_fsrc <= _GEN_2921;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h3 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_3_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h4 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_4_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_4_debug_inst <= _GEN_9641;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h4 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_4_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_4_debug_inst <= _GEN_9641;
      end
    end else begin
      rob_uop_4_debug_inst <= _GEN_9641;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_108) begin // @[rob.scala 455:7]
      rob_uop_4_br_mask <= _GEN_4618;
    end else if (rob_val_4) begin // @[rob.scala 458:32]
      rob_uop_4_br_mask <= _T_110; // @[rob.scala 460:28]
    end else begin
      rob_uop_4_br_mask <= _GEN_4618;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h4 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_4_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_4_taken <= _GEN_4458;
      end
    end else begin
      rob_uop_4_taken <= _GEN_4458;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h4 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_4_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_4_debug_fsrc <= _GEN_2922;
      end
    end else begin
      rob_uop_4_debug_fsrc <= _GEN_2922;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h4 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_4_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h5 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_5_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_5_debug_inst <= _GEN_9645;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h5 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_5_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_5_debug_inst <= _GEN_9645;
      end
    end else begin
      rob_uop_5_debug_inst <= _GEN_9645;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_112) begin // @[rob.scala 455:7]
      rob_uop_5_br_mask <= _GEN_4619;
    end else if (rob_val_5) begin // @[rob.scala 458:32]
      rob_uop_5_br_mask <= _T_114; // @[rob.scala 460:28]
    end else begin
      rob_uop_5_br_mask <= _GEN_4619;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h5 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_5_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_5_taken <= _GEN_4459;
      end
    end else begin
      rob_uop_5_taken <= _GEN_4459;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h5 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_5_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_5_debug_fsrc <= _GEN_2923;
      end
    end else begin
      rob_uop_5_debug_fsrc <= _GEN_2923;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h5 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_5_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h6 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_6_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_6_debug_inst <= _GEN_9649;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h6 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_6_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_6_debug_inst <= _GEN_9649;
      end
    end else begin
      rob_uop_6_debug_inst <= _GEN_9649;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_116) begin // @[rob.scala 455:7]
      rob_uop_6_br_mask <= _GEN_4620;
    end else if (rob_val_6) begin // @[rob.scala 458:32]
      rob_uop_6_br_mask <= _T_118; // @[rob.scala 460:28]
    end else begin
      rob_uop_6_br_mask <= _GEN_4620;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h6 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_6_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_6_taken <= _GEN_4460;
      end
    end else begin
      rob_uop_6_taken <= _GEN_4460;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h6 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_6_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_6_debug_fsrc <= _GEN_2924;
      end
    end else begin
      rob_uop_6_debug_fsrc <= _GEN_2924;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h6 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_6_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h7 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_7_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_7_debug_inst <= _GEN_9653;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h7 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_7_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_7_debug_inst <= _GEN_9653;
      end
    end else begin
      rob_uop_7_debug_inst <= _GEN_9653;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_120) begin // @[rob.scala 455:7]
      rob_uop_7_br_mask <= _GEN_4621;
    end else if (rob_val_7) begin // @[rob.scala 458:32]
      rob_uop_7_br_mask <= _T_122; // @[rob.scala 460:28]
    end else begin
      rob_uop_7_br_mask <= _GEN_4621;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h7 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_7_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_7_taken <= _GEN_4461;
      end
    end else begin
      rob_uop_7_taken <= _GEN_4461;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h7 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_7_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_7_debug_fsrc <= _GEN_2925;
      end
    end else begin
      rob_uop_7_debug_fsrc <= _GEN_2925;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h7 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_7_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h8 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_8_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_8_debug_inst <= _GEN_9657;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h8 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_8_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_8_debug_inst <= _GEN_9657;
      end
    end else begin
      rob_uop_8_debug_inst <= _GEN_9657;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_124) begin // @[rob.scala 455:7]
      rob_uop_8_br_mask <= _GEN_4622;
    end else if (rob_val_8) begin // @[rob.scala 458:32]
      rob_uop_8_br_mask <= _T_126; // @[rob.scala 460:28]
    end else begin
      rob_uop_8_br_mask <= _GEN_4622;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h8 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_8_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_8_taken <= _GEN_4462;
      end
    end else begin
      rob_uop_8_taken <= _GEN_4462;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h8 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_8_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_8_debug_fsrc <= _GEN_2926;
      end
    end else begin
      rob_uop_8_debug_fsrc <= _GEN_2926;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h8 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_8_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h9 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_9_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_9_debug_inst <= _GEN_9661;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h9 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_9_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_9_debug_inst <= _GEN_9661;
      end
    end else begin
      rob_uop_9_debug_inst <= _GEN_9661;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_128) begin // @[rob.scala 455:7]
      rob_uop_9_br_mask <= _GEN_4623;
    end else if (rob_val_9) begin // @[rob.scala 458:32]
      rob_uop_9_br_mask <= _T_130; // @[rob.scala 460:28]
    end else begin
      rob_uop_9_br_mask <= _GEN_4623;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h9 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_9_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_9_taken <= _GEN_4463;
      end
    end else begin
      rob_uop_9_taken <= _GEN_4463;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h9 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_9_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_9_debug_fsrc <= _GEN_2927;
      end
    end else begin
      rob_uop_9_debug_fsrc <= _GEN_2927;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h9 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_9_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'ha == rob_head) begin // @[rob.scala 498:36]
        rob_uop_10_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_10_debug_inst <= _GEN_9665;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'ha == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_10_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_10_debug_inst <= _GEN_9665;
      end
    end else begin
      rob_uop_10_debug_inst <= _GEN_9665;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_132) begin // @[rob.scala 455:7]
      rob_uop_10_br_mask <= _GEN_4624;
    end else if (rob_val_10) begin // @[rob.scala 458:32]
      rob_uop_10_br_mask <= _T_134; // @[rob.scala 460:28]
    end else begin
      rob_uop_10_br_mask <= _GEN_4624;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'ha == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_10_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_10_taken <= _GEN_4464;
      end
    end else begin
      rob_uop_10_taken <= _GEN_4464;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'ha == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_10_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_10_debug_fsrc <= _GEN_2928;
      end
    end else begin
      rob_uop_10_debug_fsrc <= _GEN_2928;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'ha == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_10_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'hb == rob_head) begin // @[rob.scala 498:36]
        rob_uop_11_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_11_debug_inst <= _GEN_9669;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'hb == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_11_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_11_debug_inst <= _GEN_9669;
      end
    end else begin
      rob_uop_11_debug_inst <= _GEN_9669;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_136) begin // @[rob.scala 455:7]
      rob_uop_11_br_mask <= _GEN_4625;
    end else if (rob_val_11) begin // @[rob.scala 458:32]
      rob_uop_11_br_mask <= _T_138; // @[rob.scala 460:28]
    end else begin
      rob_uop_11_br_mask <= _GEN_4625;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'hb == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_11_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_11_taken <= _GEN_4465;
      end
    end else begin
      rob_uop_11_taken <= _GEN_4465;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'hb == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_11_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_11_debug_fsrc <= _GEN_2929;
      end
    end else begin
      rob_uop_11_debug_fsrc <= _GEN_2929;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hb == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_11_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'hc == rob_head) begin // @[rob.scala 498:36]
        rob_uop_12_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_12_debug_inst <= _GEN_9673;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'hc == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_12_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_12_debug_inst <= _GEN_9673;
      end
    end else begin
      rob_uop_12_debug_inst <= _GEN_9673;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_140) begin // @[rob.scala 455:7]
      rob_uop_12_br_mask <= _GEN_4626;
    end else if (rob_val_12) begin // @[rob.scala 458:32]
      rob_uop_12_br_mask <= _T_142; // @[rob.scala 460:28]
    end else begin
      rob_uop_12_br_mask <= _GEN_4626;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'hc == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_12_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_12_taken <= _GEN_4466;
      end
    end else begin
      rob_uop_12_taken <= _GEN_4466;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'hc == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_12_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_12_debug_fsrc <= _GEN_2930;
      end
    end else begin
      rob_uop_12_debug_fsrc <= _GEN_2930;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hc == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_12_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'hd == rob_head) begin // @[rob.scala 498:36]
        rob_uop_13_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_13_debug_inst <= _GEN_9677;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'hd == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_13_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_13_debug_inst <= _GEN_9677;
      end
    end else begin
      rob_uop_13_debug_inst <= _GEN_9677;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_144) begin // @[rob.scala 455:7]
      rob_uop_13_br_mask <= _GEN_4627;
    end else if (rob_val_13) begin // @[rob.scala 458:32]
      rob_uop_13_br_mask <= _T_146; // @[rob.scala 460:28]
    end else begin
      rob_uop_13_br_mask <= _GEN_4627;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'hd == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_13_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_13_taken <= _GEN_4467;
      end
    end else begin
      rob_uop_13_taken <= _GEN_4467;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'hd == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_13_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_13_debug_fsrc <= _GEN_2931;
      end
    end else begin
      rob_uop_13_debug_fsrc <= _GEN_2931;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hd == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_13_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'he == rob_head) begin // @[rob.scala 498:36]
        rob_uop_14_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_14_debug_inst <= _GEN_9681;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'he == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_14_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_14_debug_inst <= _GEN_9681;
      end
    end else begin
      rob_uop_14_debug_inst <= _GEN_9681;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_148) begin // @[rob.scala 455:7]
      rob_uop_14_br_mask <= _GEN_4628;
    end else if (rob_val_14) begin // @[rob.scala 458:32]
      rob_uop_14_br_mask <= _T_150; // @[rob.scala 460:28]
    end else begin
      rob_uop_14_br_mask <= _GEN_4628;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'he == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_14_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_14_taken <= _GEN_4468;
      end
    end else begin
      rob_uop_14_taken <= _GEN_4468;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'he == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_14_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_14_debug_fsrc <= _GEN_2932;
      end
    end else begin
      rob_uop_14_debug_fsrc <= _GEN_2932;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'he == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_14_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'hf == rob_head) begin // @[rob.scala 498:36]
        rob_uop_15_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_15_debug_inst <= _GEN_9685;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'hf == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_15_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_15_debug_inst <= _GEN_9685;
      end
    end else begin
      rob_uop_15_debug_inst <= _GEN_9685;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_152) begin // @[rob.scala 455:7]
      rob_uop_15_br_mask <= _GEN_4629;
    end else if (rob_val_15) begin // @[rob.scala 458:32]
      rob_uop_15_br_mask <= _T_154; // @[rob.scala 460:28]
    end else begin
      rob_uop_15_br_mask <= _GEN_4629;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'hf == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_15_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_15_taken <= _GEN_4469;
      end
    end else begin
      rob_uop_15_taken <= _GEN_4469;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'hf == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_15_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_15_debug_fsrc <= _GEN_2933;
      end
    end else begin
      rob_uop_15_debug_fsrc <= _GEN_2933;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'hf == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_15_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h10 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_16_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_16_debug_inst <= _GEN_9689;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h10 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_16_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_16_debug_inst <= _GEN_9689;
      end
    end else begin
      rob_uop_16_debug_inst <= _GEN_9689;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_156) begin // @[rob.scala 455:7]
      rob_uop_16_br_mask <= _GEN_4630;
    end else if (rob_val_16) begin // @[rob.scala 458:32]
      rob_uop_16_br_mask <= _T_158; // @[rob.scala 460:28]
    end else begin
      rob_uop_16_br_mask <= _GEN_4630;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h10 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_16_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_16_taken <= _GEN_4470;
      end
    end else begin
      rob_uop_16_taken <= _GEN_4470;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h10 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_16_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_16_debug_fsrc <= _GEN_2934;
      end
    end else begin
      rob_uop_16_debug_fsrc <= _GEN_2934;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h10 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_16_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h11 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_17_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_17_debug_inst <= _GEN_9693;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h11 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_17_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_17_debug_inst <= _GEN_9693;
      end
    end else begin
      rob_uop_17_debug_inst <= _GEN_9693;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_160) begin // @[rob.scala 455:7]
      rob_uop_17_br_mask <= _GEN_4631;
    end else if (rob_val_17) begin // @[rob.scala 458:32]
      rob_uop_17_br_mask <= _T_162; // @[rob.scala 460:28]
    end else begin
      rob_uop_17_br_mask <= _GEN_4631;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h11 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_17_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_17_taken <= _GEN_4471;
      end
    end else begin
      rob_uop_17_taken <= _GEN_4471;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h11 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_17_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_17_debug_fsrc <= _GEN_2935;
      end
    end else begin
      rob_uop_17_debug_fsrc <= _GEN_2935;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h11 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_17_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h12 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_18_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_18_debug_inst <= _GEN_9697;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h12 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_18_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_18_debug_inst <= _GEN_9697;
      end
    end else begin
      rob_uop_18_debug_inst <= _GEN_9697;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_164) begin // @[rob.scala 455:7]
      rob_uop_18_br_mask <= _GEN_4632;
    end else if (rob_val_18) begin // @[rob.scala 458:32]
      rob_uop_18_br_mask <= _T_166; // @[rob.scala 460:28]
    end else begin
      rob_uop_18_br_mask <= _GEN_4632;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h12 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_18_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_18_taken <= _GEN_4472;
      end
    end else begin
      rob_uop_18_taken <= _GEN_4472;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h12 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_18_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_18_debug_fsrc <= _GEN_2936;
      end
    end else begin
      rob_uop_18_debug_fsrc <= _GEN_2936;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h12 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_18_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h13 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_19_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_19_debug_inst <= _GEN_9701;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h13 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_19_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_19_debug_inst <= _GEN_9701;
      end
    end else begin
      rob_uop_19_debug_inst <= _GEN_9701;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_168) begin // @[rob.scala 455:7]
      rob_uop_19_br_mask <= _GEN_4633;
    end else if (rob_val_19) begin // @[rob.scala 458:32]
      rob_uop_19_br_mask <= _T_170; // @[rob.scala 460:28]
    end else begin
      rob_uop_19_br_mask <= _GEN_4633;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h13 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_19_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_19_taken <= _GEN_4473;
      end
    end else begin
      rob_uop_19_taken <= _GEN_4473;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h13 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_19_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_19_debug_fsrc <= _GEN_2937;
      end
    end else begin
      rob_uop_19_debug_fsrc <= _GEN_2937;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h13 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_19_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h14 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_20_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_20_debug_inst <= _GEN_9705;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h14 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_20_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_20_debug_inst <= _GEN_9705;
      end
    end else begin
      rob_uop_20_debug_inst <= _GEN_9705;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_172) begin // @[rob.scala 455:7]
      rob_uop_20_br_mask <= _GEN_4634;
    end else if (rob_val_20) begin // @[rob.scala 458:32]
      rob_uop_20_br_mask <= _T_174; // @[rob.scala 460:28]
    end else begin
      rob_uop_20_br_mask <= _GEN_4634;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h14 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_20_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_20_taken <= _GEN_4474;
      end
    end else begin
      rob_uop_20_taken <= _GEN_4474;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h14 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_20_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_20_debug_fsrc <= _GEN_2938;
      end
    end else begin
      rob_uop_20_debug_fsrc <= _GEN_2938;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h14 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_20_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h15 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_21_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_21_debug_inst <= _GEN_9709;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h15 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_21_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_21_debug_inst <= _GEN_9709;
      end
    end else begin
      rob_uop_21_debug_inst <= _GEN_9709;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_176) begin // @[rob.scala 455:7]
      rob_uop_21_br_mask <= _GEN_4635;
    end else if (rob_val_21) begin // @[rob.scala 458:32]
      rob_uop_21_br_mask <= _T_178; // @[rob.scala 460:28]
    end else begin
      rob_uop_21_br_mask <= _GEN_4635;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h15 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_21_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_21_taken <= _GEN_4475;
      end
    end else begin
      rob_uop_21_taken <= _GEN_4475;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h15 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_21_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_21_debug_fsrc <= _GEN_2939;
      end
    end else begin
      rob_uop_21_debug_fsrc <= _GEN_2939;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h15 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_21_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h16 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_22_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_22_debug_inst <= _GEN_9713;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h16 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_22_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_22_debug_inst <= _GEN_9713;
      end
    end else begin
      rob_uop_22_debug_inst <= _GEN_9713;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_180) begin // @[rob.scala 455:7]
      rob_uop_22_br_mask <= _GEN_4636;
    end else if (rob_val_22) begin // @[rob.scala 458:32]
      rob_uop_22_br_mask <= _T_182; // @[rob.scala 460:28]
    end else begin
      rob_uop_22_br_mask <= _GEN_4636;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h16 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_22_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_22_taken <= _GEN_4476;
      end
    end else begin
      rob_uop_22_taken <= _GEN_4476;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h16 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_22_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_22_debug_fsrc <= _GEN_2940;
      end
    end else begin
      rob_uop_22_debug_fsrc <= _GEN_2940;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h16 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_22_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h17 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_23_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_23_debug_inst <= _GEN_9717;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h17 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_23_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_23_debug_inst <= _GEN_9717;
      end
    end else begin
      rob_uop_23_debug_inst <= _GEN_9717;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_184) begin // @[rob.scala 455:7]
      rob_uop_23_br_mask <= _GEN_4637;
    end else if (rob_val_23) begin // @[rob.scala 458:32]
      rob_uop_23_br_mask <= _T_186; // @[rob.scala 460:28]
    end else begin
      rob_uop_23_br_mask <= _GEN_4637;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h17 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_23_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_23_taken <= _GEN_4477;
      end
    end else begin
      rob_uop_23_taken <= _GEN_4477;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h17 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_23_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_23_debug_fsrc <= _GEN_2941;
      end
    end else begin
      rob_uop_23_debug_fsrc <= _GEN_2941;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h17 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_23_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h18 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_24_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_24_debug_inst <= _GEN_9721;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h18 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_24_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_24_debug_inst <= _GEN_9721;
      end
    end else begin
      rob_uop_24_debug_inst <= _GEN_9721;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_188) begin // @[rob.scala 455:7]
      rob_uop_24_br_mask <= _GEN_4638;
    end else if (rob_val_24) begin // @[rob.scala 458:32]
      rob_uop_24_br_mask <= _T_190; // @[rob.scala 460:28]
    end else begin
      rob_uop_24_br_mask <= _GEN_4638;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h18 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_24_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_24_taken <= _GEN_4478;
      end
    end else begin
      rob_uop_24_taken <= _GEN_4478;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h18 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_24_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_24_debug_fsrc <= _GEN_2942;
      end
    end else begin
      rob_uop_24_debug_fsrc <= _GEN_2942;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h18 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_24_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h19 == rob_head) begin // @[rob.scala 498:36]
        rob_uop_25_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_25_debug_inst <= _GEN_9725;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h19 == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_25_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_25_debug_inst <= _GEN_9725;
      end
    end else begin
      rob_uop_25_debug_inst <= _GEN_9725;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_192) begin // @[rob.scala 455:7]
      rob_uop_25_br_mask <= _GEN_4639;
    end else if (rob_val_25) begin // @[rob.scala 458:32]
      rob_uop_25_br_mask <= _T_194; // @[rob.scala 460:28]
    end else begin
      rob_uop_25_br_mask <= _GEN_4639;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h19 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_25_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_25_taken <= _GEN_4479;
      end
    end else begin
      rob_uop_25_taken <= _GEN_4479;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h19 == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_25_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_25_debug_fsrc <= _GEN_2943;
      end
    end else begin
      rob_uop_25_debug_fsrc <= _GEN_2943;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h19 == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_25_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h1a == rob_head) begin // @[rob.scala 498:36]
        rob_uop_26_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_26_debug_inst <= _GEN_9729;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h1a == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_26_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_26_debug_inst <= _GEN_9729;
      end
    end else begin
      rob_uop_26_debug_inst <= _GEN_9729;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_196) begin // @[rob.scala 455:7]
      rob_uop_26_br_mask <= _GEN_4640;
    end else if (rob_val_26) begin // @[rob.scala 458:32]
      rob_uop_26_br_mask <= _T_198; // @[rob.scala 460:28]
    end else begin
      rob_uop_26_br_mask <= _GEN_4640;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h1a == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_26_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_26_taken <= _GEN_4480;
      end
    end else begin
      rob_uop_26_taken <= _GEN_4480;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h1a == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_26_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_26_debug_fsrc <= _GEN_2944;
      end
    end else begin
      rob_uop_26_debug_fsrc <= _GEN_2944;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1a == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_26_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h1b == rob_head) begin // @[rob.scala 498:36]
        rob_uop_27_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_27_debug_inst <= _GEN_9733;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h1b == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_27_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_27_debug_inst <= _GEN_9733;
      end
    end else begin
      rob_uop_27_debug_inst <= _GEN_9733;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_200) begin // @[rob.scala 455:7]
      rob_uop_27_br_mask <= _GEN_4641;
    end else if (rob_val_27) begin // @[rob.scala 458:32]
      rob_uop_27_br_mask <= _T_202; // @[rob.scala 460:28]
    end else begin
      rob_uop_27_br_mask <= _GEN_4641;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h1b == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_27_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_27_taken <= _GEN_4481;
      end
    end else begin
      rob_uop_27_taken <= _GEN_4481;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h1b == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_27_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_27_debug_fsrc <= _GEN_2945;
      end
    end else begin
      rob_uop_27_debug_fsrc <= _GEN_2945;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1b == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_27_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h1c == rob_head) begin // @[rob.scala 498:36]
        rob_uop_28_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_28_debug_inst <= _GEN_9737;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h1c == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_28_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_28_debug_inst <= _GEN_9737;
      end
    end else begin
      rob_uop_28_debug_inst <= _GEN_9737;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_204) begin // @[rob.scala 455:7]
      rob_uop_28_br_mask <= _GEN_4642;
    end else if (rob_val_28) begin // @[rob.scala 458:32]
      rob_uop_28_br_mask <= _T_206; // @[rob.scala 460:28]
    end else begin
      rob_uop_28_br_mask <= _GEN_4642;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h1c == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_28_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_28_taken <= _GEN_4482;
      end
    end else begin
      rob_uop_28_taken <= _GEN_4482;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h1c == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_28_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_28_debug_fsrc <= _GEN_2946;
      end
    end else begin
      rob_uop_28_debug_fsrc <= _GEN_2946;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1c == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_28_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h1d == rob_head) begin // @[rob.scala 498:36]
        rob_uop_29_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_29_debug_inst <= _GEN_9741;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h1d == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_29_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_29_debug_inst <= _GEN_9741;
      end
    end else begin
      rob_uop_29_debug_inst <= _GEN_9741;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_208) begin // @[rob.scala 455:7]
      rob_uop_29_br_mask <= _GEN_4643;
    end else if (rob_val_29) begin // @[rob.scala 458:32]
      rob_uop_29_br_mask <= _T_210; // @[rob.scala 460:28]
    end else begin
      rob_uop_29_br_mask <= _GEN_4643;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h1d == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_29_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_29_taken <= _GEN_4483;
      end
    end else begin
      rob_uop_29_taken <= _GEN_4483;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h1d == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_29_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_29_debug_fsrc <= _GEN_2947;
      end
    end else begin
      rob_uop_29_debug_fsrc <= _GEN_2947;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1d == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_29_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h1e == rob_head) begin // @[rob.scala 498:36]
        rob_uop_30_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_30_debug_inst <= _GEN_9745;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h1e == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_30_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_30_debug_inst <= _GEN_9745;
      end
    end else begin
      rob_uop_30_debug_inst <= _GEN_9745;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_212) begin // @[rob.scala 455:7]
      rob_uop_30_br_mask <= _GEN_4644;
    end else if (rob_val_30) begin // @[rob.scala 458:32]
      rob_uop_30_br_mask <= _T_214; // @[rob.scala 460:28]
    end else begin
      rob_uop_30_br_mask <= _GEN_4644;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h1e == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_30_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_30_taken <= _GEN_4484;
      end
    end else begin
      rob_uop_30_taken <= _GEN_4484;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h1e == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_30_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_30_debug_fsrc <= _GEN_2948;
      end
    end else begin
      rob_uop_30_debug_fsrc <= _GEN_2948;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1e == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_30_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_uopc <= io_enq_uops_0_uopc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_inst <= io_enq_uops_0_inst; // @[rob.scala 328:31]
      end
    end
    if (will_commit_0) begin // @[rob.scala 497:27]
      if (5'h1f == rob_head) begin // @[rob.scala 498:36]
        rob_uop_31_debug_inst <= 32'h4033; // @[rob.scala 498:36]
      end else begin
        rob_uop_31_debug_inst <= _GEN_9749;
      end
    end else if (rbk_row) begin // @[rob.scala 500:5]
      if (5'h1f == rob_tail) begin // @[rob.scala 501:36]
        rob_uop_31_debug_inst <= 32'h4033; // @[rob.scala 501:36]
      end else begin
        rob_uop_31_debug_inst <= _GEN_9749;
      end
    end else begin
      rob_uop_31_debug_inst <= _GEN_9749;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_is_rvc <= io_enq_uops_0_is_rvc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_debug_pc <= io_enq_uops_0_debug_pc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_iq_type <= io_enq_uops_0_iq_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_fu_code <= io_enq_uops_0_fu_code; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_ctrl_br_type <= io_enq_uops_0_ctrl_br_type; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_ctrl_op1_sel <= io_enq_uops_0_ctrl_op1_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_ctrl_op2_sel <= io_enq_uops_0_ctrl_op2_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_ctrl_imm_sel <= io_enq_uops_0_ctrl_imm_sel; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_ctrl_op_fcn <= io_enq_uops_0_ctrl_op_fcn; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_ctrl_fcn_dw <= io_enq_uops_0_ctrl_fcn_dw; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_ctrl_csr_cmd <= io_enq_uops_0_ctrl_csr_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_ctrl_is_load <= io_enq_uops_0_ctrl_is_load; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_ctrl_is_sta <= io_enq_uops_0_ctrl_is_sta; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_ctrl_is_std <= io_enq_uops_0_ctrl_is_std; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_iw_state <= io_enq_uops_0_iw_state; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_iw_p1_poisoned <= io_enq_uops_0_iw_p1_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_iw_p2_poisoned <= io_enq_uops_0_iw_p2_poisoned; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_is_br <= io_enq_uops_0_is_br; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_is_jalr <= io_enq_uops_0_is_jalr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_is_jal <= io_enq_uops_0_is_jal; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_is_sfb <= io_enq_uops_0_is_sfb; // @[rob.scala 328:31]
      end
    end
    if (_T_216) begin // @[rob.scala 455:7]
      rob_uop_31_br_mask <= _GEN_4645;
    end else if (rob_val_31) begin // @[rob.scala 458:32]
      rob_uop_31_br_mask <= _T_218; // @[rob.scala 460:28]
    end else begin
      rob_uop_31_br_mask <= _GEN_4645;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_br_tag <= io_enq_uops_0_br_tag; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_ftq_idx <= io_enq_uops_0_ftq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_edge_inst <= io_enq_uops_0_edge_inst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_pc_lob <= io_enq_uops_0_pc_lob; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h1f == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 470:65]
        rob_uop_31_taken <= io_brupdate_b2_taken; // @[rob.scala 470:65]
      end else begin
        rob_uop_31_taken <= _GEN_4485;
      end
    end else begin
      rob_uop_31_taken <= _GEN_4485;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_imm_packed <= io_enq_uops_0_imm_packed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_csr_addr <= io_enq_uops_0_csr_addr; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_rob_idx <= io_enq_uops_0_rob_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_ldq_idx <= io_enq_uops_0_ldq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_stq_idx <= io_enq_uops_0_stq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_rxq_idx <= io_enq_uops_0_rxq_idx; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_pdst <= io_enq_uops_0_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_prs1 <= io_enq_uops_0_prs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_prs2 <= io_enq_uops_0_prs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_prs3 <= io_enq_uops_0_prs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_ppred <= io_enq_uops_0_ppred; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_prs1_busy <= io_enq_uops_0_prs1_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_prs2_busy <= io_enq_uops_0_prs2_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_prs3_busy <= io_enq_uops_0_prs3_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_ppred_busy <= io_enq_uops_0_ppred_busy; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_stale_pdst <= io_enq_uops_0_stale_pdst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_exception <= io_enq_uops_0_exception; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_exc_cause <= io_enq_uops_0_exc_cause; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_bypassable <= io_enq_uops_0_bypassable; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_mem_cmd <= io_enq_uops_0_mem_cmd; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_mem_size <= io_enq_uops_0_mem_size; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_mem_signed <= io_enq_uops_0_mem_signed; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_is_fence <= io_enq_uops_0_is_fence; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_is_fencei <= io_enq_uops_0_is_fencei; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_is_amo <= io_enq_uops_0_is_amo; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_uses_ldq <= io_enq_uops_0_uses_ldq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_uses_stq <= io_enq_uops_0_uses_stq; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_is_unique <= io_enq_uops_0_is_unique; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_flush_on_commit <= io_enq_uops_0_flush_on_commit; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_ldst_is_rs1 <= io_enq_uops_0_ldst_is_rs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_ldst <= io_enq_uops_0_ldst; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_lrs1 <= io_enq_uops_0_lrs1; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_lrs2 <= io_enq_uops_0_lrs2; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_lrs3 <= io_enq_uops_0_lrs3; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_ldst_val <= io_enq_uops_0_ldst_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_dst_rtype <= io_enq_uops_0_dst_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_lrs1_rtype <= io_enq_uops_0_lrs1_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_lrs2_rtype <= io_enq_uops_0_lrs2_rtype; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_frs3_en <= io_enq_uops_0_frs3_en; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_fp_val <= io_enq_uops_0_fp_val; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_fp_single <= io_enq_uops_0_fp_single; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_xcpt_pf_if <= io_enq_uops_0_xcpt_pf_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_xcpt_ae_if <= io_enq_uops_0_xcpt_ae_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_xcpt_ma_if <= io_enq_uops_0_xcpt_ma_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_bp_debug_if <= io_enq_uops_0_bp_debug_if; // @[rob.scala 328:31]
      end
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_bp_xcpt_if <= io_enq_uops_0_bp_xcpt_if; // @[rob.scala 328:31]
      end
    end
    if (io_brupdate_b2_mispredict) begin // @[rob.scala 468:58]
      if (5'h1f == io_brupdate_b2_uop_rob_idx) begin // @[rob.scala 469:65]
        rob_uop_31_debug_fsrc <= 2'h3; // @[rob.scala 469:65]
      end else begin
        rob_uop_31_debug_fsrc <= _GEN_2949;
      end
    end else begin
      rob_uop_31_debug_fsrc <= _GEN_2949;
    end
    if (io_enq_valids_0) begin // @[rob.scala 323:29]
      if (5'h1f == rob_tail) begin // @[rob.scala 328:31]
        rob_uop_31_debug_tsrc <= io_enq_uops_0_debug_tsrc; // @[rob.scala 328:31]
      end
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h0 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_0 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_0 <= _GEN_6027;
      end
    end else begin
      rob_predicated_0 <= _GEN_6027;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h1 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_1 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_1 <= _GEN_6028;
      end
    end else begin
      rob_predicated_1 <= _GEN_6028;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h2 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_2 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_2 <= _GEN_6029;
      end
    end else begin
      rob_predicated_2 <= _GEN_6029;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h3 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_3 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_3 <= _GEN_6030;
      end
    end else begin
      rob_predicated_3 <= _GEN_6030;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h4 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_4 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_4 <= _GEN_6031;
      end
    end else begin
      rob_predicated_4 <= _GEN_6031;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h5 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_5 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_5 <= _GEN_6032;
      end
    end else begin
      rob_predicated_5 <= _GEN_6032;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h6 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_6 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_6 <= _GEN_6033;
      end
    end else begin
      rob_predicated_6 <= _GEN_6033;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h7 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_7 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_7 <= _GEN_6034;
      end
    end else begin
      rob_predicated_7 <= _GEN_6034;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h8 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_8 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_8 <= _GEN_6035;
      end
    end else begin
      rob_predicated_8 <= _GEN_6035;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h9 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_9 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_9 <= _GEN_6036;
      end
    end else begin
      rob_predicated_9 <= _GEN_6036;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'ha == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_10 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_10 <= _GEN_6037;
      end
    end else begin
      rob_predicated_10 <= _GEN_6037;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'hb == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_11 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_11 <= _GEN_6038;
      end
    end else begin
      rob_predicated_11 <= _GEN_6038;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'hc == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_12 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_12 <= _GEN_6039;
      end
    end else begin
      rob_predicated_12 <= _GEN_6039;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'hd == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_13 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_13 <= _GEN_6040;
      end
    end else begin
      rob_predicated_13 <= _GEN_6040;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'he == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_14 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_14 <= _GEN_6041;
      end
    end else begin
      rob_predicated_14 <= _GEN_6041;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'hf == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_15 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_15 <= _GEN_6042;
      end
    end else begin
      rob_predicated_15 <= _GEN_6042;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h10 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_16 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_16 <= _GEN_6043;
      end
    end else begin
      rob_predicated_16 <= _GEN_6043;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h11 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_17 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_17 <= _GEN_6044;
      end
    end else begin
      rob_predicated_17 <= _GEN_6044;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h12 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_18 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_18 <= _GEN_6045;
      end
    end else begin
      rob_predicated_18 <= _GEN_6045;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h13 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_19 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_19 <= _GEN_6046;
      end
    end else begin
      rob_predicated_19 <= _GEN_6046;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h14 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_20 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_20 <= _GEN_6047;
      end
    end else begin
      rob_predicated_20 <= _GEN_6047;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h15 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_21 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_21 <= _GEN_6048;
      end
    end else begin
      rob_predicated_21 <= _GEN_6048;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h16 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_22 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_22 <= _GEN_6049;
      end
    end else begin
      rob_predicated_22 <= _GEN_6049;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h17 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_23 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_23 <= _GEN_6050;
      end
    end else begin
      rob_predicated_23 <= _GEN_6050;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h18 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_24 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_24 <= _GEN_6051;
      end
    end else begin
      rob_predicated_24 <= _GEN_6051;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h19 == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_25 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_25 <= _GEN_6052;
      end
    end else begin
      rob_predicated_25 <= _GEN_6052;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h1a == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_26 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_26 <= _GEN_6053;
      end
    end else begin
      rob_predicated_26 <= _GEN_6053;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h1b == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_27 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_27 <= _GEN_6054;
      end
    end else begin
      rob_predicated_27 <= _GEN_6054;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h1c == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_28 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_28 <= _GEN_6055;
      end
    end else begin
      rob_predicated_28 <= _GEN_6055;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h1d == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_29 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_29 <= _GEN_6056;
      end
    end else begin
      rob_predicated_29 <= _GEN_6056;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h1e == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_30 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_30 <= _GEN_6057;
      end
    end else begin
      rob_predicated_30 <= _GEN_6057;
    end
    if (io_wb_resps_3_valid) begin // @[rob.scala 346:69]
      if (5'h1f == io_wb_resps_3_bits_uop_rob_idx) begin // @[rob.scala 349:34]
        rob_predicated_31 <= io_wb_resps_3_bits_predicated; // @[rob.scala 349:34]
      end else begin
        rob_predicated_31 <= _GEN_6058;
      end
    end else begin
      rob_predicated_31 <= _GEN_6058;
    end
    _T_406 <= can_throw_exception_0 & _T_415; // @[rob.scala 545:52]
    if (reset) begin // @[rob.scala 677:30]
      r_partial_row <= 1'h0; // @[rob.scala 677:30]
    end else if (io_enq_valids_0) begin // @[rob.scala 679:36]
      r_partial_row <= io_enq_partial_stall; // @[rob.scala 680:19]
    end
    if (reset) begin // @[rob.scala 714:36]
      pnr_maybe_at_tail <= 1'h0; // @[rob.scala 714:36]
    end else begin
      pnr_maybe_at_tail <= ~rob_deq & (do_inc_row | pnr_maybe_at_tail); // @[rob.scala 736:23]
    end
    _T_609 <= can_throw_exception_0 & _T_415; // @[rob.scala 545:52]
    _T_610 <= _T_609; // @[rob.scala 808:22]
    _T_614 <= can_throw_exception_0 & _T_415; // @[rob.scala 545:52]
    _T_618 <= rob_head_uses_ldq_0 & _T_616; // @[rob.scala 865:98]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_enq_valids_0 & ~(~rob_tail_vals_0 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:333 assert (rob_val(rob_tail) === false.B, \"[rob] overwriting a valid entry.\")\n"
            ); // @[rob.scala 333:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_enq_valids_0 & ~(~rob_tail_vals_0 | reset)) begin
          $fatal; // @[rob.scala 333:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_enq_valids_0 & ~(io_enq_uops_0_rob_idx == rob_tail | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at rob.scala:334 assert ((io.enq_uops(w).rob_idx >> log2Ceil(coreWidth)) === rob_tail)\n"
            ); // @[rob.scala 334:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_enq_valids_0 & ~(io_enq_uops_0_rob_idx == rob_tail | reset)) begin
          $fatal; // @[rob.scala 334:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_lsu_clr_bsy_0_valid & ~(_GEN_6346 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n"
            ); // @[rob.scala 365:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_lsu_clr_bsy_0_valid & ~(_GEN_6346 | reset)) begin
          $fatal; // @[rob.scala 365:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_lsu_clr_bsy_0_valid & ~(_GEN_6378 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n"
            ); // @[rob.scala 366:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_lsu_clr_bsy_0_valid & ~(_GEN_6378 | reset)) begin
          $fatal; // @[rob.scala 366:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_lsu_clr_bsy_1_valid & ~(_GEN_6538 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n"
            ); // @[rob.scala 365:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_lsu_clr_bsy_1_valid & ~(_GEN_6538 | reset)) begin
          $fatal; // @[rob.scala 365:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_lsu_clr_bsy_1_valid & ~(_GEN_6570 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n"
            ); // @[rob.scala 366:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_lsu_clr_bsy_1_valid & ~(_GEN_6570 | reset)) begin
          $fatal; // @[rob.scala 366:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_lxcpt_valid & _T_65 & ~(_GEN_6772 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: An instruction marked as safe is causing an exception\n    at rob.scala:394 assert(rob_unsafe(GetRowIdx(io.lxcpt.bits.uop.rob_idx)),\n"
            ); // @[rob.scala 394:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_lxcpt_valid & _T_65 & ~(_GEN_6772 | reset)) begin
          $fatal; // @[rob.scala 394:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_commit_valids_0 & io_commit_rbk_valids_0) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: com_valids and rbk_valids are mutually exclusive\n    at rob.scala:430 assert (!(io.commit.valids.reduce(_||_) && io.commit.rbk_valids.reduce(_||_)),\n"
            ); // @[rob.scala 430:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_commit_valids_0 & io_commit_rbk_valids_0) | reset)) begin
          $fatal; // @[rob.scala 430:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_wb_resps_0_valid & _T_293) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 514:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_wb_resps_0_valid & _T_293) | reset)) begin
          $fatal; // @[rob.scala 514:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_wb_resps_0_valid & _T_301) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 517:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_wb_resps_0_valid & _T_301) | reset)) begin
          $fatal; // @[rob.scala 517:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~_T_311 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 520:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~_T_311 | reset)) begin
          $fatal; // @[rob.scala 520:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_wb_resps_1_valid & _T_321) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 514:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_wb_resps_1_valid & _T_321) | reset)) begin
          $fatal; // @[rob.scala 514:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_wb_resps_1_valid & _T_329) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 517:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_wb_resps_1_valid & _T_329) | reset)) begin
          $fatal; // @[rob.scala 517:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~_T_339 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 520:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~_T_339 | reset)) begin
          $fatal; // @[rob.scala 520:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_wb_resps_2_valid & _T_349) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 514:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_wb_resps_2_valid & _T_349) | reset)) begin
          $fatal; // @[rob.scala 514:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_wb_resps_2_valid & _T_357) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 517:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_wb_resps_2_valid & _T_357) | reset)) begin
          $fatal; // @[rob.scala 517:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~_T_367 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 520:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~_T_367 | reset)) begin
          $fatal; // @[rob.scala 520:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_wb_resps_3_valid & _T_377) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 514:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_wb_resps_3_valid & _T_377) | reset)) begin
          $fatal; // @[rob.scala 514:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_wb_resps_3_valid & _T_385) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 517:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_wb_resps_3_valid & _T_385) | reset)) begin
          $fatal; // @[rob.scala 517:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~_T_395 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 520:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~_T_395 | reset)) begin
          $fatal; // @[rob.scala 520:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~_T_447 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:607 assert (!(io.commit.valids(w) &&\n"
            ); // @[rob.scala 607:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~_T_447 | reset)) begin
          $fatal; // @[rob.scala 607:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~_T_456 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:611 assert (!(io.commit.valids(w) &&\n"
            ); // @[rob.scala 611:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~_T_456 | reset)) begin
          $fatal; // @[rob.scala 611:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(will_throw_exception & _T_466) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB trying to throw an exception, but it doesn't have a valid xcpt_cause\n    at rob.scala:658 assert (!(exception_thrown && !r_xcpt_val),\n"
            ); // @[rob.scala 658:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(will_throw_exception & _T_466) | reset)) begin
          $fatal; // @[rob.scala 658:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(empty & r_xcpt_val) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB is empty, but believes it has an outstanding exception.\n    at rob.scala:661 assert (!(empty && r_xcpt_val),\n"
            ); // @[rob.scala 661:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(empty & r_xcpt_val) | reset)) begin
          $fatal; // @[rob.scala 661:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(will_throw_exception & r_xcpt_uop_rob_idx != rob_head) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB is throwing an exception, but the stored exception information's rob_idx does not match the rob_head\n    at rob.scala:664 assert (!(will_throw_exception && (GetRowIdx(r_xcpt_uop.rob_idx) =/= rob_head)),\n"
            ); // @[rob.scala 664:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(will_throw_exception & r_xcpt_uop_rob_idx != rob_head) | reset)) begin
          $fatal; // @[rob.scala 664:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~_T_549 | rob_pnr == rob_tail | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at rob.scala:740 assert(!IsOlder(rob_pnr_idx, rob_head_idx, rob_tail_idx) || rob_pnr_idx === rob_tail_idx)\n"
            ); // @[rob.scala 740:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~_T_549 | rob_pnr == rob_tail | reset)) begin
          $fatal; // @[rob.scala 740:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~_T_560 | full | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at rob.scala:743 assert(!IsOlder(rob_tail_idx, rob_pnr_idx, rob_head_idx) || full)\n"
            ); // @[rob.scala 743:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~_T_560 | full | reset)) begin
          $fatal; // @[rob.scala 743:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    rob_debug_inst_mem_0[initvar] = _RAND_0[31:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    rob_fflags[initvar] = _RAND_3[4:0];
  _RAND_4 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    rob_debug_wdata[initvar] = _RAND_4[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rob_debug_inst_mem_0_rob_debug_inst_rdata_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  rob_debug_inst_mem_0_rob_debug_inst_rdata_addr_pipe_0 = _RAND_2[4:0];
  _RAND_5 = {1{`RANDOM}};
  rob_state = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  rob_head = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  rob_tail = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  rob_pnr = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  maybe_full = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  r_xcpt_val = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  r_xcpt_uop_br_mask = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  r_xcpt_uop_rob_idx = _RAND_12[4:0];
  _RAND_13 = {2{`RANDOM}};
  r_xcpt_uop_exc_cause = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  r_xcpt_badvaddr = _RAND_14[39:0];
  _RAND_15 = {1{`RANDOM}};
  rob_val_31 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  rob_val_30 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  rob_val_29 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  rob_val_28 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  rob_val_27 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  rob_val_26 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  rob_val_25 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  rob_val_24 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  rob_val_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  rob_val_22 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  rob_val_21 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  rob_val_20 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  rob_val_19 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  rob_val_18 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  rob_val_17 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  rob_val_16 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  rob_val_15 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  rob_val_14 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  rob_val_13 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  rob_val_12 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  rob_val_11 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  rob_val_10 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  rob_val_9 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  rob_val_8 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  rob_val_7 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  rob_val_6 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  rob_val_5 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  rob_val_4 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  rob_val_3 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  rob_val_2 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  rob_val_1 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  rob_val_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  rob_bsy_31 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  rob_bsy_30 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  rob_bsy_29 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  rob_bsy_28 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  rob_bsy_27 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  rob_bsy_26 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  rob_bsy_25 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  rob_bsy_24 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  rob_bsy_23 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  rob_bsy_22 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  rob_bsy_21 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  rob_bsy_20 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  rob_bsy_19 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  rob_bsy_18 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  rob_bsy_17 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  rob_bsy_16 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  rob_bsy_15 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  rob_bsy_14 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  rob_bsy_13 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  rob_bsy_12 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  rob_bsy_11 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  rob_bsy_10 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  rob_bsy_9 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  rob_bsy_8 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  rob_bsy_7 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  rob_bsy_6 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  rob_bsy_5 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  rob_bsy_4 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  rob_bsy_3 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  rob_bsy_2 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  rob_bsy_1 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  rob_bsy_0 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  rob_exception_31 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  rob_exception_30 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  rob_exception_29 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  rob_exception_28 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  rob_exception_27 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  rob_exception_26 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  rob_exception_25 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  rob_exception_24 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  rob_exception_23 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  rob_exception_22 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  rob_exception_21 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  rob_exception_20 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  rob_exception_19 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  rob_exception_18 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  rob_exception_17 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  rob_exception_16 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  rob_exception_15 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  rob_exception_14 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  rob_exception_13 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  rob_exception_12 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  rob_exception_11 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  rob_exception_10 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  rob_exception_9 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  rob_exception_8 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  rob_exception_7 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  rob_exception_6 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  rob_exception_5 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  rob_exception_4 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  rob_exception_3 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  rob_exception_2 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  rob_exception_1 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  rob_exception_0 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  _T_404 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  _T_407 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  rob_unsafe_0 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  rob_unsafe_1 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  rob_unsafe_2 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  rob_unsafe_3 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  rob_unsafe_4 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  rob_unsafe_5 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  rob_unsafe_6 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  rob_unsafe_7 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  rob_unsafe_8 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  rob_unsafe_9 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  rob_unsafe_10 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  rob_unsafe_11 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  rob_unsafe_12 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  rob_unsafe_13 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  rob_unsafe_14 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  rob_unsafe_15 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  rob_unsafe_16 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  rob_unsafe_17 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  rob_unsafe_18 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  rob_unsafe_19 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  rob_unsafe_20 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  rob_unsafe_21 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  rob_unsafe_22 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  rob_unsafe_23 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  rob_unsafe_24 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  rob_unsafe_25 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  rob_unsafe_26 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  rob_unsafe_27 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  rob_unsafe_28 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  rob_unsafe_29 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  rob_unsafe_30 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  rob_unsafe_31 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  rob_uop_0_uopc = _RAND_145[6:0];
  _RAND_146 = {1{`RANDOM}};
  rob_uop_0_inst = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  rob_uop_0_debug_inst = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  rob_uop_0_is_rvc = _RAND_148[0:0];
  _RAND_149 = {2{`RANDOM}};
  rob_uop_0_debug_pc = _RAND_149[39:0];
  _RAND_150 = {1{`RANDOM}};
  rob_uop_0_iq_type = _RAND_150[2:0];
  _RAND_151 = {1{`RANDOM}};
  rob_uop_0_fu_code = _RAND_151[9:0];
  _RAND_152 = {1{`RANDOM}};
  rob_uop_0_ctrl_br_type = _RAND_152[3:0];
  _RAND_153 = {1{`RANDOM}};
  rob_uop_0_ctrl_op1_sel = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  rob_uop_0_ctrl_op2_sel = _RAND_154[2:0];
  _RAND_155 = {1{`RANDOM}};
  rob_uop_0_ctrl_imm_sel = _RAND_155[2:0];
  _RAND_156 = {1{`RANDOM}};
  rob_uop_0_ctrl_op_fcn = _RAND_156[3:0];
  _RAND_157 = {1{`RANDOM}};
  rob_uop_0_ctrl_fcn_dw = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  rob_uop_0_ctrl_csr_cmd = _RAND_158[2:0];
  _RAND_159 = {1{`RANDOM}};
  rob_uop_0_ctrl_is_load = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  rob_uop_0_ctrl_is_sta = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  rob_uop_0_ctrl_is_std = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  rob_uop_0_iw_state = _RAND_162[1:0];
  _RAND_163 = {1{`RANDOM}};
  rob_uop_0_iw_p1_poisoned = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  rob_uop_0_iw_p2_poisoned = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  rob_uop_0_is_br = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  rob_uop_0_is_jalr = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  rob_uop_0_is_jal = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  rob_uop_0_is_sfb = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  rob_uop_0_br_mask = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  rob_uop_0_br_tag = _RAND_170[2:0];
  _RAND_171 = {1{`RANDOM}};
  rob_uop_0_ftq_idx = _RAND_171[3:0];
  _RAND_172 = {1{`RANDOM}};
  rob_uop_0_edge_inst = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  rob_uop_0_pc_lob = _RAND_173[5:0];
  _RAND_174 = {1{`RANDOM}};
  rob_uop_0_taken = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  rob_uop_0_imm_packed = _RAND_175[19:0];
  _RAND_176 = {1{`RANDOM}};
  rob_uop_0_csr_addr = _RAND_176[11:0];
  _RAND_177 = {1{`RANDOM}};
  rob_uop_0_rob_idx = _RAND_177[4:0];
  _RAND_178 = {1{`RANDOM}};
  rob_uop_0_ldq_idx = _RAND_178[2:0];
  _RAND_179 = {1{`RANDOM}};
  rob_uop_0_stq_idx = _RAND_179[2:0];
  _RAND_180 = {1{`RANDOM}};
  rob_uop_0_rxq_idx = _RAND_180[1:0];
  _RAND_181 = {1{`RANDOM}};
  rob_uop_0_pdst = _RAND_181[5:0];
  _RAND_182 = {1{`RANDOM}};
  rob_uop_0_prs1 = _RAND_182[5:0];
  _RAND_183 = {1{`RANDOM}};
  rob_uop_0_prs2 = _RAND_183[5:0];
  _RAND_184 = {1{`RANDOM}};
  rob_uop_0_prs3 = _RAND_184[5:0];
  _RAND_185 = {1{`RANDOM}};
  rob_uop_0_ppred = _RAND_185[3:0];
  _RAND_186 = {1{`RANDOM}};
  rob_uop_0_prs1_busy = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  rob_uop_0_prs2_busy = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  rob_uop_0_prs3_busy = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  rob_uop_0_ppred_busy = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  rob_uop_0_stale_pdst = _RAND_190[5:0];
  _RAND_191 = {1{`RANDOM}};
  rob_uop_0_exception = _RAND_191[0:0];
  _RAND_192 = {2{`RANDOM}};
  rob_uop_0_exc_cause = _RAND_192[63:0];
  _RAND_193 = {1{`RANDOM}};
  rob_uop_0_bypassable = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  rob_uop_0_mem_cmd = _RAND_194[4:0];
  _RAND_195 = {1{`RANDOM}};
  rob_uop_0_mem_size = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  rob_uop_0_mem_signed = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  rob_uop_0_is_fence = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  rob_uop_0_is_fencei = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  rob_uop_0_is_amo = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  rob_uop_0_uses_ldq = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  rob_uop_0_uses_stq = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  rob_uop_0_is_sys_pc2epc = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  rob_uop_0_is_unique = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  rob_uop_0_flush_on_commit = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  rob_uop_0_ldst_is_rs1 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  rob_uop_0_ldst = _RAND_206[5:0];
  _RAND_207 = {1{`RANDOM}};
  rob_uop_0_lrs1 = _RAND_207[5:0];
  _RAND_208 = {1{`RANDOM}};
  rob_uop_0_lrs2 = _RAND_208[5:0];
  _RAND_209 = {1{`RANDOM}};
  rob_uop_0_lrs3 = _RAND_209[5:0];
  _RAND_210 = {1{`RANDOM}};
  rob_uop_0_ldst_val = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  rob_uop_0_dst_rtype = _RAND_211[1:0];
  _RAND_212 = {1{`RANDOM}};
  rob_uop_0_lrs1_rtype = _RAND_212[1:0];
  _RAND_213 = {1{`RANDOM}};
  rob_uop_0_lrs2_rtype = _RAND_213[1:0];
  _RAND_214 = {1{`RANDOM}};
  rob_uop_0_frs3_en = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  rob_uop_0_fp_val = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  rob_uop_0_fp_single = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  rob_uop_0_xcpt_pf_if = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  rob_uop_0_xcpt_ae_if = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  rob_uop_0_xcpt_ma_if = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  rob_uop_0_bp_debug_if = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  rob_uop_0_bp_xcpt_if = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  rob_uop_0_debug_fsrc = _RAND_222[1:0];
  _RAND_223 = {1{`RANDOM}};
  rob_uop_0_debug_tsrc = _RAND_223[1:0];
  _RAND_224 = {1{`RANDOM}};
  rob_uop_1_uopc = _RAND_224[6:0];
  _RAND_225 = {1{`RANDOM}};
  rob_uop_1_inst = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  rob_uop_1_debug_inst = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  rob_uop_1_is_rvc = _RAND_227[0:0];
  _RAND_228 = {2{`RANDOM}};
  rob_uop_1_debug_pc = _RAND_228[39:0];
  _RAND_229 = {1{`RANDOM}};
  rob_uop_1_iq_type = _RAND_229[2:0];
  _RAND_230 = {1{`RANDOM}};
  rob_uop_1_fu_code = _RAND_230[9:0];
  _RAND_231 = {1{`RANDOM}};
  rob_uop_1_ctrl_br_type = _RAND_231[3:0];
  _RAND_232 = {1{`RANDOM}};
  rob_uop_1_ctrl_op1_sel = _RAND_232[1:0];
  _RAND_233 = {1{`RANDOM}};
  rob_uop_1_ctrl_op2_sel = _RAND_233[2:0];
  _RAND_234 = {1{`RANDOM}};
  rob_uop_1_ctrl_imm_sel = _RAND_234[2:0];
  _RAND_235 = {1{`RANDOM}};
  rob_uop_1_ctrl_op_fcn = _RAND_235[3:0];
  _RAND_236 = {1{`RANDOM}};
  rob_uop_1_ctrl_fcn_dw = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  rob_uop_1_ctrl_csr_cmd = _RAND_237[2:0];
  _RAND_238 = {1{`RANDOM}};
  rob_uop_1_ctrl_is_load = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  rob_uop_1_ctrl_is_sta = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  rob_uop_1_ctrl_is_std = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  rob_uop_1_iw_state = _RAND_241[1:0];
  _RAND_242 = {1{`RANDOM}};
  rob_uop_1_iw_p1_poisoned = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  rob_uop_1_iw_p2_poisoned = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  rob_uop_1_is_br = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  rob_uop_1_is_jalr = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  rob_uop_1_is_jal = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  rob_uop_1_is_sfb = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  rob_uop_1_br_mask = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  rob_uop_1_br_tag = _RAND_249[2:0];
  _RAND_250 = {1{`RANDOM}};
  rob_uop_1_ftq_idx = _RAND_250[3:0];
  _RAND_251 = {1{`RANDOM}};
  rob_uop_1_edge_inst = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  rob_uop_1_pc_lob = _RAND_252[5:0];
  _RAND_253 = {1{`RANDOM}};
  rob_uop_1_taken = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  rob_uop_1_imm_packed = _RAND_254[19:0];
  _RAND_255 = {1{`RANDOM}};
  rob_uop_1_csr_addr = _RAND_255[11:0];
  _RAND_256 = {1{`RANDOM}};
  rob_uop_1_rob_idx = _RAND_256[4:0];
  _RAND_257 = {1{`RANDOM}};
  rob_uop_1_ldq_idx = _RAND_257[2:0];
  _RAND_258 = {1{`RANDOM}};
  rob_uop_1_stq_idx = _RAND_258[2:0];
  _RAND_259 = {1{`RANDOM}};
  rob_uop_1_rxq_idx = _RAND_259[1:0];
  _RAND_260 = {1{`RANDOM}};
  rob_uop_1_pdst = _RAND_260[5:0];
  _RAND_261 = {1{`RANDOM}};
  rob_uop_1_prs1 = _RAND_261[5:0];
  _RAND_262 = {1{`RANDOM}};
  rob_uop_1_prs2 = _RAND_262[5:0];
  _RAND_263 = {1{`RANDOM}};
  rob_uop_1_prs3 = _RAND_263[5:0];
  _RAND_264 = {1{`RANDOM}};
  rob_uop_1_ppred = _RAND_264[3:0];
  _RAND_265 = {1{`RANDOM}};
  rob_uop_1_prs1_busy = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  rob_uop_1_prs2_busy = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  rob_uop_1_prs3_busy = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  rob_uop_1_ppred_busy = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  rob_uop_1_stale_pdst = _RAND_269[5:0];
  _RAND_270 = {1{`RANDOM}};
  rob_uop_1_exception = _RAND_270[0:0];
  _RAND_271 = {2{`RANDOM}};
  rob_uop_1_exc_cause = _RAND_271[63:0];
  _RAND_272 = {1{`RANDOM}};
  rob_uop_1_bypassable = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  rob_uop_1_mem_cmd = _RAND_273[4:0];
  _RAND_274 = {1{`RANDOM}};
  rob_uop_1_mem_size = _RAND_274[1:0];
  _RAND_275 = {1{`RANDOM}};
  rob_uop_1_mem_signed = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  rob_uop_1_is_fence = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  rob_uop_1_is_fencei = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  rob_uop_1_is_amo = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  rob_uop_1_uses_ldq = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  rob_uop_1_uses_stq = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  rob_uop_1_is_sys_pc2epc = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  rob_uop_1_is_unique = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  rob_uop_1_flush_on_commit = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  rob_uop_1_ldst_is_rs1 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  rob_uop_1_ldst = _RAND_285[5:0];
  _RAND_286 = {1{`RANDOM}};
  rob_uop_1_lrs1 = _RAND_286[5:0];
  _RAND_287 = {1{`RANDOM}};
  rob_uop_1_lrs2 = _RAND_287[5:0];
  _RAND_288 = {1{`RANDOM}};
  rob_uop_1_lrs3 = _RAND_288[5:0];
  _RAND_289 = {1{`RANDOM}};
  rob_uop_1_ldst_val = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  rob_uop_1_dst_rtype = _RAND_290[1:0];
  _RAND_291 = {1{`RANDOM}};
  rob_uop_1_lrs1_rtype = _RAND_291[1:0];
  _RAND_292 = {1{`RANDOM}};
  rob_uop_1_lrs2_rtype = _RAND_292[1:0];
  _RAND_293 = {1{`RANDOM}};
  rob_uop_1_frs3_en = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  rob_uop_1_fp_val = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  rob_uop_1_fp_single = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  rob_uop_1_xcpt_pf_if = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  rob_uop_1_xcpt_ae_if = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  rob_uop_1_xcpt_ma_if = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  rob_uop_1_bp_debug_if = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  rob_uop_1_bp_xcpt_if = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  rob_uop_1_debug_fsrc = _RAND_301[1:0];
  _RAND_302 = {1{`RANDOM}};
  rob_uop_1_debug_tsrc = _RAND_302[1:0];
  _RAND_303 = {1{`RANDOM}};
  rob_uop_2_uopc = _RAND_303[6:0];
  _RAND_304 = {1{`RANDOM}};
  rob_uop_2_inst = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  rob_uop_2_debug_inst = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  rob_uop_2_is_rvc = _RAND_306[0:0];
  _RAND_307 = {2{`RANDOM}};
  rob_uop_2_debug_pc = _RAND_307[39:0];
  _RAND_308 = {1{`RANDOM}};
  rob_uop_2_iq_type = _RAND_308[2:0];
  _RAND_309 = {1{`RANDOM}};
  rob_uop_2_fu_code = _RAND_309[9:0];
  _RAND_310 = {1{`RANDOM}};
  rob_uop_2_ctrl_br_type = _RAND_310[3:0];
  _RAND_311 = {1{`RANDOM}};
  rob_uop_2_ctrl_op1_sel = _RAND_311[1:0];
  _RAND_312 = {1{`RANDOM}};
  rob_uop_2_ctrl_op2_sel = _RAND_312[2:0];
  _RAND_313 = {1{`RANDOM}};
  rob_uop_2_ctrl_imm_sel = _RAND_313[2:0];
  _RAND_314 = {1{`RANDOM}};
  rob_uop_2_ctrl_op_fcn = _RAND_314[3:0];
  _RAND_315 = {1{`RANDOM}};
  rob_uop_2_ctrl_fcn_dw = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  rob_uop_2_ctrl_csr_cmd = _RAND_316[2:0];
  _RAND_317 = {1{`RANDOM}};
  rob_uop_2_ctrl_is_load = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  rob_uop_2_ctrl_is_sta = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  rob_uop_2_ctrl_is_std = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  rob_uop_2_iw_state = _RAND_320[1:0];
  _RAND_321 = {1{`RANDOM}};
  rob_uop_2_iw_p1_poisoned = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  rob_uop_2_iw_p2_poisoned = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  rob_uop_2_is_br = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  rob_uop_2_is_jalr = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  rob_uop_2_is_jal = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  rob_uop_2_is_sfb = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  rob_uop_2_br_mask = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  rob_uop_2_br_tag = _RAND_328[2:0];
  _RAND_329 = {1{`RANDOM}};
  rob_uop_2_ftq_idx = _RAND_329[3:0];
  _RAND_330 = {1{`RANDOM}};
  rob_uop_2_edge_inst = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  rob_uop_2_pc_lob = _RAND_331[5:0];
  _RAND_332 = {1{`RANDOM}};
  rob_uop_2_taken = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  rob_uop_2_imm_packed = _RAND_333[19:0];
  _RAND_334 = {1{`RANDOM}};
  rob_uop_2_csr_addr = _RAND_334[11:0];
  _RAND_335 = {1{`RANDOM}};
  rob_uop_2_rob_idx = _RAND_335[4:0];
  _RAND_336 = {1{`RANDOM}};
  rob_uop_2_ldq_idx = _RAND_336[2:0];
  _RAND_337 = {1{`RANDOM}};
  rob_uop_2_stq_idx = _RAND_337[2:0];
  _RAND_338 = {1{`RANDOM}};
  rob_uop_2_rxq_idx = _RAND_338[1:0];
  _RAND_339 = {1{`RANDOM}};
  rob_uop_2_pdst = _RAND_339[5:0];
  _RAND_340 = {1{`RANDOM}};
  rob_uop_2_prs1 = _RAND_340[5:0];
  _RAND_341 = {1{`RANDOM}};
  rob_uop_2_prs2 = _RAND_341[5:0];
  _RAND_342 = {1{`RANDOM}};
  rob_uop_2_prs3 = _RAND_342[5:0];
  _RAND_343 = {1{`RANDOM}};
  rob_uop_2_ppred = _RAND_343[3:0];
  _RAND_344 = {1{`RANDOM}};
  rob_uop_2_prs1_busy = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  rob_uop_2_prs2_busy = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  rob_uop_2_prs3_busy = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  rob_uop_2_ppred_busy = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  rob_uop_2_stale_pdst = _RAND_348[5:0];
  _RAND_349 = {1{`RANDOM}};
  rob_uop_2_exception = _RAND_349[0:0];
  _RAND_350 = {2{`RANDOM}};
  rob_uop_2_exc_cause = _RAND_350[63:0];
  _RAND_351 = {1{`RANDOM}};
  rob_uop_2_bypassable = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  rob_uop_2_mem_cmd = _RAND_352[4:0];
  _RAND_353 = {1{`RANDOM}};
  rob_uop_2_mem_size = _RAND_353[1:0];
  _RAND_354 = {1{`RANDOM}};
  rob_uop_2_mem_signed = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  rob_uop_2_is_fence = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  rob_uop_2_is_fencei = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  rob_uop_2_is_amo = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  rob_uop_2_uses_ldq = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  rob_uop_2_uses_stq = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  rob_uop_2_is_sys_pc2epc = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  rob_uop_2_is_unique = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  rob_uop_2_flush_on_commit = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  rob_uop_2_ldst_is_rs1 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  rob_uop_2_ldst = _RAND_364[5:0];
  _RAND_365 = {1{`RANDOM}};
  rob_uop_2_lrs1 = _RAND_365[5:0];
  _RAND_366 = {1{`RANDOM}};
  rob_uop_2_lrs2 = _RAND_366[5:0];
  _RAND_367 = {1{`RANDOM}};
  rob_uop_2_lrs3 = _RAND_367[5:0];
  _RAND_368 = {1{`RANDOM}};
  rob_uop_2_ldst_val = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  rob_uop_2_dst_rtype = _RAND_369[1:0];
  _RAND_370 = {1{`RANDOM}};
  rob_uop_2_lrs1_rtype = _RAND_370[1:0];
  _RAND_371 = {1{`RANDOM}};
  rob_uop_2_lrs2_rtype = _RAND_371[1:0];
  _RAND_372 = {1{`RANDOM}};
  rob_uop_2_frs3_en = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  rob_uop_2_fp_val = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  rob_uop_2_fp_single = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  rob_uop_2_xcpt_pf_if = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  rob_uop_2_xcpt_ae_if = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  rob_uop_2_xcpt_ma_if = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  rob_uop_2_bp_debug_if = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  rob_uop_2_bp_xcpt_if = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  rob_uop_2_debug_fsrc = _RAND_380[1:0];
  _RAND_381 = {1{`RANDOM}};
  rob_uop_2_debug_tsrc = _RAND_381[1:0];
  _RAND_382 = {1{`RANDOM}};
  rob_uop_3_uopc = _RAND_382[6:0];
  _RAND_383 = {1{`RANDOM}};
  rob_uop_3_inst = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  rob_uop_3_debug_inst = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  rob_uop_3_is_rvc = _RAND_385[0:0];
  _RAND_386 = {2{`RANDOM}};
  rob_uop_3_debug_pc = _RAND_386[39:0];
  _RAND_387 = {1{`RANDOM}};
  rob_uop_3_iq_type = _RAND_387[2:0];
  _RAND_388 = {1{`RANDOM}};
  rob_uop_3_fu_code = _RAND_388[9:0];
  _RAND_389 = {1{`RANDOM}};
  rob_uop_3_ctrl_br_type = _RAND_389[3:0];
  _RAND_390 = {1{`RANDOM}};
  rob_uop_3_ctrl_op1_sel = _RAND_390[1:0];
  _RAND_391 = {1{`RANDOM}};
  rob_uop_3_ctrl_op2_sel = _RAND_391[2:0];
  _RAND_392 = {1{`RANDOM}};
  rob_uop_3_ctrl_imm_sel = _RAND_392[2:0];
  _RAND_393 = {1{`RANDOM}};
  rob_uop_3_ctrl_op_fcn = _RAND_393[3:0];
  _RAND_394 = {1{`RANDOM}};
  rob_uop_3_ctrl_fcn_dw = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  rob_uop_3_ctrl_csr_cmd = _RAND_395[2:0];
  _RAND_396 = {1{`RANDOM}};
  rob_uop_3_ctrl_is_load = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  rob_uop_3_ctrl_is_sta = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  rob_uop_3_ctrl_is_std = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  rob_uop_3_iw_state = _RAND_399[1:0];
  _RAND_400 = {1{`RANDOM}};
  rob_uop_3_iw_p1_poisoned = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  rob_uop_3_iw_p2_poisoned = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  rob_uop_3_is_br = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  rob_uop_3_is_jalr = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  rob_uop_3_is_jal = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  rob_uop_3_is_sfb = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  rob_uop_3_br_mask = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  rob_uop_3_br_tag = _RAND_407[2:0];
  _RAND_408 = {1{`RANDOM}};
  rob_uop_3_ftq_idx = _RAND_408[3:0];
  _RAND_409 = {1{`RANDOM}};
  rob_uop_3_edge_inst = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  rob_uop_3_pc_lob = _RAND_410[5:0];
  _RAND_411 = {1{`RANDOM}};
  rob_uop_3_taken = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  rob_uop_3_imm_packed = _RAND_412[19:0];
  _RAND_413 = {1{`RANDOM}};
  rob_uop_3_csr_addr = _RAND_413[11:0];
  _RAND_414 = {1{`RANDOM}};
  rob_uop_3_rob_idx = _RAND_414[4:0];
  _RAND_415 = {1{`RANDOM}};
  rob_uop_3_ldq_idx = _RAND_415[2:0];
  _RAND_416 = {1{`RANDOM}};
  rob_uop_3_stq_idx = _RAND_416[2:0];
  _RAND_417 = {1{`RANDOM}};
  rob_uop_3_rxq_idx = _RAND_417[1:0];
  _RAND_418 = {1{`RANDOM}};
  rob_uop_3_pdst = _RAND_418[5:0];
  _RAND_419 = {1{`RANDOM}};
  rob_uop_3_prs1 = _RAND_419[5:0];
  _RAND_420 = {1{`RANDOM}};
  rob_uop_3_prs2 = _RAND_420[5:0];
  _RAND_421 = {1{`RANDOM}};
  rob_uop_3_prs3 = _RAND_421[5:0];
  _RAND_422 = {1{`RANDOM}};
  rob_uop_3_ppred = _RAND_422[3:0];
  _RAND_423 = {1{`RANDOM}};
  rob_uop_3_prs1_busy = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  rob_uop_3_prs2_busy = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  rob_uop_3_prs3_busy = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  rob_uop_3_ppred_busy = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  rob_uop_3_stale_pdst = _RAND_427[5:0];
  _RAND_428 = {1{`RANDOM}};
  rob_uop_3_exception = _RAND_428[0:0];
  _RAND_429 = {2{`RANDOM}};
  rob_uop_3_exc_cause = _RAND_429[63:0];
  _RAND_430 = {1{`RANDOM}};
  rob_uop_3_bypassable = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  rob_uop_3_mem_cmd = _RAND_431[4:0];
  _RAND_432 = {1{`RANDOM}};
  rob_uop_3_mem_size = _RAND_432[1:0];
  _RAND_433 = {1{`RANDOM}};
  rob_uop_3_mem_signed = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  rob_uop_3_is_fence = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  rob_uop_3_is_fencei = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  rob_uop_3_is_amo = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  rob_uop_3_uses_ldq = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  rob_uop_3_uses_stq = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  rob_uop_3_is_sys_pc2epc = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  rob_uop_3_is_unique = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  rob_uop_3_flush_on_commit = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  rob_uop_3_ldst_is_rs1 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  rob_uop_3_ldst = _RAND_443[5:0];
  _RAND_444 = {1{`RANDOM}};
  rob_uop_3_lrs1 = _RAND_444[5:0];
  _RAND_445 = {1{`RANDOM}};
  rob_uop_3_lrs2 = _RAND_445[5:0];
  _RAND_446 = {1{`RANDOM}};
  rob_uop_3_lrs3 = _RAND_446[5:0];
  _RAND_447 = {1{`RANDOM}};
  rob_uop_3_ldst_val = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  rob_uop_3_dst_rtype = _RAND_448[1:0];
  _RAND_449 = {1{`RANDOM}};
  rob_uop_3_lrs1_rtype = _RAND_449[1:0];
  _RAND_450 = {1{`RANDOM}};
  rob_uop_3_lrs2_rtype = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  rob_uop_3_frs3_en = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  rob_uop_3_fp_val = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  rob_uop_3_fp_single = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  rob_uop_3_xcpt_pf_if = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  rob_uop_3_xcpt_ae_if = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  rob_uop_3_xcpt_ma_if = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  rob_uop_3_bp_debug_if = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  rob_uop_3_bp_xcpt_if = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  rob_uop_3_debug_fsrc = _RAND_459[1:0];
  _RAND_460 = {1{`RANDOM}};
  rob_uop_3_debug_tsrc = _RAND_460[1:0];
  _RAND_461 = {1{`RANDOM}};
  rob_uop_4_uopc = _RAND_461[6:0];
  _RAND_462 = {1{`RANDOM}};
  rob_uop_4_inst = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  rob_uop_4_debug_inst = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  rob_uop_4_is_rvc = _RAND_464[0:0];
  _RAND_465 = {2{`RANDOM}};
  rob_uop_4_debug_pc = _RAND_465[39:0];
  _RAND_466 = {1{`RANDOM}};
  rob_uop_4_iq_type = _RAND_466[2:0];
  _RAND_467 = {1{`RANDOM}};
  rob_uop_4_fu_code = _RAND_467[9:0];
  _RAND_468 = {1{`RANDOM}};
  rob_uop_4_ctrl_br_type = _RAND_468[3:0];
  _RAND_469 = {1{`RANDOM}};
  rob_uop_4_ctrl_op1_sel = _RAND_469[1:0];
  _RAND_470 = {1{`RANDOM}};
  rob_uop_4_ctrl_op2_sel = _RAND_470[2:0];
  _RAND_471 = {1{`RANDOM}};
  rob_uop_4_ctrl_imm_sel = _RAND_471[2:0];
  _RAND_472 = {1{`RANDOM}};
  rob_uop_4_ctrl_op_fcn = _RAND_472[3:0];
  _RAND_473 = {1{`RANDOM}};
  rob_uop_4_ctrl_fcn_dw = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  rob_uop_4_ctrl_csr_cmd = _RAND_474[2:0];
  _RAND_475 = {1{`RANDOM}};
  rob_uop_4_ctrl_is_load = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  rob_uop_4_ctrl_is_sta = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  rob_uop_4_ctrl_is_std = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  rob_uop_4_iw_state = _RAND_478[1:0];
  _RAND_479 = {1{`RANDOM}};
  rob_uop_4_iw_p1_poisoned = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  rob_uop_4_iw_p2_poisoned = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  rob_uop_4_is_br = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  rob_uop_4_is_jalr = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  rob_uop_4_is_jal = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  rob_uop_4_is_sfb = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  rob_uop_4_br_mask = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  rob_uop_4_br_tag = _RAND_486[2:0];
  _RAND_487 = {1{`RANDOM}};
  rob_uop_4_ftq_idx = _RAND_487[3:0];
  _RAND_488 = {1{`RANDOM}};
  rob_uop_4_edge_inst = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  rob_uop_4_pc_lob = _RAND_489[5:0];
  _RAND_490 = {1{`RANDOM}};
  rob_uop_4_taken = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  rob_uop_4_imm_packed = _RAND_491[19:0];
  _RAND_492 = {1{`RANDOM}};
  rob_uop_4_csr_addr = _RAND_492[11:0];
  _RAND_493 = {1{`RANDOM}};
  rob_uop_4_rob_idx = _RAND_493[4:0];
  _RAND_494 = {1{`RANDOM}};
  rob_uop_4_ldq_idx = _RAND_494[2:0];
  _RAND_495 = {1{`RANDOM}};
  rob_uop_4_stq_idx = _RAND_495[2:0];
  _RAND_496 = {1{`RANDOM}};
  rob_uop_4_rxq_idx = _RAND_496[1:0];
  _RAND_497 = {1{`RANDOM}};
  rob_uop_4_pdst = _RAND_497[5:0];
  _RAND_498 = {1{`RANDOM}};
  rob_uop_4_prs1 = _RAND_498[5:0];
  _RAND_499 = {1{`RANDOM}};
  rob_uop_4_prs2 = _RAND_499[5:0];
  _RAND_500 = {1{`RANDOM}};
  rob_uop_4_prs3 = _RAND_500[5:0];
  _RAND_501 = {1{`RANDOM}};
  rob_uop_4_ppred = _RAND_501[3:0];
  _RAND_502 = {1{`RANDOM}};
  rob_uop_4_prs1_busy = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  rob_uop_4_prs2_busy = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  rob_uop_4_prs3_busy = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  rob_uop_4_ppred_busy = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  rob_uop_4_stale_pdst = _RAND_506[5:0];
  _RAND_507 = {1{`RANDOM}};
  rob_uop_4_exception = _RAND_507[0:0];
  _RAND_508 = {2{`RANDOM}};
  rob_uop_4_exc_cause = _RAND_508[63:0];
  _RAND_509 = {1{`RANDOM}};
  rob_uop_4_bypassable = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  rob_uop_4_mem_cmd = _RAND_510[4:0];
  _RAND_511 = {1{`RANDOM}};
  rob_uop_4_mem_size = _RAND_511[1:0];
  _RAND_512 = {1{`RANDOM}};
  rob_uop_4_mem_signed = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  rob_uop_4_is_fence = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  rob_uop_4_is_fencei = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  rob_uop_4_is_amo = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  rob_uop_4_uses_ldq = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  rob_uop_4_uses_stq = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  rob_uop_4_is_sys_pc2epc = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  rob_uop_4_is_unique = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  rob_uop_4_flush_on_commit = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  rob_uop_4_ldst_is_rs1 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  rob_uop_4_ldst = _RAND_522[5:0];
  _RAND_523 = {1{`RANDOM}};
  rob_uop_4_lrs1 = _RAND_523[5:0];
  _RAND_524 = {1{`RANDOM}};
  rob_uop_4_lrs2 = _RAND_524[5:0];
  _RAND_525 = {1{`RANDOM}};
  rob_uop_4_lrs3 = _RAND_525[5:0];
  _RAND_526 = {1{`RANDOM}};
  rob_uop_4_ldst_val = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  rob_uop_4_dst_rtype = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  rob_uop_4_lrs1_rtype = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  rob_uop_4_lrs2_rtype = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  rob_uop_4_frs3_en = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  rob_uop_4_fp_val = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  rob_uop_4_fp_single = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  rob_uop_4_xcpt_pf_if = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  rob_uop_4_xcpt_ae_if = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  rob_uop_4_xcpt_ma_if = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  rob_uop_4_bp_debug_if = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  rob_uop_4_bp_xcpt_if = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  rob_uop_4_debug_fsrc = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  rob_uop_4_debug_tsrc = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  rob_uop_5_uopc = _RAND_540[6:0];
  _RAND_541 = {1{`RANDOM}};
  rob_uop_5_inst = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  rob_uop_5_debug_inst = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  rob_uop_5_is_rvc = _RAND_543[0:0];
  _RAND_544 = {2{`RANDOM}};
  rob_uop_5_debug_pc = _RAND_544[39:0];
  _RAND_545 = {1{`RANDOM}};
  rob_uop_5_iq_type = _RAND_545[2:0];
  _RAND_546 = {1{`RANDOM}};
  rob_uop_5_fu_code = _RAND_546[9:0];
  _RAND_547 = {1{`RANDOM}};
  rob_uop_5_ctrl_br_type = _RAND_547[3:0];
  _RAND_548 = {1{`RANDOM}};
  rob_uop_5_ctrl_op1_sel = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  rob_uop_5_ctrl_op2_sel = _RAND_549[2:0];
  _RAND_550 = {1{`RANDOM}};
  rob_uop_5_ctrl_imm_sel = _RAND_550[2:0];
  _RAND_551 = {1{`RANDOM}};
  rob_uop_5_ctrl_op_fcn = _RAND_551[3:0];
  _RAND_552 = {1{`RANDOM}};
  rob_uop_5_ctrl_fcn_dw = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  rob_uop_5_ctrl_csr_cmd = _RAND_553[2:0];
  _RAND_554 = {1{`RANDOM}};
  rob_uop_5_ctrl_is_load = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  rob_uop_5_ctrl_is_sta = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  rob_uop_5_ctrl_is_std = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  rob_uop_5_iw_state = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  rob_uop_5_iw_p1_poisoned = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  rob_uop_5_iw_p2_poisoned = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  rob_uop_5_is_br = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  rob_uop_5_is_jalr = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  rob_uop_5_is_jal = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  rob_uop_5_is_sfb = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  rob_uop_5_br_mask = _RAND_564[7:0];
  _RAND_565 = {1{`RANDOM}};
  rob_uop_5_br_tag = _RAND_565[2:0];
  _RAND_566 = {1{`RANDOM}};
  rob_uop_5_ftq_idx = _RAND_566[3:0];
  _RAND_567 = {1{`RANDOM}};
  rob_uop_5_edge_inst = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  rob_uop_5_pc_lob = _RAND_568[5:0];
  _RAND_569 = {1{`RANDOM}};
  rob_uop_5_taken = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  rob_uop_5_imm_packed = _RAND_570[19:0];
  _RAND_571 = {1{`RANDOM}};
  rob_uop_5_csr_addr = _RAND_571[11:0];
  _RAND_572 = {1{`RANDOM}};
  rob_uop_5_rob_idx = _RAND_572[4:0];
  _RAND_573 = {1{`RANDOM}};
  rob_uop_5_ldq_idx = _RAND_573[2:0];
  _RAND_574 = {1{`RANDOM}};
  rob_uop_5_stq_idx = _RAND_574[2:0];
  _RAND_575 = {1{`RANDOM}};
  rob_uop_5_rxq_idx = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  rob_uop_5_pdst = _RAND_576[5:0];
  _RAND_577 = {1{`RANDOM}};
  rob_uop_5_prs1 = _RAND_577[5:0];
  _RAND_578 = {1{`RANDOM}};
  rob_uop_5_prs2 = _RAND_578[5:0];
  _RAND_579 = {1{`RANDOM}};
  rob_uop_5_prs3 = _RAND_579[5:0];
  _RAND_580 = {1{`RANDOM}};
  rob_uop_5_ppred = _RAND_580[3:0];
  _RAND_581 = {1{`RANDOM}};
  rob_uop_5_prs1_busy = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  rob_uop_5_prs2_busy = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  rob_uop_5_prs3_busy = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  rob_uop_5_ppred_busy = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  rob_uop_5_stale_pdst = _RAND_585[5:0];
  _RAND_586 = {1{`RANDOM}};
  rob_uop_5_exception = _RAND_586[0:0];
  _RAND_587 = {2{`RANDOM}};
  rob_uop_5_exc_cause = _RAND_587[63:0];
  _RAND_588 = {1{`RANDOM}};
  rob_uop_5_bypassable = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  rob_uop_5_mem_cmd = _RAND_589[4:0];
  _RAND_590 = {1{`RANDOM}};
  rob_uop_5_mem_size = _RAND_590[1:0];
  _RAND_591 = {1{`RANDOM}};
  rob_uop_5_mem_signed = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  rob_uop_5_is_fence = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  rob_uop_5_is_fencei = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  rob_uop_5_is_amo = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  rob_uop_5_uses_ldq = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  rob_uop_5_uses_stq = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  rob_uop_5_is_sys_pc2epc = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  rob_uop_5_is_unique = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  rob_uop_5_flush_on_commit = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  rob_uop_5_ldst_is_rs1 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  rob_uop_5_ldst = _RAND_601[5:0];
  _RAND_602 = {1{`RANDOM}};
  rob_uop_5_lrs1 = _RAND_602[5:0];
  _RAND_603 = {1{`RANDOM}};
  rob_uop_5_lrs2 = _RAND_603[5:0];
  _RAND_604 = {1{`RANDOM}};
  rob_uop_5_lrs3 = _RAND_604[5:0];
  _RAND_605 = {1{`RANDOM}};
  rob_uop_5_ldst_val = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  rob_uop_5_dst_rtype = _RAND_606[1:0];
  _RAND_607 = {1{`RANDOM}};
  rob_uop_5_lrs1_rtype = _RAND_607[1:0];
  _RAND_608 = {1{`RANDOM}};
  rob_uop_5_lrs2_rtype = _RAND_608[1:0];
  _RAND_609 = {1{`RANDOM}};
  rob_uop_5_frs3_en = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  rob_uop_5_fp_val = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  rob_uop_5_fp_single = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  rob_uop_5_xcpt_pf_if = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  rob_uop_5_xcpt_ae_if = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  rob_uop_5_xcpt_ma_if = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  rob_uop_5_bp_debug_if = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  rob_uop_5_bp_xcpt_if = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  rob_uop_5_debug_fsrc = _RAND_617[1:0];
  _RAND_618 = {1{`RANDOM}};
  rob_uop_5_debug_tsrc = _RAND_618[1:0];
  _RAND_619 = {1{`RANDOM}};
  rob_uop_6_uopc = _RAND_619[6:0];
  _RAND_620 = {1{`RANDOM}};
  rob_uop_6_inst = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  rob_uop_6_debug_inst = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  rob_uop_6_is_rvc = _RAND_622[0:0];
  _RAND_623 = {2{`RANDOM}};
  rob_uop_6_debug_pc = _RAND_623[39:0];
  _RAND_624 = {1{`RANDOM}};
  rob_uop_6_iq_type = _RAND_624[2:0];
  _RAND_625 = {1{`RANDOM}};
  rob_uop_6_fu_code = _RAND_625[9:0];
  _RAND_626 = {1{`RANDOM}};
  rob_uop_6_ctrl_br_type = _RAND_626[3:0];
  _RAND_627 = {1{`RANDOM}};
  rob_uop_6_ctrl_op1_sel = _RAND_627[1:0];
  _RAND_628 = {1{`RANDOM}};
  rob_uop_6_ctrl_op2_sel = _RAND_628[2:0];
  _RAND_629 = {1{`RANDOM}};
  rob_uop_6_ctrl_imm_sel = _RAND_629[2:0];
  _RAND_630 = {1{`RANDOM}};
  rob_uop_6_ctrl_op_fcn = _RAND_630[3:0];
  _RAND_631 = {1{`RANDOM}};
  rob_uop_6_ctrl_fcn_dw = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  rob_uop_6_ctrl_csr_cmd = _RAND_632[2:0];
  _RAND_633 = {1{`RANDOM}};
  rob_uop_6_ctrl_is_load = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  rob_uop_6_ctrl_is_sta = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  rob_uop_6_ctrl_is_std = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  rob_uop_6_iw_state = _RAND_636[1:0];
  _RAND_637 = {1{`RANDOM}};
  rob_uop_6_iw_p1_poisoned = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  rob_uop_6_iw_p2_poisoned = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  rob_uop_6_is_br = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  rob_uop_6_is_jalr = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  rob_uop_6_is_jal = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  rob_uop_6_is_sfb = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  rob_uop_6_br_mask = _RAND_643[7:0];
  _RAND_644 = {1{`RANDOM}};
  rob_uop_6_br_tag = _RAND_644[2:0];
  _RAND_645 = {1{`RANDOM}};
  rob_uop_6_ftq_idx = _RAND_645[3:0];
  _RAND_646 = {1{`RANDOM}};
  rob_uop_6_edge_inst = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  rob_uop_6_pc_lob = _RAND_647[5:0];
  _RAND_648 = {1{`RANDOM}};
  rob_uop_6_taken = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  rob_uop_6_imm_packed = _RAND_649[19:0];
  _RAND_650 = {1{`RANDOM}};
  rob_uop_6_csr_addr = _RAND_650[11:0];
  _RAND_651 = {1{`RANDOM}};
  rob_uop_6_rob_idx = _RAND_651[4:0];
  _RAND_652 = {1{`RANDOM}};
  rob_uop_6_ldq_idx = _RAND_652[2:0];
  _RAND_653 = {1{`RANDOM}};
  rob_uop_6_stq_idx = _RAND_653[2:0];
  _RAND_654 = {1{`RANDOM}};
  rob_uop_6_rxq_idx = _RAND_654[1:0];
  _RAND_655 = {1{`RANDOM}};
  rob_uop_6_pdst = _RAND_655[5:0];
  _RAND_656 = {1{`RANDOM}};
  rob_uop_6_prs1 = _RAND_656[5:0];
  _RAND_657 = {1{`RANDOM}};
  rob_uop_6_prs2 = _RAND_657[5:0];
  _RAND_658 = {1{`RANDOM}};
  rob_uop_6_prs3 = _RAND_658[5:0];
  _RAND_659 = {1{`RANDOM}};
  rob_uop_6_ppred = _RAND_659[3:0];
  _RAND_660 = {1{`RANDOM}};
  rob_uop_6_prs1_busy = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  rob_uop_6_prs2_busy = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  rob_uop_6_prs3_busy = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  rob_uop_6_ppred_busy = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  rob_uop_6_stale_pdst = _RAND_664[5:0];
  _RAND_665 = {1{`RANDOM}};
  rob_uop_6_exception = _RAND_665[0:0];
  _RAND_666 = {2{`RANDOM}};
  rob_uop_6_exc_cause = _RAND_666[63:0];
  _RAND_667 = {1{`RANDOM}};
  rob_uop_6_bypassable = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  rob_uop_6_mem_cmd = _RAND_668[4:0];
  _RAND_669 = {1{`RANDOM}};
  rob_uop_6_mem_size = _RAND_669[1:0];
  _RAND_670 = {1{`RANDOM}};
  rob_uop_6_mem_signed = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  rob_uop_6_is_fence = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  rob_uop_6_is_fencei = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  rob_uop_6_is_amo = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  rob_uop_6_uses_ldq = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  rob_uop_6_uses_stq = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  rob_uop_6_is_sys_pc2epc = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  rob_uop_6_is_unique = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  rob_uop_6_flush_on_commit = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  rob_uop_6_ldst_is_rs1 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  rob_uop_6_ldst = _RAND_680[5:0];
  _RAND_681 = {1{`RANDOM}};
  rob_uop_6_lrs1 = _RAND_681[5:0];
  _RAND_682 = {1{`RANDOM}};
  rob_uop_6_lrs2 = _RAND_682[5:0];
  _RAND_683 = {1{`RANDOM}};
  rob_uop_6_lrs3 = _RAND_683[5:0];
  _RAND_684 = {1{`RANDOM}};
  rob_uop_6_ldst_val = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  rob_uop_6_dst_rtype = _RAND_685[1:0];
  _RAND_686 = {1{`RANDOM}};
  rob_uop_6_lrs1_rtype = _RAND_686[1:0];
  _RAND_687 = {1{`RANDOM}};
  rob_uop_6_lrs2_rtype = _RAND_687[1:0];
  _RAND_688 = {1{`RANDOM}};
  rob_uop_6_frs3_en = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  rob_uop_6_fp_val = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  rob_uop_6_fp_single = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  rob_uop_6_xcpt_pf_if = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  rob_uop_6_xcpt_ae_if = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  rob_uop_6_xcpt_ma_if = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  rob_uop_6_bp_debug_if = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  rob_uop_6_bp_xcpt_if = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  rob_uop_6_debug_fsrc = _RAND_696[1:0];
  _RAND_697 = {1{`RANDOM}};
  rob_uop_6_debug_tsrc = _RAND_697[1:0];
  _RAND_698 = {1{`RANDOM}};
  rob_uop_7_uopc = _RAND_698[6:0];
  _RAND_699 = {1{`RANDOM}};
  rob_uop_7_inst = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  rob_uop_7_debug_inst = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  rob_uop_7_is_rvc = _RAND_701[0:0];
  _RAND_702 = {2{`RANDOM}};
  rob_uop_7_debug_pc = _RAND_702[39:0];
  _RAND_703 = {1{`RANDOM}};
  rob_uop_7_iq_type = _RAND_703[2:0];
  _RAND_704 = {1{`RANDOM}};
  rob_uop_7_fu_code = _RAND_704[9:0];
  _RAND_705 = {1{`RANDOM}};
  rob_uop_7_ctrl_br_type = _RAND_705[3:0];
  _RAND_706 = {1{`RANDOM}};
  rob_uop_7_ctrl_op1_sel = _RAND_706[1:0];
  _RAND_707 = {1{`RANDOM}};
  rob_uop_7_ctrl_op2_sel = _RAND_707[2:0];
  _RAND_708 = {1{`RANDOM}};
  rob_uop_7_ctrl_imm_sel = _RAND_708[2:0];
  _RAND_709 = {1{`RANDOM}};
  rob_uop_7_ctrl_op_fcn = _RAND_709[3:0];
  _RAND_710 = {1{`RANDOM}};
  rob_uop_7_ctrl_fcn_dw = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  rob_uop_7_ctrl_csr_cmd = _RAND_711[2:0];
  _RAND_712 = {1{`RANDOM}};
  rob_uop_7_ctrl_is_load = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  rob_uop_7_ctrl_is_sta = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  rob_uop_7_ctrl_is_std = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  rob_uop_7_iw_state = _RAND_715[1:0];
  _RAND_716 = {1{`RANDOM}};
  rob_uop_7_iw_p1_poisoned = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  rob_uop_7_iw_p2_poisoned = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  rob_uop_7_is_br = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  rob_uop_7_is_jalr = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  rob_uop_7_is_jal = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  rob_uop_7_is_sfb = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  rob_uop_7_br_mask = _RAND_722[7:0];
  _RAND_723 = {1{`RANDOM}};
  rob_uop_7_br_tag = _RAND_723[2:0];
  _RAND_724 = {1{`RANDOM}};
  rob_uop_7_ftq_idx = _RAND_724[3:0];
  _RAND_725 = {1{`RANDOM}};
  rob_uop_7_edge_inst = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  rob_uop_7_pc_lob = _RAND_726[5:0];
  _RAND_727 = {1{`RANDOM}};
  rob_uop_7_taken = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  rob_uop_7_imm_packed = _RAND_728[19:0];
  _RAND_729 = {1{`RANDOM}};
  rob_uop_7_csr_addr = _RAND_729[11:0];
  _RAND_730 = {1{`RANDOM}};
  rob_uop_7_rob_idx = _RAND_730[4:0];
  _RAND_731 = {1{`RANDOM}};
  rob_uop_7_ldq_idx = _RAND_731[2:0];
  _RAND_732 = {1{`RANDOM}};
  rob_uop_7_stq_idx = _RAND_732[2:0];
  _RAND_733 = {1{`RANDOM}};
  rob_uop_7_rxq_idx = _RAND_733[1:0];
  _RAND_734 = {1{`RANDOM}};
  rob_uop_7_pdst = _RAND_734[5:0];
  _RAND_735 = {1{`RANDOM}};
  rob_uop_7_prs1 = _RAND_735[5:0];
  _RAND_736 = {1{`RANDOM}};
  rob_uop_7_prs2 = _RAND_736[5:0];
  _RAND_737 = {1{`RANDOM}};
  rob_uop_7_prs3 = _RAND_737[5:0];
  _RAND_738 = {1{`RANDOM}};
  rob_uop_7_ppred = _RAND_738[3:0];
  _RAND_739 = {1{`RANDOM}};
  rob_uop_7_prs1_busy = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  rob_uop_7_prs2_busy = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  rob_uop_7_prs3_busy = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  rob_uop_7_ppred_busy = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  rob_uop_7_stale_pdst = _RAND_743[5:0];
  _RAND_744 = {1{`RANDOM}};
  rob_uop_7_exception = _RAND_744[0:0];
  _RAND_745 = {2{`RANDOM}};
  rob_uop_7_exc_cause = _RAND_745[63:0];
  _RAND_746 = {1{`RANDOM}};
  rob_uop_7_bypassable = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  rob_uop_7_mem_cmd = _RAND_747[4:0];
  _RAND_748 = {1{`RANDOM}};
  rob_uop_7_mem_size = _RAND_748[1:0];
  _RAND_749 = {1{`RANDOM}};
  rob_uop_7_mem_signed = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  rob_uop_7_is_fence = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  rob_uop_7_is_fencei = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  rob_uop_7_is_amo = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  rob_uop_7_uses_ldq = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  rob_uop_7_uses_stq = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  rob_uop_7_is_sys_pc2epc = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  rob_uop_7_is_unique = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  rob_uop_7_flush_on_commit = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  rob_uop_7_ldst_is_rs1 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  rob_uop_7_ldst = _RAND_759[5:0];
  _RAND_760 = {1{`RANDOM}};
  rob_uop_7_lrs1 = _RAND_760[5:0];
  _RAND_761 = {1{`RANDOM}};
  rob_uop_7_lrs2 = _RAND_761[5:0];
  _RAND_762 = {1{`RANDOM}};
  rob_uop_7_lrs3 = _RAND_762[5:0];
  _RAND_763 = {1{`RANDOM}};
  rob_uop_7_ldst_val = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  rob_uop_7_dst_rtype = _RAND_764[1:0];
  _RAND_765 = {1{`RANDOM}};
  rob_uop_7_lrs1_rtype = _RAND_765[1:0];
  _RAND_766 = {1{`RANDOM}};
  rob_uop_7_lrs2_rtype = _RAND_766[1:0];
  _RAND_767 = {1{`RANDOM}};
  rob_uop_7_frs3_en = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  rob_uop_7_fp_val = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  rob_uop_7_fp_single = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  rob_uop_7_xcpt_pf_if = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  rob_uop_7_xcpt_ae_if = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  rob_uop_7_xcpt_ma_if = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  rob_uop_7_bp_debug_if = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  rob_uop_7_bp_xcpt_if = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  rob_uop_7_debug_fsrc = _RAND_775[1:0];
  _RAND_776 = {1{`RANDOM}};
  rob_uop_7_debug_tsrc = _RAND_776[1:0];
  _RAND_777 = {1{`RANDOM}};
  rob_uop_8_uopc = _RAND_777[6:0];
  _RAND_778 = {1{`RANDOM}};
  rob_uop_8_inst = _RAND_778[31:0];
  _RAND_779 = {1{`RANDOM}};
  rob_uop_8_debug_inst = _RAND_779[31:0];
  _RAND_780 = {1{`RANDOM}};
  rob_uop_8_is_rvc = _RAND_780[0:0];
  _RAND_781 = {2{`RANDOM}};
  rob_uop_8_debug_pc = _RAND_781[39:0];
  _RAND_782 = {1{`RANDOM}};
  rob_uop_8_iq_type = _RAND_782[2:0];
  _RAND_783 = {1{`RANDOM}};
  rob_uop_8_fu_code = _RAND_783[9:0];
  _RAND_784 = {1{`RANDOM}};
  rob_uop_8_ctrl_br_type = _RAND_784[3:0];
  _RAND_785 = {1{`RANDOM}};
  rob_uop_8_ctrl_op1_sel = _RAND_785[1:0];
  _RAND_786 = {1{`RANDOM}};
  rob_uop_8_ctrl_op2_sel = _RAND_786[2:0];
  _RAND_787 = {1{`RANDOM}};
  rob_uop_8_ctrl_imm_sel = _RAND_787[2:0];
  _RAND_788 = {1{`RANDOM}};
  rob_uop_8_ctrl_op_fcn = _RAND_788[3:0];
  _RAND_789 = {1{`RANDOM}};
  rob_uop_8_ctrl_fcn_dw = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  rob_uop_8_ctrl_csr_cmd = _RAND_790[2:0];
  _RAND_791 = {1{`RANDOM}};
  rob_uop_8_ctrl_is_load = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  rob_uop_8_ctrl_is_sta = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  rob_uop_8_ctrl_is_std = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  rob_uop_8_iw_state = _RAND_794[1:0];
  _RAND_795 = {1{`RANDOM}};
  rob_uop_8_iw_p1_poisoned = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  rob_uop_8_iw_p2_poisoned = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  rob_uop_8_is_br = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  rob_uop_8_is_jalr = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  rob_uop_8_is_jal = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  rob_uop_8_is_sfb = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  rob_uop_8_br_mask = _RAND_801[7:0];
  _RAND_802 = {1{`RANDOM}};
  rob_uop_8_br_tag = _RAND_802[2:0];
  _RAND_803 = {1{`RANDOM}};
  rob_uop_8_ftq_idx = _RAND_803[3:0];
  _RAND_804 = {1{`RANDOM}};
  rob_uop_8_edge_inst = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  rob_uop_8_pc_lob = _RAND_805[5:0];
  _RAND_806 = {1{`RANDOM}};
  rob_uop_8_taken = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  rob_uop_8_imm_packed = _RAND_807[19:0];
  _RAND_808 = {1{`RANDOM}};
  rob_uop_8_csr_addr = _RAND_808[11:0];
  _RAND_809 = {1{`RANDOM}};
  rob_uop_8_rob_idx = _RAND_809[4:0];
  _RAND_810 = {1{`RANDOM}};
  rob_uop_8_ldq_idx = _RAND_810[2:0];
  _RAND_811 = {1{`RANDOM}};
  rob_uop_8_stq_idx = _RAND_811[2:0];
  _RAND_812 = {1{`RANDOM}};
  rob_uop_8_rxq_idx = _RAND_812[1:0];
  _RAND_813 = {1{`RANDOM}};
  rob_uop_8_pdst = _RAND_813[5:0];
  _RAND_814 = {1{`RANDOM}};
  rob_uop_8_prs1 = _RAND_814[5:0];
  _RAND_815 = {1{`RANDOM}};
  rob_uop_8_prs2 = _RAND_815[5:0];
  _RAND_816 = {1{`RANDOM}};
  rob_uop_8_prs3 = _RAND_816[5:0];
  _RAND_817 = {1{`RANDOM}};
  rob_uop_8_ppred = _RAND_817[3:0];
  _RAND_818 = {1{`RANDOM}};
  rob_uop_8_prs1_busy = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  rob_uop_8_prs2_busy = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  rob_uop_8_prs3_busy = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  rob_uop_8_ppred_busy = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  rob_uop_8_stale_pdst = _RAND_822[5:0];
  _RAND_823 = {1{`RANDOM}};
  rob_uop_8_exception = _RAND_823[0:0];
  _RAND_824 = {2{`RANDOM}};
  rob_uop_8_exc_cause = _RAND_824[63:0];
  _RAND_825 = {1{`RANDOM}};
  rob_uop_8_bypassable = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  rob_uop_8_mem_cmd = _RAND_826[4:0];
  _RAND_827 = {1{`RANDOM}};
  rob_uop_8_mem_size = _RAND_827[1:0];
  _RAND_828 = {1{`RANDOM}};
  rob_uop_8_mem_signed = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  rob_uop_8_is_fence = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  rob_uop_8_is_fencei = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  rob_uop_8_is_amo = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  rob_uop_8_uses_ldq = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  rob_uop_8_uses_stq = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  rob_uop_8_is_sys_pc2epc = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  rob_uop_8_is_unique = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  rob_uop_8_flush_on_commit = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  rob_uop_8_ldst_is_rs1 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  rob_uop_8_ldst = _RAND_838[5:0];
  _RAND_839 = {1{`RANDOM}};
  rob_uop_8_lrs1 = _RAND_839[5:0];
  _RAND_840 = {1{`RANDOM}};
  rob_uop_8_lrs2 = _RAND_840[5:0];
  _RAND_841 = {1{`RANDOM}};
  rob_uop_8_lrs3 = _RAND_841[5:0];
  _RAND_842 = {1{`RANDOM}};
  rob_uop_8_ldst_val = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  rob_uop_8_dst_rtype = _RAND_843[1:0];
  _RAND_844 = {1{`RANDOM}};
  rob_uop_8_lrs1_rtype = _RAND_844[1:0];
  _RAND_845 = {1{`RANDOM}};
  rob_uop_8_lrs2_rtype = _RAND_845[1:0];
  _RAND_846 = {1{`RANDOM}};
  rob_uop_8_frs3_en = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  rob_uop_8_fp_val = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  rob_uop_8_fp_single = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  rob_uop_8_xcpt_pf_if = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  rob_uop_8_xcpt_ae_if = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  rob_uop_8_xcpt_ma_if = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  rob_uop_8_bp_debug_if = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  rob_uop_8_bp_xcpt_if = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  rob_uop_8_debug_fsrc = _RAND_854[1:0];
  _RAND_855 = {1{`RANDOM}};
  rob_uop_8_debug_tsrc = _RAND_855[1:0];
  _RAND_856 = {1{`RANDOM}};
  rob_uop_9_uopc = _RAND_856[6:0];
  _RAND_857 = {1{`RANDOM}};
  rob_uop_9_inst = _RAND_857[31:0];
  _RAND_858 = {1{`RANDOM}};
  rob_uop_9_debug_inst = _RAND_858[31:0];
  _RAND_859 = {1{`RANDOM}};
  rob_uop_9_is_rvc = _RAND_859[0:0];
  _RAND_860 = {2{`RANDOM}};
  rob_uop_9_debug_pc = _RAND_860[39:0];
  _RAND_861 = {1{`RANDOM}};
  rob_uop_9_iq_type = _RAND_861[2:0];
  _RAND_862 = {1{`RANDOM}};
  rob_uop_9_fu_code = _RAND_862[9:0];
  _RAND_863 = {1{`RANDOM}};
  rob_uop_9_ctrl_br_type = _RAND_863[3:0];
  _RAND_864 = {1{`RANDOM}};
  rob_uop_9_ctrl_op1_sel = _RAND_864[1:0];
  _RAND_865 = {1{`RANDOM}};
  rob_uop_9_ctrl_op2_sel = _RAND_865[2:0];
  _RAND_866 = {1{`RANDOM}};
  rob_uop_9_ctrl_imm_sel = _RAND_866[2:0];
  _RAND_867 = {1{`RANDOM}};
  rob_uop_9_ctrl_op_fcn = _RAND_867[3:0];
  _RAND_868 = {1{`RANDOM}};
  rob_uop_9_ctrl_fcn_dw = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  rob_uop_9_ctrl_csr_cmd = _RAND_869[2:0];
  _RAND_870 = {1{`RANDOM}};
  rob_uop_9_ctrl_is_load = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  rob_uop_9_ctrl_is_sta = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  rob_uop_9_ctrl_is_std = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  rob_uop_9_iw_state = _RAND_873[1:0];
  _RAND_874 = {1{`RANDOM}};
  rob_uop_9_iw_p1_poisoned = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  rob_uop_9_iw_p2_poisoned = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  rob_uop_9_is_br = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  rob_uop_9_is_jalr = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  rob_uop_9_is_jal = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  rob_uop_9_is_sfb = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  rob_uop_9_br_mask = _RAND_880[7:0];
  _RAND_881 = {1{`RANDOM}};
  rob_uop_9_br_tag = _RAND_881[2:0];
  _RAND_882 = {1{`RANDOM}};
  rob_uop_9_ftq_idx = _RAND_882[3:0];
  _RAND_883 = {1{`RANDOM}};
  rob_uop_9_edge_inst = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  rob_uop_9_pc_lob = _RAND_884[5:0];
  _RAND_885 = {1{`RANDOM}};
  rob_uop_9_taken = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  rob_uop_9_imm_packed = _RAND_886[19:0];
  _RAND_887 = {1{`RANDOM}};
  rob_uop_9_csr_addr = _RAND_887[11:0];
  _RAND_888 = {1{`RANDOM}};
  rob_uop_9_rob_idx = _RAND_888[4:0];
  _RAND_889 = {1{`RANDOM}};
  rob_uop_9_ldq_idx = _RAND_889[2:0];
  _RAND_890 = {1{`RANDOM}};
  rob_uop_9_stq_idx = _RAND_890[2:0];
  _RAND_891 = {1{`RANDOM}};
  rob_uop_9_rxq_idx = _RAND_891[1:0];
  _RAND_892 = {1{`RANDOM}};
  rob_uop_9_pdst = _RAND_892[5:0];
  _RAND_893 = {1{`RANDOM}};
  rob_uop_9_prs1 = _RAND_893[5:0];
  _RAND_894 = {1{`RANDOM}};
  rob_uop_9_prs2 = _RAND_894[5:0];
  _RAND_895 = {1{`RANDOM}};
  rob_uop_9_prs3 = _RAND_895[5:0];
  _RAND_896 = {1{`RANDOM}};
  rob_uop_9_ppred = _RAND_896[3:0];
  _RAND_897 = {1{`RANDOM}};
  rob_uop_9_prs1_busy = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  rob_uop_9_prs2_busy = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  rob_uop_9_prs3_busy = _RAND_899[0:0];
  _RAND_900 = {1{`RANDOM}};
  rob_uop_9_ppred_busy = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  rob_uop_9_stale_pdst = _RAND_901[5:0];
  _RAND_902 = {1{`RANDOM}};
  rob_uop_9_exception = _RAND_902[0:0];
  _RAND_903 = {2{`RANDOM}};
  rob_uop_9_exc_cause = _RAND_903[63:0];
  _RAND_904 = {1{`RANDOM}};
  rob_uop_9_bypassable = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  rob_uop_9_mem_cmd = _RAND_905[4:0];
  _RAND_906 = {1{`RANDOM}};
  rob_uop_9_mem_size = _RAND_906[1:0];
  _RAND_907 = {1{`RANDOM}};
  rob_uop_9_mem_signed = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  rob_uop_9_is_fence = _RAND_908[0:0];
  _RAND_909 = {1{`RANDOM}};
  rob_uop_9_is_fencei = _RAND_909[0:0];
  _RAND_910 = {1{`RANDOM}};
  rob_uop_9_is_amo = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  rob_uop_9_uses_ldq = _RAND_911[0:0];
  _RAND_912 = {1{`RANDOM}};
  rob_uop_9_uses_stq = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  rob_uop_9_is_sys_pc2epc = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  rob_uop_9_is_unique = _RAND_914[0:0];
  _RAND_915 = {1{`RANDOM}};
  rob_uop_9_flush_on_commit = _RAND_915[0:0];
  _RAND_916 = {1{`RANDOM}};
  rob_uop_9_ldst_is_rs1 = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  rob_uop_9_ldst = _RAND_917[5:0];
  _RAND_918 = {1{`RANDOM}};
  rob_uop_9_lrs1 = _RAND_918[5:0];
  _RAND_919 = {1{`RANDOM}};
  rob_uop_9_lrs2 = _RAND_919[5:0];
  _RAND_920 = {1{`RANDOM}};
  rob_uop_9_lrs3 = _RAND_920[5:0];
  _RAND_921 = {1{`RANDOM}};
  rob_uop_9_ldst_val = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  rob_uop_9_dst_rtype = _RAND_922[1:0];
  _RAND_923 = {1{`RANDOM}};
  rob_uop_9_lrs1_rtype = _RAND_923[1:0];
  _RAND_924 = {1{`RANDOM}};
  rob_uop_9_lrs2_rtype = _RAND_924[1:0];
  _RAND_925 = {1{`RANDOM}};
  rob_uop_9_frs3_en = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  rob_uop_9_fp_val = _RAND_926[0:0];
  _RAND_927 = {1{`RANDOM}};
  rob_uop_9_fp_single = _RAND_927[0:0];
  _RAND_928 = {1{`RANDOM}};
  rob_uop_9_xcpt_pf_if = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  rob_uop_9_xcpt_ae_if = _RAND_929[0:0];
  _RAND_930 = {1{`RANDOM}};
  rob_uop_9_xcpt_ma_if = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  rob_uop_9_bp_debug_if = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  rob_uop_9_bp_xcpt_if = _RAND_932[0:0];
  _RAND_933 = {1{`RANDOM}};
  rob_uop_9_debug_fsrc = _RAND_933[1:0];
  _RAND_934 = {1{`RANDOM}};
  rob_uop_9_debug_tsrc = _RAND_934[1:0];
  _RAND_935 = {1{`RANDOM}};
  rob_uop_10_uopc = _RAND_935[6:0];
  _RAND_936 = {1{`RANDOM}};
  rob_uop_10_inst = _RAND_936[31:0];
  _RAND_937 = {1{`RANDOM}};
  rob_uop_10_debug_inst = _RAND_937[31:0];
  _RAND_938 = {1{`RANDOM}};
  rob_uop_10_is_rvc = _RAND_938[0:0];
  _RAND_939 = {2{`RANDOM}};
  rob_uop_10_debug_pc = _RAND_939[39:0];
  _RAND_940 = {1{`RANDOM}};
  rob_uop_10_iq_type = _RAND_940[2:0];
  _RAND_941 = {1{`RANDOM}};
  rob_uop_10_fu_code = _RAND_941[9:0];
  _RAND_942 = {1{`RANDOM}};
  rob_uop_10_ctrl_br_type = _RAND_942[3:0];
  _RAND_943 = {1{`RANDOM}};
  rob_uop_10_ctrl_op1_sel = _RAND_943[1:0];
  _RAND_944 = {1{`RANDOM}};
  rob_uop_10_ctrl_op2_sel = _RAND_944[2:0];
  _RAND_945 = {1{`RANDOM}};
  rob_uop_10_ctrl_imm_sel = _RAND_945[2:0];
  _RAND_946 = {1{`RANDOM}};
  rob_uop_10_ctrl_op_fcn = _RAND_946[3:0];
  _RAND_947 = {1{`RANDOM}};
  rob_uop_10_ctrl_fcn_dw = _RAND_947[0:0];
  _RAND_948 = {1{`RANDOM}};
  rob_uop_10_ctrl_csr_cmd = _RAND_948[2:0];
  _RAND_949 = {1{`RANDOM}};
  rob_uop_10_ctrl_is_load = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  rob_uop_10_ctrl_is_sta = _RAND_950[0:0];
  _RAND_951 = {1{`RANDOM}};
  rob_uop_10_ctrl_is_std = _RAND_951[0:0];
  _RAND_952 = {1{`RANDOM}};
  rob_uop_10_iw_state = _RAND_952[1:0];
  _RAND_953 = {1{`RANDOM}};
  rob_uop_10_iw_p1_poisoned = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  rob_uop_10_iw_p2_poisoned = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  rob_uop_10_is_br = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  rob_uop_10_is_jalr = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  rob_uop_10_is_jal = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  rob_uop_10_is_sfb = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  rob_uop_10_br_mask = _RAND_959[7:0];
  _RAND_960 = {1{`RANDOM}};
  rob_uop_10_br_tag = _RAND_960[2:0];
  _RAND_961 = {1{`RANDOM}};
  rob_uop_10_ftq_idx = _RAND_961[3:0];
  _RAND_962 = {1{`RANDOM}};
  rob_uop_10_edge_inst = _RAND_962[0:0];
  _RAND_963 = {1{`RANDOM}};
  rob_uop_10_pc_lob = _RAND_963[5:0];
  _RAND_964 = {1{`RANDOM}};
  rob_uop_10_taken = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  rob_uop_10_imm_packed = _RAND_965[19:0];
  _RAND_966 = {1{`RANDOM}};
  rob_uop_10_csr_addr = _RAND_966[11:0];
  _RAND_967 = {1{`RANDOM}};
  rob_uop_10_rob_idx = _RAND_967[4:0];
  _RAND_968 = {1{`RANDOM}};
  rob_uop_10_ldq_idx = _RAND_968[2:0];
  _RAND_969 = {1{`RANDOM}};
  rob_uop_10_stq_idx = _RAND_969[2:0];
  _RAND_970 = {1{`RANDOM}};
  rob_uop_10_rxq_idx = _RAND_970[1:0];
  _RAND_971 = {1{`RANDOM}};
  rob_uop_10_pdst = _RAND_971[5:0];
  _RAND_972 = {1{`RANDOM}};
  rob_uop_10_prs1 = _RAND_972[5:0];
  _RAND_973 = {1{`RANDOM}};
  rob_uop_10_prs2 = _RAND_973[5:0];
  _RAND_974 = {1{`RANDOM}};
  rob_uop_10_prs3 = _RAND_974[5:0];
  _RAND_975 = {1{`RANDOM}};
  rob_uop_10_ppred = _RAND_975[3:0];
  _RAND_976 = {1{`RANDOM}};
  rob_uop_10_prs1_busy = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  rob_uop_10_prs2_busy = _RAND_977[0:0];
  _RAND_978 = {1{`RANDOM}};
  rob_uop_10_prs3_busy = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  rob_uop_10_ppred_busy = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  rob_uop_10_stale_pdst = _RAND_980[5:0];
  _RAND_981 = {1{`RANDOM}};
  rob_uop_10_exception = _RAND_981[0:0];
  _RAND_982 = {2{`RANDOM}};
  rob_uop_10_exc_cause = _RAND_982[63:0];
  _RAND_983 = {1{`RANDOM}};
  rob_uop_10_bypassable = _RAND_983[0:0];
  _RAND_984 = {1{`RANDOM}};
  rob_uop_10_mem_cmd = _RAND_984[4:0];
  _RAND_985 = {1{`RANDOM}};
  rob_uop_10_mem_size = _RAND_985[1:0];
  _RAND_986 = {1{`RANDOM}};
  rob_uop_10_mem_signed = _RAND_986[0:0];
  _RAND_987 = {1{`RANDOM}};
  rob_uop_10_is_fence = _RAND_987[0:0];
  _RAND_988 = {1{`RANDOM}};
  rob_uop_10_is_fencei = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  rob_uop_10_is_amo = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  rob_uop_10_uses_ldq = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  rob_uop_10_uses_stq = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  rob_uop_10_is_sys_pc2epc = _RAND_992[0:0];
  _RAND_993 = {1{`RANDOM}};
  rob_uop_10_is_unique = _RAND_993[0:0];
  _RAND_994 = {1{`RANDOM}};
  rob_uop_10_flush_on_commit = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  rob_uop_10_ldst_is_rs1 = _RAND_995[0:0];
  _RAND_996 = {1{`RANDOM}};
  rob_uop_10_ldst = _RAND_996[5:0];
  _RAND_997 = {1{`RANDOM}};
  rob_uop_10_lrs1 = _RAND_997[5:0];
  _RAND_998 = {1{`RANDOM}};
  rob_uop_10_lrs2 = _RAND_998[5:0];
  _RAND_999 = {1{`RANDOM}};
  rob_uop_10_lrs3 = _RAND_999[5:0];
  _RAND_1000 = {1{`RANDOM}};
  rob_uop_10_ldst_val = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  rob_uop_10_dst_rtype = _RAND_1001[1:0];
  _RAND_1002 = {1{`RANDOM}};
  rob_uop_10_lrs1_rtype = _RAND_1002[1:0];
  _RAND_1003 = {1{`RANDOM}};
  rob_uop_10_lrs2_rtype = _RAND_1003[1:0];
  _RAND_1004 = {1{`RANDOM}};
  rob_uop_10_frs3_en = _RAND_1004[0:0];
  _RAND_1005 = {1{`RANDOM}};
  rob_uop_10_fp_val = _RAND_1005[0:0];
  _RAND_1006 = {1{`RANDOM}};
  rob_uop_10_fp_single = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  rob_uop_10_xcpt_pf_if = _RAND_1007[0:0];
  _RAND_1008 = {1{`RANDOM}};
  rob_uop_10_xcpt_ae_if = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  rob_uop_10_xcpt_ma_if = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  rob_uop_10_bp_debug_if = _RAND_1010[0:0];
  _RAND_1011 = {1{`RANDOM}};
  rob_uop_10_bp_xcpt_if = _RAND_1011[0:0];
  _RAND_1012 = {1{`RANDOM}};
  rob_uop_10_debug_fsrc = _RAND_1012[1:0];
  _RAND_1013 = {1{`RANDOM}};
  rob_uop_10_debug_tsrc = _RAND_1013[1:0];
  _RAND_1014 = {1{`RANDOM}};
  rob_uop_11_uopc = _RAND_1014[6:0];
  _RAND_1015 = {1{`RANDOM}};
  rob_uop_11_inst = _RAND_1015[31:0];
  _RAND_1016 = {1{`RANDOM}};
  rob_uop_11_debug_inst = _RAND_1016[31:0];
  _RAND_1017 = {1{`RANDOM}};
  rob_uop_11_is_rvc = _RAND_1017[0:0];
  _RAND_1018 = {2{`RANDOM}};
  rob_uop_11_debug_pc = _RAND_1018[39:0];
  _RAND_1019 = {1{`RANDOM}};
  rob_uop_11_iq_type = _RAND_1019[2:0];
  _RAND_1020 = {1{`RANDOM}};
  rob_uop_11_fu_code = _RAND_1020[9:0];
  _RAND_1021 = {1{`RANDOM}};
  rob_uop_11_ctrl_br_type = _RAND_1021[3:0];
  _RAND_1022 = {1{`RANDOM}};
  rob_uop_11_ctrl_op1_sel = _RAND_1022[1:0];
  _RAND_1023 = {1{`RANDOM}};
  rob_uop_11_ctrl_op2_sel = _RAND_1023[2:0];
  _RAND_1024 = {1{`RANDOM}};
  rob_uop_11_ctrl_imm_sel = _RAND_1024[2:0];
  _RAND_1025 = {1{`RANDOM}};
  rob_uop_11_ctrl_op_fcn = _RAND_1025[3:0];
  _RAND_1026 = {1{`RANDOM}};
  rob_uop_11_ctrl_fcn_dw = _RAND_1026[0:0];
  _RAND_1027 = {1{`RANDOM}};
  rob_uop_11_ctrl_csr_cmd = _RAND_1027[2:0];
  _RAND_1028 = {1{`RANDOM}};
  rob_uop_11_ctrl_is_load = _RAND_1028[0:0];
  _RAND_1029 = {1{`RANDOM}};
  rob_uop_11_ctrl_is_sta = _RAND_1029[0:0];
  _RAND_1030 = {1{`RANDOM}};
  rob_uop_11_ctrl_is_std = _RAND_1030[0:0];
  _RAND_1031 = {1{`RANDOM}};
  rob_uop_11_iw_state = _RAND_1031[1:0];
  _RAND_1032 = {1{`RANDOM}};
  rob_uop_11_iw_p1_poisoned = _RAND_1032[0:0];
  _RAND_1033 = {1{`RANDOM}};
  rob_uop_11_iw_p2_poisoned = _RAND_1033[0:0];
  _RAND_1034 = {1{`RANDOM}};
  rob_uop_11_is_br = _RAND_1034[0:0];
  _RAND_1035 = {1{`RANDOM}};
  rob_uop_11_is_jalr = _RAND_1035[0:0];
  _RAND_1036 = {1{`RANDOM}};
  rob_uop_11_is_jal = _RAND_1036[0:0];
  _RAND_1037 = {1{`RANDOM}};
  rob_uop_11_is_sfb = _RAND_1037[0:0];
  _RAND_1038 = {1{`RANDOM}};
  rob_uop_11_br_mask = _RAND_1038[7:0];
  _RAND_1039 = {1{`RANDOM}};
  rob_uop_11_br_tag = _RAND_1039[2:0];
  _RAND_1040 = {1{`RANDOM}};
  rob_uop_11_ftq_idx = _RAND_1040[3:0];
  _RAND_1041 = {1{`RANDOM}};
  rob_uop_11_edge_inst = _RAND_1041[0:0];
  _RAND_1042 = {1{`RANDOM}};
  rob_uop_11_pc_lob = _RAND_1042[5:0];
  _RAND_1043 = {1{`RANDOM}};
  rob_uop_11_taken = _RAND_1043[0:0];
  _RAND_1044 = {1{`RANDOM}};
  rob_uop_11_imm_packed = _RAND_1044[19:0];
  _RAND_1045 = {1{`RANDOM}};
  rob_uop_11_csr_addr = _RAND_1045[11:0];
  _RAND_1046 = {1{`RANDOM}};
  rob_uop_11_rob_idx = _RAND_1046[4:0];
  _RAND_1047 = {1{`RANDOM}};
  rob_uop_11_ldq_idx = _RAND_1047[2:0];
  _RAND_1048 = {1{`RANDOM}};
  rob_uop_11_stq_idx = _RAND_1048[2:0];
  _RAND_1049 = {1{`RANDOM}};
  rob_uop_11_rxq_idx = _RAND_1049[1:0];
  _RAND_1050 = {1{`RANDOM}};
  rob_uop_11_pdst = _RAND_1050[5:0];
  _RAND_1051 = {1{`RANDOM}};
  rob_uop_11_prs1 = _RAND_1051[5:0];
  _RAND_1052 = {1{`RANDOM}};
  rob_uop_11_prs2 = _RAND_1052[5:0];
  _RAND_1053 = {1{`RANDOM}};
  rob_uop_11_prs3 = _RAND_1053[5:0];
  _RAND_1054 = {1{`RANDOM}};
  rob_uop_11_ppred = _RAND_1054[3:0];
  _RAND_1055 = {1{`RANDOM}};
  rob_uop_11_prs1_busy = _RAND_1055[0:0];
  _RAND_1056 = {1{`RANDOM}};
  rob_uop_11_prs2_busy = _RAND_1056[0:0];
  _RAND_1057 = {1{`RANDOM}};
  rob_uop_11_prs3_busy = _RAND_1057[0:0];
  _RAND_1058 = {1{`RANDOM}};
  rob_uop_11_ppred_busy = _RAND_1058[0:0];
  _RAND_1059 = {1{`RANDOM}};
  rob_uop_11_stale_pdst = _RAND_1059[5:0];
  _RAND_1060 = {1{`RANDOM}};
  rob_uop_11_exception = _RAND_1060[0:0];
  _RAND_1061 = {2{`RANDOM}};
  rob_uop_11_exc_cause = _RAND_1061[63:0];
  _RAND_1062 = {1{`RANDOM}};
  rob_uop_11_bypassable = _RAND_1062[0:0];
  _RAND_1063 = {1{`RANDOM}};
  rob_uop_11_mem_cmd = _RAND_1063[4:0];
  _RAND_1064 = {1{`RANDOM}};
  rob_uop_11_mem_size = _RAND_1064[1:0];
  _RAND_1065 = {1{`RANDOM}};
  rob_uop_11_mem_signed = _RAND_1065[0:0];
  _RAND_1066 = {1{`RANDOM}};
  rob_uop_11_is_fence = _RAND_1066[0:0];
  _RAND_1067 = {1{`RANDOM}};
  rob_uop_11_is_fencei = _RAND_1067[0:0];
  _RAND_1068 = {1{`RANDOM}};
  rob_uop_11_is_amo = _RAND_1068[0:0];
  _RAND_1069 = {1{`RANDOM}};
  rob_uop_11_uses_ldq = _RAND_1069[0:0];
  _RAND_1070 = {1{`RANDOM}};
  rob_uop_11_uses_stq = _RAND_1070[0:0];
  _RAND_1071 = {1{`RANDOM}};
  rob_uop_11_is_sys_pc2epc = _RAND_1071[0:0];
  _RAND_1072 = {1{`RANDOM}};
  rob_uop_11_is_unique = _RAND_1072[0:0];
  _RAND_1073 = {1{`RANDOM}};
  rob_uop_11_flush_on_commit = _RAND_1073[0:0];
  _RAND_1074 = {1{`RANDOM}};
  rob_uop_11_ldst_is_rs1 = _RAND_1074[0:0];
  _RAND_1075 = {1{`RANDOM}};
  rob_uop_11_ldst = _RAND_1075[5:0];
  _RAND_1076 = {1{`RANDOM}};
  rob_uop_11_lrs1 = _RAND_1076[5:0];
  _RAND_1077 = {1{`RANDOM}};
  rob_uop_11_lrs2 = _RAND_1077[5:0];
  _RAND_1078 = {1{`RANDOM}};
  rob_uop_11_lrs3 = _RAND_1078[5:0];
  _RAND_1079 = {1{`RANDOM}};
  rob_uop_11_ldst_val = _RAND_1079[0:0];
  _RAND_1080 = {1{`RANDOM}};
  rob_uop_11_dst_rtype = _RAND_1080[1:0];
  _RAND_1081 = {1{`RANDOM}};
  rob_uop_11_lrs1_rtype = _RAND_1081[1:0];
  _RAND_1082 = {1{`RANDOM}};
  rob_uop_11_lrs2_rtype = _RAND_1082[1:0];
  _RAND_1083 = {1{`RANDOM}};
  rob_uop_11_frs3_en = _RAND_1083[0:0];
  _RAND_1084 = {1{`RANDOM}};
  rob_uop_11_fp_val = _RAND_1084[0:0];
  _RAND_1085 = {1{`RANDOM}};
  rob_uop_11_fp_single = _RAND_1085[0:0];
  _RAND_1086 = {1{`RANDOM}};
  rob_uop_11_xcpt_pf_if = _RAND_1086[0:0];
  _RAND_1087 = {1{`RANDOM}};
  rob_uop_11_xcpt_ae_if = _RAND_1087[0:0];
  _RAND_1088 = {1{`RANDOM}};
  rob_uop_11_xcpt_ma_if = _RAND_1088[0:0];
  _RAND_1089 = {1{`RANDOM}};
  rob_uop_11_bp_debug_if = _RAND_1089[0:0];
  _RAND_1090 = {1{`RANDOM}};
  rob_uop_11_bp_xcpt_if = _RAND_1090[0:0];
  _RAND_1091 = {1{`RANDOM}};
  rob_uop_11_debug_fsrc = _RAND_1091[1:0];
  _RAND_1092 = {1{`RANDOM}};
  rob_uop_11_debug_tsrc = _RAND_1092[1:0];
  _RAND_1093 = {1{`RANDOM}};
  rob_uop_12_uopc = _RAND_1093[6:0];
  _RAND_1094 = {1{`RANDOM}};
  rob_uop_12_inst = _RAND_1094[31:0];
  _RAND_1095 = {1{`RANDOM}};
  rob_uop_12_debug_inst = _RAND_1095[31:0];
  _RAND_1096 = {1{`RANDOM}};
  rob_uop_12_is_rvc = _RAND_1096[0:0];
  _RAND_1097 = {2{`RANDOM}};
  rob_uop_12_debug_pc = _RAND_1097[39:0];
  _RAND_1098 = {1{`RANDOM}};
  rob_uop_12_iq_type = _RAND_1098[2:0];
  _RAND_1099 = {1{`RANDOM}};
  rob_uop_12_fu_code = _RAND_1099[9:0];
  _RAND_1100 = {1{`RANDOM}};
  rob_uop_12_ctrl_br_type = _RAND_1100[3:0];
  _RAND_1101 = {1{`RANDOM}};
  rob_uop_12_ctrl_op1_sel = _RAND_1101[1:0];
  _RAND_1102 = {1{`RANDOM}};
  rob_uop_12_ctrl_op2_sel = _RAND_1102[2:0];
  _RAND_1103 = {1{`RANDOM}};
  rob_uop_12_ctrl_imm_sel = _RAND_1103[2:0];
  _RAND_1104 = {1{`RANDOM}};
  rob_uop_12_ctrl_op_fcn = _RAND_1104[3:0];
  _RAND_1105 = {1{`RANDOM}};
  rob_uop_12_ctrl_fcn_dw = _RAND_1105[0:0];
  _RAND_1106 = {1{`RANDOM}};
  rob_uop_12_ctrl_csr_cmd = _RAND_1106[2:0];
  _RAND_1107 = {1{`RANDOM}};
  rob_uop_12_ctrl_is_load = _RAND_1107[0:0];
  _RAND_1108 = {1{`RANDOM}};
  rob_uop_12_ctrl_is_sta = _RAND_1108[0:0];
  _RAND_1109 = {1{`RANDOM}};
  rob_uop_12_ctrl_is_std = _RAND_1109[0:0];
  _RAND_1110 = {1{`RANDOM}};
  rob_uop_12_iw_state = _RAND_1110[1:0];
  _RAND_1111 = {1{`RANDOM}};
  rob_uop_12_iw_p1_poisoned = _RAND_1111[0:0];
  _RAND_1112 = {1{`RANDOM}};
  rob_uop_12_iw_p2_poisoned = _RAND_1112[0:0];
  _RAND_1113 = {1{`RANDOM}};
  rob_uop_12_is_br = _RAND_1113[0:0];
  _RAND_1114 = {1{`RANDOM}};
  rob_uop_12_is_jalr = _RAND_1114[0:0];
  _RAND_1115 = {1{`RANDOM}};
  rob_uop_12_is_jal = _RAND_1115[0:0];
  _RAND_1116 = {1{`RANDOM}};
  rob_uop_12_is_sfb = _RAND_1116[0:0];
  _RAND_1117 = {1{`RANDOM}};
  rob_uop_12_br_mask = _RAND_1117[7:0];
  _RAND_1118 = {1{`RANDOM}};
  rob_uop_12_br_tag = _RAND_1118[2:0];
  _RAND_1119 = {1{`RANDOM}};
  rob_uop_12_ftq_idx = _RAND_1119[3:0];
  _RAND_1120 = {1{`RANDOM}};
  rob_uop_12_edge_inst = _RAND_1120[0:0];
  _RAND_1121 = {1{`RANDOM}};
  rob_uop_12_pc_lob = _RAND_1121[5:0];
  _RAND_1122 = {1{`RANDOM}};
  rob_uop_12_taken = _RAND_1122[0:0];
  _RAND_1123 = {1{`RANDOM}};
  rob_uop_12_imm_packed = _RAND_1123[19:0];
  _RAND_1124 = {1{`RANDOM}};
  rob_uop_12_csr_addr = _RAND_1124[11:0];
  _RAND_1125 = {1{`RANDOM}};
  rob_uop_12_rob_idx = _RAND_1125[4:0];
  _RAND_1126 = {1{`RANDOM}};
  rob_uop_12_ldq_idx = _RAND_1126[2:0];
  _RAND_1127 = {1{`RANDOM}};
  rob_uop_12_stq_idx = _RAND_1127[2:0];
  _RAND_1128 = {1{`RANDOM}};
  rob_uop_12_rxq_idx = _RAND_1128[1:0];
  _RAND_1129 = {1{`RANDOM}};
  rob_uop_12_pdst = _RAND_1129[5:0];
  _RAND_1130 = {1{`RANDOM}};
  rob_uop_12_prs1 = _RAND_1130[5:0];
  _RAND_1131 = {1{`RANDOM}};
  rob_uop_12_prs2 = _RAND_1131[5:0];
  _RAND_1132 = {1{`RANDOM}};
  rob_uop_12_prs3 = _RAND_1132[5:0];
  _RAND_1133 = {1{`RANDOM}};
  rob_uop_12_ppred = _RAND_1133[3:0];
  _RAND_1134 = {1{`RANDOM}};
  rob_uop_12_prs1_busy = _RAND_1134[0:0];
  _RAND_1135 = {1{`RANDOM}};
  rob_uop_12_prs2_busy = _RAND_1135[0:0];
  _RAND_1136 = {1{`RANDOM}};
  rob_uop_12_prs3_busy = _RAND_1136[0:0];
  _RAND_1137 = {1{`RANDOM}};
  rob_uop_12_ppred_busy = _RAND_1137[0:0];
  _RAND_1138 = {1{`RANDOM}};
  rob_uop_12_stale_pdst = _RAND_1138[5:0];
  _RAND_1139 = {1{`RANDOM}};
  rob_uop_12_exception = _RAND_1139[0:0];
  _RAND_1140 = {2{`RANDOM}};
  rob_uop_12_exc_cause = _RAND_1140[63:0];
  _RAND_1141 = {1{`RANDOM}};
  rob_uop_12_bypassable = _RAND_1141[0:0];
  _RAND_1142 = {1{`RANDOM}};
  rob_uop_12_mem_cmd = _RAND_1142[4:0];
  _RAND_1143 = {1{`RANDOM}};
  rob_uop_12_mem_size = _RAND_1143[1:0];
  _RAND_1144 = {1{`RANDOM}};
  rob_uop_12_mem_signed = _RAND_1144[0:0];
  _RAND_1145 = {1{`RANDOM}};
  rob_uop_12_is_fence = _RAND_1145[0:0];
  _RAND_1146 = {1{`RANDOM}};
  rob_uop_12_is_fencei = _RAND_1146[0:0];
  _RAND_1147 = {1{`RANDOM}};
  rob_uop_12_is_amo = _RAND_1147[0:0];
  _RAND_1148 = {1{`RANDOM}};
  rob_uop_12_uses_ldq = _RAND_1148[0:0];
  _RAND_1149 = {1{`RANDOM}};
  rob_uop_12_uses_stq = _RAND_1149[0:0];
  _RAND_1150 = {1{`RANDOM}};
  rob_uop_12_is_sys_pc2epc = _RAND_1150[0:0];
  _RAND_1151 = {1{`RANDOM}};
  rob_uop_12_is_unique = _RAND_1151[0:0];
  _RAND_1152 = {1{`RANDOM}};
  rob_uop_12_flush_on_commit = _RAND_1152[0:0];
  _RAND_1153 = {1{`RANDOM}};
  rob_uop_12_ldst_is_rs1 = _RAND_1153[0:0];
  _RAND_1154 = {1{`RANDOM}};
  rob_uop_12_ldst = _RAND_1154[5:0];
  _RAND_1155 = {1{`RANDOM}};
  rob_uop_12_lrs1 = _RAND_1155[5:0];
  _RAND_1156 = {1{`RANDOM}};
  rob_uop_12_lrs2 = _RAND_1156[5:0];
  _RAND_1157 = {1{`RANDOM}};
  rob_uop_12_lrs3 = _RAND_1157[5:0];
  _RAND_1158 = {1{`RANDOM}};
  rob_uop_12_ldst_val = _RAND_1158[0:0];
  _RAND_1159 = {1{`RANDOM}};
  rob_uop_12_dst_rtype = _RAND_1159[1:0];
  _RAND_1160 = {1{`RANDOM}};
  rob_uop_12_lrs1_rtype = _RAND_1160[1:0];
  _RAND_1161 = {1{`RANDOM}};
  rob_uop_12_lrs2_rtype = _RAND_1161[1:0];
  _RAND_1162 = {1{`RANDOM}};
  rob_uop_12_frs3_en = _RAND_1162[0:0];
  _RAND_1163 = {1{`RANDOM}};
  rob_uop_12_fp_val = _RAND_1163[0:0];
  _RAND_1164 = {1{`RANDOM}};
  rob_uop_12_fp_single = _RAND_1164[0:0];
  _RAND_1165 = {1{`RANDOM}};
  rob_uop_12_xcpt_pf_if = _RAND_1165[0:0];
  _RAND_1166 = {1{`RANDOM}};
  rob_uop_12_xcpt_ae_if = _RAND_1166[0:0];
  _RAND_1167 = {1{`RANDOM}};
  rob_uop_12_xcpt_ma_if = _RAND_1167[0:0];
  _RAND_1168 = {1{`RANDOM}};
  rob_uop_12_bp_debug_if = _RAND_1168[0:0];
  _RAND_1169 = {1{`RANDOM}};
  rob_uop_12_bp_xcpt_if = _RAND_1169[0:0];
  _RAND_1170 = {1{`RANDOM}};
  rob_uop_12_debug_fsrc = _RAND_1170[1:0];
  _RAND_1171 = {1{`RANDOM}};
  rob_uop_12_debug_tsrc = _RAND_1171[1:0];
  _RAND_1172 = {1{`RANDOM}};
  rob_uop_13_uopc = _RAND_1172[6:0];
  _RAND_1173 = {1{`RANDOM}};
  rob_uop_13_inst = _RAND_1173[31:0];
  _RAND_1174 = {1{`RANDOM}};
  rob_uop_13_debug_inst = _RAND_1174[31:0];
  _RAND_1175 = {1{`RANDOM}};
  rob_uop_13_is_rvc = _RAND_1175[0:0];
  _RAND_1176 = {2{`RANDOM}};
  rob_uop_13_debug_pc = _RAND_1176[39:0];
  _RAND_1177 = {1{`RANDOM}};
  rob_uop_13_iq_type = _RAND_1177[2:0];
  _RAND_1178 = {1{`RANDOM}};
  rob_uop_13_fu_code = _RAND_1178[9:0];
  _RAND_1179 = {1{`RANDOM}};
  rob_uop_13_ctrl_br_type = _RAND_1179[3:0];
  _RAND_1180 = {1{`RANDOM}};
  rob_uop_13_ctrl_op1_sel = _RAND_1180[1:0];
  _RAND_1181 = {1{`RANDOM}};
  rob_uop_13_ctrl_op2_sel = _RAND_1181[2:0];
  _RAND_1182 = {1{`RANDOM}};
  rob_uop_13_ctrl_imm_sel = _RAND_1182[2:0];
  _RAND_1183 = {1{`RANDOM}};
  rob_uop_13_ctrl_op_fcn = _RAND_1183[3:0];
  _RAND_1184 = {1{`RANDOM}};
  rob_uop_13_ctrl_fcn_dw = _RAND_1184[0:0];
  _RAND_1185 = {1{`RANDOM}};
  rob_uop_13_ctrl_csr_cmd = _RAND_1185[2:0];
  _RAND_1186 = {1{`RANDOM}};
  rob_uop_13_ctrl_is_load = _RAND_1186[0:0];
  _RAND_1187 = {1{`RANDOM}};
  rob_uop_13_ctrl_is_sta = _RAND_1187[0:0];
  _RAND_1188 = {1{`RANDOM}};
  rob_uop_13_ctrl_is_std = _RAND_1188[0:0];
  _RAND_1189 = {1{`RANDOM}};
  rob_uop_13_iw_state = _RAND_1189[1:0];
  _RAND_1190 = {1{`RANDOM}};
  rob_uop_13_iw_p1_poisoned = _RAND_1190[0:0];
  _RAND_1191 = {1{`RANDOM}};
  rob_uop_13_iw_p2_poisoned = _RAND_1191[0:0];
  _RAND_1192 = {1{`RANDOM}};
  rob_uop_13_is_br = _RAND_1192[0:0];
  _RAND_1193 = {1{`RANDOM}};
  rob_uop_13_is_jalr = _RAND_1193[0:0];
  _RAND_1194 = {1{`RANDOM}};
  rob_uop_13_is_jal = _RAND_1194[0:0];
  _RAND_1195 = {1{`RANDOM}};
  rob_uop_13_is_sfb = _RAND_1195[0:0];
  _RAND_1196 = {1{`RANDOM}};
  rob_uop_13_br_mask = _RAND_1196[7:0];
  _RAND_1197 = {1{`RANDOM}};
  rob_uop_13_br_tag = _RAND_1197[2:0];
  _RAND_1198 = {1{`RANDOM}};
  rob_uop_13_ftq_idx = _RAND_1198[3:0];
  _RAND_1199 = {1{`RANDOM}};
  rob_uop_13_edge_inst = _RAND_1199[0:0];
  _RAND_1200 = {1{`RANDOM}};
  rob_uop_13_pc_lob = _RAND_1200[5:0];
  _RAND_1201 = {1{`RANDOM}};
  rob_uop_13_taken = _RAND_1201[0:0];
  _RAND_1202 = {1{`RANDOM}};
  rob_uop_13_imm_packed = _RAND_1202[19:0];
  _RAND_1203 = {1{`RANDOM}};
  rob_uop_13_csr_addr = _RAND_1203[11:0];
  _RAND_1204 = {1{`RANDOM}};
  rob_uop_13_rob_idx = _RAND_1204[4:0];
  _RAND_1205 = {1{`RANDOM}};
  rob_uop_13_ldq_idx = _RAND_1205[2:0];
  _RAND_1206 = {1{`RANDOM}};
  rob_uop_13_stq_idx = _RAND_1206[2:0];
  _RAND_1207 = {1{`RANDOM}};
  rob_uop_13_rxq_idx = _RAND_1207[1:0];
  _RAND_1208 = {1{`RANDOM}};
  rob_uop_13_pdst = _RAND_1208[5:0];
  _RAND_1209 = {1{`RANDOM}};
  rob_uop_13_prs1 = _RAND_1209[5:0];
  _RAND_1210 = {1{`RANDOM}};
  rob_uop_13_prs2 = _RAND_1210[5:0];
  _RAND_1211 = {1{`RANDOM}};
  rob_uop_13_prs3 = _RAND_1211[5:0];
  _RAND_1212 = {1{`RANDOM}};
  rob_uop_13_ppred = _RAND_1212[3:0];
  _RAND_1213 = {1{`RANDOM}};
  rob_uop_13_prs1_busy = _RAND_1213[0:0];
  _RAND_1214 = {1{`RANDOM}};
  rob_uop_13_prs2_busy = _RAND_1214[0:0];
  _RAND_1215 = {1{`RANDOM}};
  rob_uop_13_prs3_busy = _RAND_1215[0:0];
  _RAND_1216 = {1{`RANDOM}};
  rob_uop_13_ppred_busy = _RAND_1216[0:0];
  _RAND_1217 = {1{`RANDOM}};
  rob_uop_13_stale_pdst = _RAND_1217[5:0];
  _RAND_1218 = {1{`RANDOM}};
  rob_uop_13_exception = _RAND_1218[0:0];
  _RAND_1219 = {2{`RANDOM}};
  rob_uop_13_exc_cause = _RAND_1219[63:0];
  _RAND_1220 = {1{`RANDOM}};
  rob_uop_13_bypassable = _RAND_1220[0:0];
  _RAND_1221 = {1{`RANDOM}};
  rob_uop_13_mem_cmd = _RAND_1221[4:0];
  _RAND_1222 = {1{`RANDOM}};
  rob_uop_13_mem_size = _RAND_1222[1:0];
  _RAND_1223 = {1{`RANDOM}};
  rob_uop_13_mem_signed = _RAND_1223[0:0];
  _RAND_1224 = {1{`RANDOM}};
  rob_uop_13_is_fence = _RAND_1224[0:0];
  _RAND_1225 = {1{`RANDOM}};
  rob_uop_13_is_fencei = _RAND_1225[0:0];
  _RAND_1226 = {1{`RANDOM}};
  rob_uop_13_is_amo = _RAND_1226[0:0];
  _RAND_1227 = {1{`RANDOM}};
  rob_uop_13_uses_ldq = _RAND_1227[0:0];
  _RAND_1228 = {1{`RANDOM}};
  rob_uop_13_uses_stq = _RAND_1228[0:0];
  _RAND_1229 = {1{`RANDOM}};
  rob_uop_13_is_sys_pc2epc = _RAND_1229[0:0];
  _RAND_1230 = {1{`RANDOM}};
  rob_uop_13_is_unique = _RAND_1230[0:0];
  _RAND_1231 = {1{`RANDOM}};
  rob_uop_13_flush_on_commit = _RAND_1231[0:0];
  _RAND_1232 = {1{`RANDOM}};
  rob_uop_13_ldst_is_rs1 = _RAND_1232[0:0];
  _RAND_1233 = {1{`RANDOM}};
  rob_uop_13_ldst = _RAND_1233[5:0];
  _RAND_1234 = {1{`RANDOM}};
  rob_uop_13_lrs1 = _RAND_1234[5:0];
  _RAND_1235 = {1{`RANDOM}};
  rob_uop_13_lrs2 = _RAND_1235[5:0];
  _RAND_1236 = {1{`RANDOM}};
  rob_uop_13_lrs3 = _RAND_1236[5:0];
  _RAND_1237 = {1{`RANDOM}};
  rob_uop_13_ldst_val = _RAND_1237[0:0];
  _RAND_1238 = {1{`RANDOM}};
  rob_uop_13_dst_rtype = _RAND_1238[1:0];
  _RAND_1239 = {1{`RANDOM}};
  rob_uop_13_lrs1_rtype = _RAND_1239[1:0];
  _RAND_1240 = {1{`RANDOM}};
  rob_uop_13_lrs2_rtype = _RAND_1240[1:0];
  _RAND_1241 = {1{`RANDOM}};
  rob_uop_13_frs3_en = _RAND_1241[0:0];
  _RAND_1242 = {1{`RANDOM}};
  rob_uop_13_fp_val = _RAND_1242[0:0];
  _RAND_1243 = {1{`RANDOM}};
  rob_uop_13_fp_single = _RAND_1243[0:0];
  _RAND_1244 = {1{`RANDOM}};
  rob_uop_13_xcpt_pf_if = _RAND_1244[0:0];
  _RAND_1245 = {1{`RANDOM}};
  rob_uop_13_xcpt_ae_if = _RAND_1245[0:0];
  _RAND_1246 = {1{`RANDOM}};
  rob_uop_13_xcpt_ma_if = _RAND_1246[0:0];
  _RAND_1247 = {1{`RANDOM}};
  rob_uop_13_bp_debug_if = _RAND_1247[0:0];
  _RAND_1248 = {1{`RANDOM}};
  rob_uop_13_bp_xcpt_if = _RAND_1248[0:0];
  _RAND_1249 = {1{`RANDOM}};
  rob_uop_13_debug_fsrc = _RAND_1249[1:0];
  _RAND_1250 = {1{`RANDOM}};
  rob_uop_13_debug_tsrc = _RAND_1250[1:0];
  _RAND_1251 = {1{`RANDOM}};
  rob_uop_14_uopc = _RAND_1251[6:0];
  _RAND_1252 = {1{`RANDOM}};
  rob_uop_14_inst = _RAND_1252[31:0];
  _RAND_1253 = {1{`RANDOM}};
  rob_uop_14_debug_inst = _RAND_1253[31:0];
  _RAND_1254 = {1{`RANDOM}};
  rob_uop_14_is_rvc = _RAND_1254[0:0];
  _RAND_1255 = {2{`RANDOM}};
  rob_uop_14_debug_pc = _RAND_1255[39:0];
  _RAND_1256 = {1{`RANDOM}};
  rob_uop_14_iq_type = _RAND_1256[2:0];
  _RAND_1257 = {1{`RANDOM}};
  rob_uop_14_fu_code = _RAND_1257[9:0];
  _RAND_1258 = {1{`RANDOM}};
  rob_uop_14_ctrl_br_type = _RAND_1258[3:0];
  _RAND_1259 = {1{`RANDOM}};
  rob_uop_14_ctrl_op1_sel = _RAND_1259[1:0];
  _RAND_1260 = {1{`RANDOM}};
  rob_uop_14_ctrl_op2_sel = _RAND_1260[2:0];
  _RAND_1261 = {1{`RANDOM}};
  rob_uop_14_ctrl_imm_sel = _RAND_1261[2:0];
  _RAND_1262 = {1{`RANDOM}};
  rob_uop_14_ctrl_op_fcn = _RAND_1262[3:0];
  _RAND_1263 = {1{`RANDOM}};
  rob_uop_14_ctrl_fcn_dw = _RAND_1263[0:0];
  _RAND_1264 = {1{`RANDOM}};
  rob_uop_14_ctrl_csr_cmd = _RAND_1264[2:0];
  _RAND_1265 = {1{`RANDOM}};
  rob_uop_14_ctrl_is_load = _RAND_1265[0:0];
  _RAND_1266 = {1{`RANDOM}};
  rob_uop_14_ctrl_is_sta = _RAND_1266[0:0];
  _RAND_1267 = {1{`RANDOM}};
  rob_uop_14_ctrl_is_std = _RAND_1267[0:0];
  _RAND_1268 = {1{`RANDOM}};
  rob_uop_14_iw_state = _RAND_1268[1:0];
  _RAND_1269 = {1{`RANDOM}};
  rob_uop_14_iw_p1_poisoned = _RAND_1269[0:0];
  _RAND_1270 = {1{`RANDOM}};
  rob_uop_14_iw_p2_poisoned = _RAND_1270[0:0];
  _RAND_1271 = {1{`RANDOM}};
  rob_uop_14_is_br = _RAND_1271[0:0];
  _RAND_1272 = {1{`RANDOM}};
  rob_uop_14_is_jalr = _RAND_1272[0:0];
  _RAND_1273 = {1{`RANDOM}};
  rob_uop_14_is_jal = _RAND_1273[0:0];
  _RAND_1274 = {1{`RANDOM}};
  rob_uop_14_is_sfb = _RAND_1274[0:0];
  _RAND_1275 = {1{`RANDOM}};
  rob_uop_14_br_mask = _RAND_1275[7:0];
  _RAND_1276 = {1{`RANDOM}};
  rob_uop_14_br_tag = _RAND_1276[2:0];
  _RAND_1277 = {1{`RANDOM}};
  rob_uop_14_ftq_idx = _RAND_1277[3:0];
  _RAND_1278 = {1{`RANDOM}};
  rob_uop_14_edge_inst = _RAND_1278[0:0];
  _RAND_1279 = {1{`RANDOM}};
  rob_uop_14_pc_lob = _RAND_1279[5:0];
  _RAND_1280 = {1{`RANDOM}};
  rob_uop_14_taken = _RAND_1280[0:0];
  _RAND_1281 = {1{`RANDOM}};
  rob_uop_14_imm_packed = _RAND_1281[19:0];
  _RAND_1282 = {1{`RANDOM}};
  rob_uop_14_csr_addr = _RAND_1282[11:0];
  _RAND_1283 = {1{`RANDOM}};
  rob_uop_14_rob_idx = _RAND_1283[4:0];
  _RAND_1284 = {1{`RANDOM}};
  rob_uop_14_ldq_idx = _RAND_1284[2:0];
  _RAND_1285 = {1{`RANDOM}};
  rob_uop_14_stq_idx = _RAND_1285[2:0];
  _RAND_1286 = {1{`RANDOM}};
  rob_uop_14_rxq_idx = _RAND_1286[1:0];
  _RAND_1287 = {1{`RANDOM}};
  rob_uop_14_pdst = _RAND_1287[5:0];
  _RAND_1288 = {1{`RANDOM}};
  rob_uop_14_prs1 = _RAND_1288[5:0];
  _RAND_1289 = {1{`RANDOM}};
  rob_uop_14_prs2 = _RAND_1289[5:0];
  _RAND_1290 = {1{`RANDOM}};
  rob_uop_14_prs3 = _RAND_1290[5:0];
  _RAND_1291 = {1{`RANDOM}};
  rob_uop_14_ppred = _RAND_1291[3:0];
  _RAND_1292 = {1{`RANDOM}};
  rob_uop_14_prs1_busy = _RAND_1292[0:0];
  _RAND_1293 = {1{`RANDOM}};
  rob_uop_14_prs2_busy = _RAND_1293[0:0];
  _RAND_1294 = {1{`RANDOM}};
  rob_uop_14_prs3_busy = _RAND_1294[0:0];
  _RAND_1295 = {1{`RANDOM}};
  rob_uop_14_ppred_busy = _RAND_1295[0:0];
  _RAND_1296 = {1{`RANDOM}};
  rob_uop_14_stale_pdst = _RAND_1296[5:0];
  _RAND_1297 = {1{`RANDOM}};
  rob_uop_14_exception = _RAND_1297[0:0];
  _RAND_1298 = {2{`RANDOM}};
  rob_uop_14_exc_cause = _RAND_1298[63:0];
  _RAND_1299 = {1{`RANDOM}};
  rob_uop_14_bypassable = _RAND_1299[0:0];
  _RAND_1300 = {1{`RANDOM}};
  rob_uop_14_mem_cmd = _RAND_1300[4:0];
  _RAND_1301 = {1{`RANDOM}};
  rob_uop_14_mem_size = _RAND_1301[1:0];
  _RAND_1302 = {1{`RANDOM}};
  rob_uop_14_mem_signed = _RAND_1302[0:0];
  _RAND_1303 = {1{`RANDOM}};
  rob_uop_14_is_fence = _RAND_1303[0:0];
  _RAND_1304 = {1{`RANDOM}};
  rob_uop_14_is_fencei = _RAND_1304[0:0];
  _RAND_1305 = {1{`RANDOM}};
  rob_uop_14_is_amo = _RAND_1305[0:0];
  _RAND_1306 = {1{`RANDOM}};
  rob_uop_14_uses_ldq = _RAND_1306[0:0];
  _RAND_1307 = {1{`RANDOM}};
  rob_uop_14_uses_stq = _RAND_1307[0:0];
  _RAND_1308 = {1{`RANDOM}};
  rob_uop_14_is_sys_pc2epc = _RAND_1308[0:0];
  _RAND_1309 = {1{`RANDOM}};
  rob_uop_14_is_unique = _RAND_1309[0:0];
  _RAND_1310 = {1{`RANDOM}};
  rob_uop_14_flush_on_commit = _RAND_1310[0:0];
  _RAND_1311 = {1{`RANDOM}};
  rob_uop_14_ldst_is_rs1 = _RAND_1311[0:0];
  _RAND_1312 = {1{`RANDOM}};
  rob_uop_14_ldst = _RAND_1312[5:0];
  _RAND_1313 = {1{`RANDOM}};
  rob_uop_14_lrs1 = _RAND_1313[5:0];
  _RAND_1314 = {1{`RANDOM}};
  rob_uop_14_lrs2 = _RAND_1314[5:0];
  _RAND_1315 = {1{`RANDOM}};
  rob_uop_14_lrs3 = _RAND_1315[5:0];
  _RAND_1316 = {1{`RANDOM}};
  rob_uop_14_ldst_val = _RAND_1316[0:0];
  _RAND_1317 = {1{`RANDOM}};
  rob_uop_14_dst_rtype = _RAND_1317[1:0];
  _RAND_1318 = {1{`RANDOM}};
  rob_uop_14_lrs1_rtype = _RAND_1318[1:0];
  _RAND_1319 = {1{`RANDOM}};
  rob_uop_14_lrs2_rtype = _RAND_1319[1:0];
  _RAND_1320 = {1{`RANDOM}};
  rob_uop_14_frs3_en = _RAND_1320[0:0];
  _RAND_1321 = {1{`RANDOM}};
  rob_uop_14_fp_val = _RAND_1321[0:0];
  _RAND_1322 = {1{`RANDOM}};
  rob_uop_14_fp_single = _RAND_1322[0:0];
  _RAND_1323 = {1{`RANDOM}};
  rob_uop_14_xcpt_pf_if = _RAND_1323[0:0];
  _RAND_1324 = {1{`RANDOM}};
  rob_uop_14_xcpt_ae_if = _RAND_1324[0:0];
  _RAND_1325 = {1{`RANDOM}};
  rob_uop_14_xcpt_ma_if = _RAND_1325[0:0];
  _RAND_1326 = {1{`RANDOM}};
  rob_uop_14_bp_debug_if = _RAND_1326[0:0];
  _RAND_1327 = {1{`RANDOM}};
  rob_uop_14_bp_xcpt_if = _RAND_1327[0:0];
  _RAND_1328 = {1{`RANDOM}};
  rob_uop_14_debug_fsrc = _RAND_1328[1:0];
  _RAND_1329 = {1{`RANDOM}};
  rob_uop_14_debug_tsrc = _RAND_1329[1:0];
  _RAND_1330 = {1{`RANDOM}};
  rob_uop_15_uopc = _RAND_1330[6:0];
  _RAND_1331 = {1{`RANDOM}};
  rob_uop_15_inst = _RAND_1331[31:0];
  _RAND_1332 = {1{`RANDOM}};
  rob_uop_15_debug_inst = _RAND_1332[31:0];
  _RAND_1333 = {1{`RANDOM}};
  rob_uop_15_is_rvc = _RAND_1333[0:0];
  _RAND_1334 = {2{`RANDOM}};
  rob_uop_15_debug_pc = _RAND_1334[39:0];
  _RAND_1335 = {1{`RANDOM}};
  rob_uop_15_iq_type = _RAND_1335[2:0];
  _RAND_1336 = {1{`RANDOM}};
  rob_uop_15_fu_code = _RAND_1336[9:0];
  _RAND_1337 = {1{`RANDOM}};
  rob_uop_15_ctrl_br_type = _RAND_1337[3:0];
  _RAND_1338 = {1{`RANDOM}};
  rob_uop_15_ctrl_op1_sel = _RAND_1338[1:0];
  _RAND_1339 = {1{`RANDOM}};
  rob_uop_15_ctrl_op2_sel = _RAND_1339[2:0];
  _RAND_1340 = {1{`RANDOM}};
  rob_uop_15_ctrl_imm_sel = _RAND_1340[2:0];
  _RAND_1341 = {1{`RANDOM}};
  rob_uop_15_ctrl_op_fcn = _RAND_1341[3:0];
  _RAND_1342 = {1{`RANDOM}};
  rob_uop_15_ctrl_fcn_dw = _RAND_1342[0:0];
  _RAND_1343 = {1{`RANDOM}};
  rob_uop_15_ctrl_csr_cmd = _RAND_1343[2:0];
  _RAND_1344 = {1{`RANDOM}};
  rob_uop_15_ctrl_is_load = _RAND_1344[0:0];
  _RAND_1345 = {1{`RANDOM}};
  rob_uop_15_ctrl_is_sta = _RAND_1345[0:0];
  _RAND_1346 = {1{`RANDOM}};
  rob_uop_15_ctrl_is_std = _RAND_1346[0:0];
  _RAND_1347 = {1{`RANDOM}};
  rob_uop_15_iw_state = _RAND_1347[1:0];
  _RAND_1348 = {1{`RANDOM}};
  rob_uop_15_iw_p1_poisoned = _RAND_1348[0:0];
  _RAND_1349 = {1{`RANDOM}};
  rob_uop_15_iw_p2_poisoned = _RAND_1349[0:0];
  _RAND_1350 = {1{`RANDOM}};
  rob_uop_15_is_br = _RAND_1350[0:0];
  _RAND_1351 = {1{`RANDOM}};
  rob_uop_15_is_jalr = _RAND_1351[0:0];
  _RAND_1352 = {1{`RANDOM}};
  rob_uop_15_is_jal = _RAND_1352[0:0];
  _RAND_1353 = {1{`RANDOM}};
  rob_uop_15_is_sfb = _RAND_1353[0:0];
  _RAND_1354 = {1{`RANDOM}};
  rob_uop_15_br_mask = _RAND_1354[7:0];
  _RAND_1355 = {1{`RANDOM}};
  rob_uop_15_br_tag = _RAND_1355[2:0];
  _RAND_1356 = {1{`RANDOM}};
  rob_uop_15_ftq_idx = _RAND_1356[3:0];
  _RAND_1357 = {1{`RANDOM}};
  rob_uop_15_edge_inst = _RAND_1357[0:0];
  _RAND_1358 = {1{`RANDOM}};
  rob_uop_15_pc_lob = _RAND_1358[5:0];
  _RAND_1359 = {1{`RANDOM}};
  rob_uop_15_taken = _RAND_1359[0:0];
  _RAND_1360 = {1{`RANDOM}};
  rob_uop_15_imm_packed = _RAND_1360[19:0];
  _RAND_1361 = {1{`RANDOM}};
  rob_uop_15_csr_addr = _RAND_1361[11:0];
  _RAND_1362 = {1{`RANDOM}};
  rob_uop_15_rob_idx = _RAND_1362[4:0];
  _RAND_1363 = {1{`RANDOM}};
  rob_uop_15_ldq_idx = _RAND_1363[2:0];
  _RAND_1364 = {1{`RANDOM}};
  rob_uop_15_stq_idx = _RAND_1364[2:0];
  _RAND_1365 = {1{`RANDOM}};
  rob_uop_15_rxq_idx = _RAND_1365[1:0];
  _RAND_1366 = {1{`RANDOM}};
  rob_uop_15_pdst = _RAND_1366[5:0];
  _RAND_1367 = {1{`RANDOM}};
  rob_uop_15_prs1 = _RAND_1367[5:0];
  _RAND_1368 = {1{`RANDOM}};
  rob_uop_15_prs2 = _RAND_1368[5:0];
  _RAND_1369 = {1{`RANDOM}};
  rob_uop_15_prs3 = _RAND_1369[5:0];
  _RAND_1370 = {1{`RANDOM}};
  rob_uop_15_ppred = _RAND_1370[3:0];
  _RAND_1371 = {1{`RANDOM}};
  rob_uop_15_prs1_busy = _RAND_1371[0:0];
  _RAND_1372 = {1{`RANDOM}};
  rob_uop_15_prs2_busy = _RAND_1372[0:0];
  _RAND_1373 = {1{`RANDOM}};
  rob_uop_15_prs3_busy = _RAND_1373[0:0];
  _RAND_1374 = {1{`RANDOM}};
  rob_uop_15_ppred_busy = _RAND_1374[0:0];
  _RAND_1375 = {1{`RANDOM}};
  rob_uop_15_stale_pdst = _RAND_1375[5:0];
  _RAND_1376 = {1{`RANDOM}};
  rob_uop_15_exception = _RAND_1376[0:0];
  _RAND_1377 = {2{`RANDOM}};
  rob_uop_15_exc_cause = _RAND_1377[63:0];
  _RAND_1378 = {1{`RANDOM}};
  rob_uop_15_bypassable = _RAND_1378[0:0];
  _RAND_1379 = {1{`RANDOM}};
  rob_uop_15_mem_cmd = _RAND_1379[4:0];
  _RAND_1380 = {1{`RANDOM}};
  rob_uop_15_mem_size = _RAND_1380[1:0];
  _RAND_1381 = {1{`RANDOM}};
  rob_uop_15_mem_signed = _RAND_1381[0:0];
  _RAND_1382 = {1{`RANDOM}};
  rob_uop_15_is_fence = _RAND_1382[0:0];
  _RAND_1383 = {1{`RANDOM}};
  rob_uop_15_is_fencei = _RAND_1383[0:0];
  _RAND_1384 = {1{`RANDOM}};
  rob_uop_15_is_amo = _RAND_1384[0:0];
  _RAND_1385 = {1{`RANDOM}};
  rob_uop_15_uses_ldq = _RAND_1385[0:0];
  _RAND_1386 = {1{`RANDOM}};
  rob_uop_15_uses_stq = _RAND_1386[0:0];
  _RAND_1387 = {1{`RANDOM}};
  rob_uop_15_is_sys_pc2epc = _RAND_1387[0:0];
  _RAND_1388 = {1{`RANDOM}};
  rob_uop_15_is_unique = _RAND_1388[0:0];
  _RAND_1389 = {1{`RANDOM}};
  rob_uop_15_flush_on_commit = _RAND_1389[0:0];
  _RAND_1390 = {1{`RANDOM}};
  rob_uop_15_ldst_is_rs1 = _RAND_1390[0:0];
  _RAND_1391 = {1{`RANDOM}};
  rob_uop_15_ldst = _RAND_1391[5:0];
  _RAND_1392 = {1{`RANDOM}};
  rob_uop_15_lrs1 = _RAND_1392[5:0];
  _RAND_1393 = {1{`RANDOM}};
  rob_uop_15_lrs2 = _RAND_1393[5:0];
  _RAND_1394 = {1{`RANDOM}};
  rob_uop_15_lrs3 = _RAND_1394[5:0];
  _RAND_1395 = {1{`RANDOM}};
  rob_uop_15_ldst_val = _RAND_1395[0:0];
  _RAND_1396 = {1{`RANDOM}};
  rob_uop_15_dst_rtype = _RAND_1396[1:0];
  _RAND_1397 = {1{`RANDOM}};
  rob_uop_15_lrs1_rtype = _RAND_1397[1:0];
  _RAND_1398 = {1{`RANDOM}};
  rob_uop_15_lrs2_rtype = _RAND_1398[1:0];
  _RAND_1399 = {1{`RANDOM}};
  rob_uop_15_frs3_en = _RAND_1399[0:0];
  _RAND_1400 = {1{`RANDOM}};
  rob_uop_15_fp_val = _RAND_1400[0:0];
  _RAND_1401 = {1{`RANDOM}};
  rob_uop_15_fp_single = _RAND_1401[0:0];
  _RAND_1402 = {1{`RANDOM}};
  rob_uop_15_xcpt_pf_if = _RAND_1402[0:0];
  _RAND_1403 = {1{`RANDOM}};
  rob_uop_15_xcpt_ae_if = _RAND_1403[0:0];
  _RAND_1404 = {1{`RANDOM}};
  rob_uop_15_xcpt_ma_if = _RAND_1404[0:0];
  _RAND_1405 = {1{`RANDOM}};
  rob_uop_15_bp_debug_if = _RAND_1405[0:0];
  _RAND_1406 = {1{`RANDOM}};
  rob_uop_15_bp_xcpt_if = _RAND_1406[0:0];
  _RAND_1407 = {1{`RANDOM}};
  rob_uop_15_debug_fsrc = _RAND_1407[1:0];
  _RAND_1408 = {1{`RANDOM}};
  rob_uop_15_debug_tsrc = _RAND_1408[1:0];
  _RAND_1409 = {1{`RANDOM}};
  rob_uop_16_uopc = _RAND_1409[6:0];
  _RAND_1410 = {1{`RANDOM}};
  rob_uop_16_inst = _RAND_1410[31:0];
  _RAND_1411 = {1{`RANDOM}};
  rob_uop_16_debug_inst = _RAND_1411[31:0];
  _RAND_1412 = {1{`RANDOM}};
  rob_uop_16_is_rvc = _RAND_1412[0:0];
  _RAND_1413 = {2{`RANDOM}};
  rob_uop_16_debug_pc = _RAND_1413[39:0];
  _RAND_1414 = {1{`RANDOM}};
  rob_uop_16_iq_type = _RAND_1414[2:0];
  _RAND_1415 = {1{`RANDOM}};
  rob_uop_16_fu_code = _RAND_1415[9:0];
  _RAND_1416 = {1{`RANDOM}};
  rob_uop_16_ctrl_br_type = _RAND_1416[3:0];
  _RAND_1417 = {1{`RANDOM}};
  rob_uop_16_ctrl_op1_sel = _RAND_1417[1:0];
  _RAND_1418 = {1{`RANDOM}};
  rob_uop_16_ctrl_op2_sel = _RAND_1418[2:0];
  _RAND_1419 = {1{`RANDOM}};
  rob_uop_16_ctrl_imm_sel = _RAND_1419[2:0];
  _RAND_1420 = {1{`RANDOM}};
  rob_uop_16_ctrl_op_fcn = _RAND_1420[3:0];
  _RAND_1421 = {1{`RANDOM}};
  rob_uop_16_ctrl_fcn_dw = _RAND_1421[0:0];
  _RAND_1422 = {1{`RANDOM}};
  rob_uop_16_ctrl_csr_cmd = _RAND_1422[2:0];
  _RAND_1423 = {1{`RANDOM}};
  rob_uop_16_ctrl_is_load = _RAND_1423[0:0];
  _RAND_1424 = {1{`RANDOM}};
  rob_uop_16_ctrl_is_sta = _RAND_1424[0:0];
  _RAND_1425 = {1{`RANDOM}};
  rob_uop_16_ctrl_is_std = _RAND_1425[0:0];
  _RAND_1426 = {1{`RANDOM}};
  rob_uop_16_iw_state = _RAND_1426[1:0];
  _RAND_1427 = {1{`RANDOM}};
  rob_uop_16_iw_p1_poisoned = _RAND_1427[0:0];
  _RAND_1428 = {1{`RANDOM}};
  rob_uop_16_iw_p2_poisoned = _RAND_1428[0:0];
  _RAND_1429 = {1{`RANDOM}};
  rob_uop_16_is_br = _RAND_1429[0:0];
  _RAND_1430 = {1{`RANDOM}};
  rob_uop_16_is_jalr = _RAND_1430[0:0];
  _RAND_1431 = {1{`RANDOM}};
  rob_uop_16_is_jal = _RAND_1431[0:0];
  _RAND_1432 = {1{`RANDOM}};
  rob_uop_16_is_sfb = _RAND_1432[0:0];
  _RAND_1433 = {1{`RANDOM}};
  rob_uop_16_br_mask = _RAND_1433[7:0];
  _RAND_1434 = {1{`RANDOM}};
  rob_uop_16_br_tag = _RAND_1434[2:0];
  _RAND_1435 = {1{`RANDOM}};
  rob_uop_16_ftq_idx = _RAND_1435[3:0];
  _RAND_1436 = {1{`RANDOM}};
  rob_uop_16_edge_inst = _RAND_1436[0:0];
  _RAND_1437 = {1{`RANDOM}};
  rob_uop_16_pc_lob = _RAND_1437[5:0];
  _RAND_1438 = {1{`RANDOM}};
  rob_uop_16_taken = _RAND_1438[0:0];
  _RAND_1439 = {1{`RANDOM}};
  rob_uop_16_imm_packed = _RAND_1439[19:0];
  _RAND_1440 = {1{`RANDOM}};
  rob_uop_16_csr_addr = _RAND_1440[11:0];
  _RAND_1441 = {1{`RANDOM}};
  rob_uop_16_rob_idx = _RAND_1441[4:0];
  _RAND_1442 = {1{`RANDOM}};
  rob_uop_16_ldq_idx = _RAND_1442[2:0];
  _RAND_1443 = {1{`RANDOM}};
  rob_uop_16_stq_idx = _RAND_1443[2:0];
  _RAND_1444 = {1{`RANDOM}};
  rob_uop_16_rxq_idx = _RAND_1444[1:0];
  _RAND_1445 = {1{`RANDOM}};
  rob_uop_16_pdst = _RAND_1445[5:0];
  _RAND_1446 = {1{`RANDOM}};
  rob_uop_16_prs1 = _RAND_1446[5:0];
  _RAND_1447 = {1{`RANDOM}};
  rob_uop_16_prs2 = _RAND_1447[5:0];
  _RAND_1448 = {1{`RANDOM}};
  rob_uop_16_prs3 = _RAND_1448[5:0];
  _RAND_1449 = {1{`RANDOM}};
  rob_uop_16_ppred = _RAND_1449[3:0];
  _RAND_1450 = {1{`RANDOM}};
  rob_uop_16_prs1_busy = _RAND_1450[0:0];
  _RAND_1451 = {1{`RANDOM}};
  rob_uop_16_prs2_busy = _RAND_1451[0:0];
  _RAND_1452 = {1{`RANDOM}};
  rob_uop_16_prs3_busy = _RAND_1452[0:0];
  _RAND_1453 = {1{`RANDOM}};
  rob_uop_16_ppred_busy = _RAND_1453[0:0];
  _RAND_1454 = {1{`RANDOM}};
  rob_uop_16_stale_pdst = _RAND_1454[5:0];
  _RAND_1455 = {1{`RANDOM}};
  rob_uop_16_exception = _RAND_1455[0:0];
  _RAND_1456 = {2{`RANDOM}};
  rob_uop_16_exc_cause = _RAND_1456[63:0];
  _RAND_1457 = {1{`RANDOM}};
  rob_uop_16_bypassable = _RAND_1457[0:0];
  _RAND_1458 = {1{`RANDOM}};
  rob_uop_16_mem_cmd = _RAND_1458[4:0];
  _RAND_1459 = {1{`RANDOM}};
  rob_uop_16_mem_size = _RAND_1459[1:0];
  _RAND_1460 = {1{`RANDOM}};
  rob_uop_16_mem_signed = _RAND_1460[0:0];
  _RAND_1461 = {1{`RANDOM}};
  rob_uop_16_is_fence = _RAND_1461[0:0];
  _RAND_1462 = {1{`RANDOM}};
  rob_uop_16_is_fencei = _RAND_1462[0:0];
  _RAND_1463 = {1{`RANDOM}};
  rob_uop_16_is_amo = _RAND_1463[0:0];
  _RAND_1464 = {1{`RANDOM}};
  rob_uop_16_uses_ldq = _RAND_1464[0:0];
  _RAND_1465 = {1{`RANDOM}};
  rob_uop_16_uses_stq = _RAND_1465[0:0];
  _RAND_1466 = {1{`RANDOM}};
  rob_uop_16_is_sys_pc2epc = _RAND_1466[0:0];
  _RAND_1467 = {1{`RANDOM}};
  rob_uop_16_is_unique = _RAND_1467[0:0];
  _RAND_1468 = {1{`RANDOM}};
  rob_uop_16_flush_on_commit = _RAND_1468[0:0];
  _RAND_1469 = {1{`RANDOM}};
  rob_uop_16_ldst_is_rs1 = _RAND_1469[0:0];
  _RAND_1470 = {1{`RANDOM}};
  rob_uop_16_ldst = _RAND_1470[5:0];
  _RAND_1471 = {1{`RANDOM}};
  rob_uop_16_lrs1 = _RAND_1471[5:0];
  _RAND_1472 = {1{`RANDOM}};
  rob_uop_16_lrs2 = _RAND_1472[5:0];
  _RAND_1473 = {1{`RANDOM}};
  rob_uop_16_lrs3 = _RAND_1473[5:0];
  _RAND_1474 = {1{`RANDOM}};
  rob_uop_16_ldst_val = _RAND_1474[0:0];
  _RAND_1475 = {1{`RANDOM}};
  rob_uop_16_dst_rtype = _RAND_1475[1:0];
  _RAND_1476 = {1{`RANDOM}};
  rob_uop_16_lrs1_rtype = _RAND_1476[1:0];
  _RAND_1477 = {1{`RANDOM}};
  rob_uop_16_lrs2_rtype = _RAND_1477[1:0];
  _RAND_1478 = {1{`RANDOM}};
  rob_uop_16_frs3_en = _RAND_1478[0:0];
  _RAND_1479 = {1{`RANDOM}};
  rob_uop_16_fp_val = _RAND_1479[0:0];
  _RAND_1480 = {1{`RANDOM}};
  rob_uop_16_fp_single = _RAND_1480[0:0];
  _RAND_1481 = {1{`RANDOM}};
  rob_uop_16_xcpt_pf_if = _RAND_1481[0:0];
  _RAND_1482 = {1{`RANDOM}};
  rob_uop_16_xcpt_ae_if = _RAND_1482[0:0];
  _RAND_1483 = {1{`RANDOM}};
  rob_uop_16_xcpt_ma_if = _RAND_1483[0:0];
  _RAND_1484 = {1{`RANDOM}};
  rob_uop_16_bp_debug_if = _RAND_1484[0:0];
  _RAND_1485 = {1{`RANDOM}};
  rob_uop_16_bp_xcpt_if = _RAND_1485[0:0];
  _RAND_1486 = {1{`RANDOM}};
  rob_uop_16_debug_fsrc = _RAND_1486[1:0];
  _RAND_1487 = {1{`RANDOM}};
  rob_uop_16_debug_tsrc = _RAND_1487[1:0];
  _RAND_1488 = {1{`RANDOM}};
  rob_uop_17_uopc = _RAND_1488[6:0];
  _RAND_1489 = {1{`RANDOM}};
  rob_uop_17_inst = _RAND_1489[31:0];
  _RAND_1490 = {1{`RANDOM}};
  rob_uop_17_debug_inst = _RAND_1490[31:0];
  _RAND_1491 = {1{`RANDOM}};
  rob_uop_17_is_rvc = _RAND_1491[0:0];
  _RAND_1492 = {2{`RANDOM}};
  rob_uop_17_debug_pc = _RAND_1492[39:0];
  _RAND_1493 = {1{`RANDOM}};
  rob_uop_17_iq_type = _RAND_1493[2:0];
  _RAND_1494 = {1{`RANDOM}};
  rob_uop_17_fu_code = _RAND_1494[9:0];
  _RAND_1495 = {1{`RANDOM}};
  rob_uop_17_ctrl_br_type = _RAND_1495[3:0];
  _RAND_1496 = {1{`RANDOM}};
  rob_uop_17_ctrl_op1_sel = _RAND_1496[1:0];
  _RAND_1497 = {1{`RANDOM}};
  rob_uop_17_ctrl_op2_sel = _RAND_1497[2:0];
  _RAND_1498 = {1{`RANDOM}};
  rob_uop_17_ctrl_imm_sel = _RAND_1498[2:0];
  _RAND_1499 = {1{`RANDOM}};
  rob_uop_17_ctrl_op_fcn = _RAND_1499[3:0];
  _RAND_1500 = {1{`RANDOM}};
  rob_uop_17_ctrl_fcn_dw = _RAND_1500[0:0];
  _RAND_1501 = {1{`RANDOM}};
  rob_uop_17_ctrl_csr_cmd = _RAND_1501[2:0];
  _RAND_1502 = {1{`RANDOM}};
  rob_uop_17_ctrl_is_load = _RAND_1502[0:0];
  _RAND_1503 = {1{`RANDOM}};
  rob_uop_17_ctrl_is_sta = _RAND_1503[0:0];
  _RAND_1504 = {1{`RANDOM}};
  rob_uop_17_ctrl_is_std = _RAND_1504[0:0];
  _RAND_1505 = {1{`RANDOM}};
  rob_uop_17_iw_state = _RAND_1505[1:0];
  _RAND_1506 = {1{`RANDOM}};
  rob_uop_17_iw_p1_poisoned = _RAND_1506[0:0];
  _RAND_1507 = {1{`RANDOM}};
  rob_uop_17_iw_p2_poisoned = _RAND_1507[0:0];
  _RAND_1508 = {1{`RANDOM}};
  rob_uop_17_is_br = _RAND_1508[0:0];
  _RAND_1509 = {1{`RANDOM}};
  rob_uop_17_is_jalr = _RAND_1509[0:0];
  _RAND_1510 = {1{`RANDOM}};
  rob_uop_17_is_jal = _RAND_1510[0:0];
  _RAND_1511 = {1{`RANDOM}};
  rob_uop_17_is_sfb = _RAND_1511[0:0];
  _RAND_1512 = {1{`RANDOM}};
  rob_uop_17_br_mask = _RAND_1512[7:0];
  _RAND_1513 = {1{`RANDOM}};
  rob_uop_17_br_tag = _RAND_1513[2:0];
  _RAND_1514 = {1{`RANDOM}};
  rob_uop_17_ftq_idx = _RAND_1514[3:0];
  _RAND_1515 = {1{`RANDOM}};
  rob_uop_17_edge_inst = _RAND_1515[0:0];
  _RAND_1516 = {1{`RANDOM}};
  rob_uop_17_pc_lob = _RAND_1516[5:0];
  _RAND_1517 = {1{`RANDOM}};
  rob_uop_17_taken = _RAND_1517[0:0];
  _RAND_1518 = {1{`RANDOM}};
  rob_uop_17_imm_packed = _RAND_1518[19:0];
  _RAND_1519 = {1{`RANDOM}};
  rob_uop_17_csr_addr = _RAND_1519[11:0];
  _RAND_1520 = {1{`RANDOM}};
  rob_uop_17_rob_idx = _RAND_1520[4:0];
  _RAND_1521 = {1{`RANDOM}};
  rob_uop_17_ldq_idx = _RAND_1521[2:0];
  _RAND_1522 = {1{`RANDOM}};
  rob_uop_17_stq_idx = _RAND_1522[2:0];
  _RAND_1523 = {1{`RANDOM}};
  rob_uop_17_rxq_idx = _RAND_1523[1:0];
  _RAND_1524 = {1{`RANDOM}};
  rob_uop_17_pdst = _RAND_1524[5:0];
  _RAND_1525 = {1{`RANDOM}};
  rob_uop_17_prs1 = _RAND_1525[5:0];
  _RAND_1526 = {1{`RANDOM}};
  rob_uop_17_prs2 = _RAND_1526[5:0];
  _RAND_1527 = {1{`RANDOM}};
  rob_uop_17_prs3 = _RAND_1527[5:0];
  _RAND_1528 = {1{`RANDOM}};
  rob_uop_17_ppred = _RAND_1528[3:0];
  _RAND_1529 = {1{`RANDOM}};
  rob_uop_17_prs1_busy = _RAND_1529[0:0];
  _RAND_1530 = {1{`RANDOM}};
  rob_uop_17_prs2_busy = _RAND_1530[0:0];
  _RAND_1531 = {1{`RANDOM}};
  rob_uop_17_prs3_busy = _RAND_1531[0:0];
  _RAND_1532 = {1{`RANDOM}};
  rob_uop_17_ppred_busy = _RAND_1532[0:0];
  _RAND_1533 = {1{`RANDOM}};
  rob_uop_17_stale_pdst = _RAND_1533[5:0];
  _RAND_1534 = {1{`RANDOM}};
  rob_uop_17_exception = _RAND_1534[0:0];
  _RAND_1535 = {2{`RANDOM}};
  rob_uop_17_exc_cause = _RAND_1535[63:0];
  _RAND_1536 = {1{`RANDOM}};
  rob_uop_17_bypassable = _RAND_1536[0:0];
  _RAND_1537 = {1{`RANDOM}};
  rob_uop_17_mem_cmd = _RAND_1537[4:0];
  _RAND_1538 = {1{`RANDOM}};
  rob_uop_17_mem_size = _RAND_1538[1:0];
  _RAND_1539 = {1{`RANDOM}};
  rob_uop_17_mem_signed = _RAND_1539[0:0];
  _RAND_1540 = {1{`RANDOM}};
  rob_uop_17_is_fence = _RAND_1540[0:0];
  _RAND_1541 = {1{`RANDOM}};
  rob_uop_17_is_fencei = _RAND_1541[0:0];
  _RAND_1542 = {1{`RANDOM}};
  rob_uop_17_is_amo = _RAND_1542[0:0];
  _RAND_1543 = {1{`RANDOM}};
  rob_uop_17_uses_ldq = _RAND_1543[0:0];
  _RAND_1544 = {1{`RANDOM}};
  rob_uop_17_uses_stq = _RAND_1544[0:0];
  _RAND_1545 = {1{`RANDOM}};
  rob_uop_17_is_sys_pc2epc = _RAND_1545[0:0];
  _RAND_1546 = {1{`RANDOM}};
  rob_uop_17_is_unique = _RAND_1546[0:0];
  _RAND_1547 = {1{`RANDOM}};
  rob_uop_17_flush_on_commit = _RAND_1547[0:0];
  _RAND_1548 = {1{`RANDOM}};
  rob_uop_17_ldst_is_rs1 = _RAND_1548[0:0];
  _RAND_1549 = {1{`RANDOM}};
  rob_uop_17_ldst = _RAND_1549[5:0];
  _RAND_1550 = {1{`RANDOM}};
  rob_uop_17_lrs1 = _RAND_1550[5:0];
  _RAND_1551 = {1{`RANDOM}};
  rob_uop_17_lrs2 = _RAND_1551[5:0];
  _RAND_1552 = {1{`RANDOM}};
  rob_uop_17_lrs3 = _RAND_1552[5:0];
  _RAND_1553 = {1{`RANDOM}};
  rob_uop_17_ldst_val = _RAND_1553[0:0];
  _RAND_1554 = {1{`RANDOM}};
  rob_uop_17_dst_rtype = _RAND_1554[1:0];
  _RAND_1555 = {1{`RANDOM}};
  rob_uop_17_lrs1_rtype = _RAND_1555[1:0];
  _RAND_1556 = {1{`RANDOM}};
  rob_uop_17_lrs2_rtype = _RAND_1556[1:0];
  _RAND_1557 = {1{`RANDOM}};
  rob_uop_17_frs3_en = _RAND_1557[0:0];
  _RAND_1558 = {1{`RANDOM}};
  rob_uop_17_fp_val = _RAND_1558[0:0];
  _RAND_1559 = {1{`RANDOM}};
  rob_uop_17_fp_single = _RAND_1559[0:0];
  _RAND_1560 = {1{`RANDOM}};
  rob_uop_17_xcpt_pf_if = _RAND_1560[0:0];
  _RAND_1561 = {1{`RANDOM}};
  rob_uop_17_xcpt_ae_if = _RAND_1561[0:0];
  _RAND_1562 = {1{`RANDOM}};
  rob_uop_17_xcpt_ma_if = _RAND_1562[0:0];
  _RAND_1563 = {1{`RANDOM}};
  rob_uop_17_bp_debug_if = _RAND_1563[0:0];
  _RAND_1564 = {1{`RANDOM}};
  rob_uop_17_bp_xcpt_if = _RAND_1564[0:0];
  _RAND_1565 = {1{`RANDOM}};
  rob_uop_17_debug_fsrc = _RAND_1565[1:0];
  _RAND_1566 = {1{`RANDOM}};
  rob_uop_17_debug_tsrc = _RAND_1566[1:0];
  _RAND_1567 = {1{`RANDOM}};
  rob_uop_18_uopc = _RAND_1567[6:0];
  _RAND_1568 = {1{`RANDOM}};
  rob_uop_18_inst = _RAND_1568[31:0];
  _RAND_1569 = {1{`RANDOM}};
  rob_uop_18_debug_inst = _RAND_1569[31:0];
  _RAND_1570 = {1{`RANDOM}};
  rob_uop_18_is_rvc = _RAND_1570[0:0];
  _RAND_1571 = {2{`RANDOM}};
  rob_uop_18_debug_pc = _RAND_1571[39:0];
  _RAND_1572 = {1{`RANDOM}};
  rob_uop_18_iq_type = _RAND_1572[2:0];
  _RAND_1573 = {1{`RANDOM}};
  rob_uop_18_fu_code = _RAND_1573[9:0];
  _RAND_1574 = {1{`RANDOM}};
  rob_uop_18_ctrl_br_type = _RAND_1574[3:0];
  _RAND_1575 = {1{`RANDOM}};
  rob_uop_18_ctrl_op1_sel = _RAND_1575[1:0];
  _RAND_1576 = {1{`RANDOM}};
  rob_uop_18_ctrl_op2_sel = _RAND_1576[2:0];
  _RAND_1577 = {1{`RANDOM}};
  rob_uop_18_ctrl_imm_sel = _RAND_1577[2:0];
  _RAND_1578 = {1{`RANDOM}};
  rob_uop_18_ctrl_op_fcn = _RAND_1578[3:0];
  _RAND_1579 = {1{`RANDOM}};
  rob_uop_18_ctrl_fcn_dw = _RAND_1579[0:0];
  _RAND_1580 = {1{`RANDOM}};
  rob_uop_18_ctrl_csr_cmd = _RAND_1580[2:0];
  _RAND_1581 = {1{`RANDOM}};
  rob_uop_18_ctrl_is_load = _RAND_1581[0:0];
  _RAND_1582 = {1{`RANDOM}};
  rob_uop_18_ctrl_is_sta = _RAND_1582[0:0];
  _RAND_1583 = {1{`RANDOM}};
  rob_uop_18_ctrl_is_std = _RAND_1583[0:0];
  _RAND_1584 = {1{`RANDOM}};
  rob_uop_18_iw_state = _RAND_1584[1:0];
  _RAND_1585 = {1{`RANDOM}};
  rob_uop_18_iw_p1_poisoned = _RAND_1585[0:0];
  _RAND_1586 = {1{`RANDOM}};
  rob_uop_18_iw_p2_poisoned = _RAND_1586[0:0];
  _RAND_1587 = {1{`RANDOM}};
  rob_uop_18_is_br = _RAND_1587[0:0];
  _RAND_1588 = {1{`RANDOM}};
  rob_uop_18_is_jalr = _RAND_1588[0:0];
  _RAND_1589 = {1{`RANDOM}};
  rob_uop_18_is_jal = _RAND_1589[0:0];
  _RAND_1590 = {1{`RANDOM}};
  rob_uop_18_is_sfb = _RAND_1590[0:0];
  _RAND_1591 = {1{`RANDOM}};
  rob_uop_18_br_mask = _RAND_1591[7:0];
  _RAND_1592 = {1{`RANDOM}};
  rob_uop_18_br_tag = _RAND_1592[2:0];
  _RAND_1593 = {1{`RANDOM}};
  rob_uop_18_ftq_idx = _RAND_1593[3:0];
  _RAND_1594 = {1{`RANDOM}};
  rob_uop_18_edge_inst = _RAND_1594[0:0];
  _RAND_1595 = {1{`RANDOM}};
  rob_uop_18_pc_lob = _RAND_1595[5:0];
  _RAND_1596 = {1{`RANDOM}};
  rob_uop_18_taken = _RAND_1596[0:0];
  _RAND_1597 = {1{`RANDOM}};
  rob_uop_18_imm_packed = _RAND_1597[19:0];
  _RAND_1598 = {1{`RANDOM}};
  rob_uop_18_csr_addr = _RAND_1598[11:0];
  _RAND_1599 = {1{`RANDOM}};
  rob_uop_18_rob_idx = _RAND_1599[4:0];
  _RAND_1600 = {1{`RANDOM}};
  rob_uop_18_ldq_idx = _RAND_1600[2:0];
  _RAND_1601 = {1{`RANDOM}};
  rob_uop_18_stq_idx = _RAND_1601[2:0];
  _RAND_1602 = {1{`RANDOM}};
  rob_uop_18_rxq_idx = _RAND_1602[1:0];
  _RAND_1603 = {1{`RANDOM}};
  rob_uop_18_pdst = _RAND_1603[5:0];
  _RAND_1604 = {1{`RANDOM}};
  rob_uop_18_prs1 = _RAND_1604[5:0];
  _RAND_1605 = {1{`RANDOM}};
  rob_uop_18_prs2 = _RAND_1605[5:0];
  _RAND_1606 = {1{`RANDOM}};
  rob_uop_18_prs3 = _RAND_1606[5:0];
  _RAND_1607 = {1{`RANDOM}};
  rob_uop_18_ppred = _RAND_1607[3:0];
  _RAND_1608 = {1{`RANDOM}};
  rob_uop_18_prs1_busy = _RAND_1608[0:0];
  _RAND_1609 = {1{`RANDOM}};
  rob_uop_18_prs2_busy = _RAND_1609[0:0];
  _RAND_1610 = {1{`RANDOM}};
  rob_uop_18_prs3_busy = _RAND_1610[0:0];
  _RAND_1611 = {1{`RANDOM}};
  rob_uop_18_ppred_busy = _RAND_1611[0:0];
  _RAND_1612 = {1{`RANDOM}};
  rob_uop_18_stale_pdst = _RAND_1612[5:0];
  _RAND_1613 = {1{`RANDOM}};
  rob_uop_18_exception = _RAND_1613[0:0];
  _RAND_1614 = {2{`RANDOM}};
  rob_uop_18_exc_cause = _RAND_1614[63:0];
  _RAND_1615 = {1{`RANDOM}};
  rob_uop_18_bypassable = _RAND_1615[0:0];
  _RAND_1616 = {1{`RANDOM}};
  rob_uop_18_mem_cmd = _RAND_1616[4:0];
  _RAND_1617 = {1{`RANDOM}};
  rob_uop_18_mem_size = _RAND_1617[1:0];
  _RAND_1618 = {1{`RANDOM}};
  rob_uop_18_mem_signed = _RAND_1618[0:0];
  _RAND_1619 = {1{`RANDOM}};
  rob_uop_18_is_fence = _RAND_1619[0:0];
  _RAND_1620 = {1{`RANDOM}};
  rob_uop_18_is_fencei = _RAND_1620[0:0];
  _RAND_1621 = {1{`RANDOM}};
  rob_uop_18_is_amo = _RAND_1621[0:0];
  _RAND_1622 = {1{`RANDOM}};
  rob_uop_18_uses_ldq = _RAND_1622[0:0];
  _RAND_1623 = {1{`RANDOM}};
  rob_uop_18_uses_stq = _RAND_1623[0:0];
  _RAND_1624 = {1{`RANDOM}};
  rob_uop_18_is_sys_pc2epc = _RAND_1624[0:0];
  _RAND_1625 = {1{`RANDOM}};
  rob_uop_18_is_unique = _RAND_1625[0:0];
  _RAND_1626 = {1{`RANDOM}};
  rob_uop_18_flush_on_commit = _RAND_1626[0:0];
  _RAND_1627 = {1{`RANDOM}};
  rob_uop_18_ldst_is_rs1 = _RAND_1627[0:0];
  _RAND_1628 = {1{`RANDOM}};
  rob_uop_18_ldst = _RAND_1628[5:0];
  _RAND_1629 = {1{`RANDOM}};
  rob_uop_18_lrs1 = _RAND_1629[5:0];
  _RAND_1630 = {1{`RANDOM}};
  rob_uop_18_lrs2 = _RAND_1630[5:0];
  _RAND_1631 = {1{`RANDOM}};
  rob_uop_18_lrs3 = _RAND_1631[5:0];
  _RAND_1632 = {1{`RANDOM}};
  rob_uop_18_ldst_val = _RAND_1632[0:0];
  _RAND_1633 = {1{`RANDOM}};
  rob_uop_18_dst_rtype = _RAND_1633[1:0];
  _RAND_1634 = {1{`RANDOM}};
  rob_uop_18_lrs1_rtype = _RAND_1634[1:0];
  _RAND_1635 = {1{`RANDOM}};
  rob_uop_18_lrs2_rtype = _RAND_1635[1:0];
  _RAND_1636 = {1{`RANDOM}};
  rob_uop_18_frs3_en = _RAND_1636[0:0];
  _RAND_1637 = {1{`RANDOM}};
  rob_uop_18_fp_val = _RAND_1637[0:0];
  _RAND_1638 = {1{`RANDOM}};
  rob_uop_18_fp_single = _RAND_1638[0:0];
  _RAND_1639 = {1{`RANDOM}};
  rob_uop_18_xcpt_pf_if = _RAND_1639[0:0];
  _RAND_1640 = {1{`RANDOM}};
  rob_uop_18_xcpt_ae_if = _RAND_1640[0:0];
  _RAND_1641 = {1{`RANDOM}};
  rob_uop_18_xcpt_ma_if = _RAND_1641[0:0];
  _RAND_1642 = {1{`RANDOM}};
  rob_uop_18_bp_debug_if = _RAND_1642[0:0];
  _RAND_1643 = {1{`RANDOM}};
  rob_uop_18_bp_xcpt_if = _RAND_1643[0:0];
  _RAND_1644 = {1{`RANDOM}};
  rob_uop_18_debug_fsrc = _RAND_1644[1:0];
  _RAND_1645 = {1{`RANDOM}};
  rob_uop_18_debug_tsrc = _RAND_1645[1:0];
  _RAND_1646 = {1{`RANDOM}};
  rob_uop_19_uopc = _RAND_1646[6:0];
  _RAND_1647 = {1{`RANDOM}};
  rob_uop_19_inst = _RAND_1647[31:0];
  _RAND_1648 = {1{`RANDOM}};
  rob_uop_19_debug_inst = _RAND_1648[31:0];
  _RAND_1649 = {1{`RANDOM}};
  rob_uop_19_is_rvc = _RAND_1649[0:0];
  _RAND_1650 = {2{`RANDOM}};
  rob_uop_19_debug_pc = _RAND_1650[39:0];
  _RAND_1651 = {1{`RANDOM}};
  rob_uop_19_iq_type = _RAND_1651[2:0];
  _RAND_1652 = {1{`RANDOM}};
  rob_uop_19_fu_code = _RAND_1652[9:0];
  _RAND_1653 = {1{`RANDOM}};
  rob_uop_19_ctrl_br_type = _RAND_1653[3:0];
  _RAND_1654 = {1{`RANDOM}};
  rob_uop_19_ctrl_op1_sel = _RAND_1654[1:0];
  _RAND_1655 = {1{`RANDOM}};
  rob_uop_19_ctrl_op2_sel = _RAND_1655[2:0];
  _RAND_1656 = {1{`RANDOM}};
  rob_uop_19_ctrl_imm_sel = _RAND_1656[2:0];
  _RAND_1657 = {1{`RANDOM}};
  rob_uop_19_ctrl_op_fcn = _RAND_1657[3:0];
  _RAND_1658 = {1{`RANDOM}};
  rob_uop_19_ctrl_fcn_dw = _RAND_1658[0:0];
  _RAND_1659 = {1{`RANDOM}};
  rob_uop_19_ctrl_csr_cmd = _RAND_1659[2:0];
  _RAND_1660 = {1{`RANDOM}};
  rob_uop_19_ctrl_is_load = _RAND_1660[0:0];
  _RAND_1661 = {1{`RANDOM}};
  rob_uop_19_ctrl_is_sta = _RAND_1661[0:0];
  _RAND_1662 = {1{`RANDOM}};
  rob_uop_19_ctrl_is_std = _RAND_1662[0:0];
  _RAND_1663 = {1{`RANDOM}};
  rob_uop_19_iw_state = _RAND_1663[1:0];
  _RAND_1664 = {1{`RANDOM}};
  rob_uop_19_iw_p1_poisoned = _RAND_1664[0:0];
  _RAND_1665 = {1{`RANDOM}};
  rob_uop_19_iw_p2_poisoned = _RAND_1665[0:0];
  _RAND_1666 = {1{`RANDOM}};
  rob_uop_19_is_br = _RAND_1666[0:0];
  _RAND_1667 = {1{`RANDOM}};
  rob_uop_19_is_jalr = _RAND_1667[0:0];
  _RAND_1668 = {1{`RANDOM}};
  rob_uop_19_is_jal = _RAND_1668[0:0];
  _RAND_1669 = {1{`RANDOM}};
  rob_uop_19_is_sfb = _RAND_1669[0:0];
  _RAND_1670 = {1{`RANDOM}};
  rob_uop_19_br_mask = _RAND_1670[7:0];
  _RAND_1671 = {1{`RANDOM}};
  rob_uop_19_br_tag = _RAND_1671[2:0];
  _RAND_1672 = {1{`RANDOM}};
  rob_uop_19_ftq_idx = _RAND_1672[3:0];
  _RAND_1673 = {1{`RANDOM}};
  rob_uop_19_edge_inst = _RAND_1673[0:0];
  _RAND_1674 = {1{`RANDOM}};
  rob_uop_19_pc_lob = _RAND_1674[5:0];
  _RAND_1675 = {1{`RANDOM}};
  rob_uop_19_taken = _RAND_1675[0:0];
  _RAND_1676 = {1{`RANDOM}};
  rob_uop_19_imm_packed = _RAND_1676[19:0];
  _RAND_1677 = {1{`RANDOM}};
  rob_uop_19_csr_addr = _RAND_1677[11:0];
  _RAND_1678 = {1{`RANDOM}};
  rob_uop_19_rob_idx = _RAND_1678[4:0];
  _RAND_1679 = {1{`RANDOM}};
  rob_uop_19_ldq_idx = _RAND_1679[2:0];
  _RAND_1680 = {1{`RANDOM}};
  rob_uop_19_stq_idx = _RAND_1680[2:0];
  _RAND_1681 = {1{`RANDOM}};
  rob_uop_19_rxq_idx = _RAND_1681[1:0];
  _RAND_1682 = {1{`RANDOM}};
  rob_uop_19_pdst = _RAND_1682[5:0];
  _RAND_1683 = {1{`RANDOM}};
  rob_uop_19_prs1 = _RAND_1683[5:0];
  _RAND_1684 = {1{`RANDOM}};
  rob_uop_19_prs2 = _RAND_1684[5:0];
  _RAND_1685 = {1{`RANDOM}};
  rob_uop_19_prs3 = _RAND_1685[5:0];
  _RAND_1686 = {1{`RANDOM}};
  rob_uop_19_ppred = _RAND_1686[3:0];
  _RAND_1687 = {1{`RANDOM}};
  rob_uop_19_prs1_busy = _RAND_1687[0:0];
  _RAND_1688 = {1{`RANDOM}};
  rob_uop_19_prs2_busy = _RAND_1688[0:0];
  _RAND_1689 = {1{`RANDOM}};
  rob_uop_19_prs3_busy = _RAND_1689[0:0];
  _RAND_1690 = {1{`RANDOM}};
  rob_uop_19_ppred_busy = _RAND_1690[0:0];
  _RAND_1691 = {1{`RANDOM}};
  rob_uop_19_stale_pdst = _RAND_1691[5:0];
  _RAND_1692 = {1{`RANDOM}};
  rob_uop_19_exception = _RAND_1692[0:0];
  _RAND_1693 = {2{`RANDOM}};
  rob_uop_19_exc_cause = _RAND_1693[63:0];
  _RAND_1694 = {1{`RANDOM}};
  rob_uop_19_bypassable = _RAND_1694[0:0];
  _RAND_1695 = {1{`RANDOM}};
  rob_uop_19_mem_cmd = _RAND_1695[4:0];
  _RAND_1696 = {1{`RANDOM}};
  rob_uop_19_mem_size = _RAND_1696[1:0];
  _RAND_1697 = {1{`RANDOM}};
  rob_uop_19_mem_signed = _RAND_1697[0:0];
  _RAND_1698 = {1{`RANDOM}};
  rob_uop_19_is_fence = _RAND_1698[0:0];
  _RAND_1699 = {1{`RANDOM}};
  rob_uop_19_is_fencei = _RAND_1699[0:0];
  _RAND_1700 = {1{`RANDOM}};
  rob_uop_19_is_amo = _RAND_1700[0:0];
  _RAND_1701 = {1{`RANDOM}};
  rob_uop_19_uses_ldq = _RAND_1701[0:0];
  _RAND_1702 = {1{`RANDOM}};
  rob_uop_19_uses_stq = _RAND_1702[0:0];
  _RAND_1703 = {1{`RANDOM}};
  rob_uop_19_is_sys_pc2epc = _RAND_1703[0:0];
  _RAND_1704 = {1{`RANDOM}};
  rob_uop_19_is_unique = _RAND_1704[0:0];
  _RAND_1705 = {1{`RANDOM}};
  rob_uop_19_flush_on_commit = _RAND_1705[0:0];
  _RAND_1706 = {1{`RANDOM}};
  rob_uop_19_ldst_is_rs1 = _RAND_1706[0:0];
  _RAND_1707 = {1{`RANDOM}};
  rob_uop_19_ldst = _RAND_1707[5:0];
  _RAND_1708 = {1{`RANDOM}};
  rob_uop_19_lrs1 = _RAND_1708[5:0];
  _RAND_1709 = {1{`RANDOM}};
  rob_uop_19_lrs2 = _RAND_1709[5:0];
  _RAND_1710 = {1{`RANDOM}};
  rob_uop_19_lrs3 = _RAND_1710[5:0];
  _RAND_1711 = {1{`RANDOM}};
  rob_uop_19_ldst_val = _RAND_1711[0:0];
  _RAND_1712 = {1{`RANDOM}};
  rob_uop_19_dst_rtype = _RAND_1712[1:0];
  _RAND_1713 = {1{`RANDOM}};
  rob_uop_19_lrs1_rtype = _RAND_1713[1:0];
  _RAND_1714 = {1{`RANDOM}};
  rob_uop_19_lrs2_rtype = _RAND_1714[1:0];
  _RAND_1715 = {1{`RANDOM}};
  rob_uop_19_frs3_en = _RAND_1715[0:0];
  _RAND_1716 = {1{`RANDOM}};
  rob_uop_19_fp_val = _RAND_1716[0:0];
  _RAND_1717 = {1{`RANDOM}};
  rob_uop_19_fp_single = _RAND_1717[0:0];
  _RAND_1718 = {1{`RANDOM}};
  rob_uop_19_xcpt_pf_if = _RAND_1718[0:0];
  _RAND_1719 = {1{`RANDOM}};
  rob_uop_19_xcpt_ae_if = _RAND_1719[0:0];
  _RAND_1720 = {1{`RANDOM}};
  rob_uop_19_xcpt_ma_if = _RAND_1720[0:0];
  _RAND_1721 = {1{`RANDOM}};
  rob_uop_19_bp_debug_if = _RAND_1721[0:0];
  _RAND_1722 = {1{`RANDOM}};
  rob_uop_19_bp_xcpt_if = _RAND_1722[0:0];
  _RAND_1723 = {1{`RANDOM}};
  rob_uop_19_debug_fsrc = _RAND_1723[1:0];
  _RAND_1724 = {1{`RANDOM}};
  rob_uop_19_debug_tsrc = _RAND_1724[1:0];
  _RAND_1725 = {1{`RANDOM}};
  rob_uop_20_uopc = _RAND_1725[6:0];
  _RAND_1726 = {1{`RANDOM}};
  rob_uop_20_inst = _RAND_1726[31:0];
  _RAND_1727 = {1{`RANDOM}};
  rob_uop_20_debug_inst = _RAND_1727[31:0];
  _RAND_1728 = {1{`RANDOM}};
  rob_uop_20_is_rvc = _RAND_1728[0:0];
  _RAND_1729 = {2{`RANDOM}};
  rob_uop_20_debug_pc = _RAND_1729[39:0];
  _RAND_1730 = {1{`RANDOM}};
  rob_uop_20_iq_type = _RAND_1730[2:0];
  _RAND_1731 = {1{`RANDOM}};
  rob_uop_20_fu_code = _RAND_1731[9:0];
  _RAND_1732 = {1{`RANDOM}};
  rob_uop_20_ctrl_br_type = _RAND_1732[3:0];
  _RAND_1733 = {1{`RANDOM}};
  rob_uop_20_ctrl_op1_sel = _RAND_1733[1:0];
  _RAND_1734 = {1{`RANDOM}};
  rob_uop_20_ctrl_op2_sel = _RAND_1734[2:0];
  _RAND_1735 = {1{`RANDOM}};
  rob_uop_20_ctrl_imm_sel = _RAND_1735[2:0];
  _RAND_1736 = {1{`RANDOM}};
  rob_uop_20_ctrl_op_fcn = _RAND_1736[3:0];
  _RAND_1737 = {1{`RANDOM}};
  rob_uop_20_ctrl_fcn_dw = _RAND_1737[0:0];
  _RAND_1738 = {1{`RANDOM}};
  rob_uop_20_ctrl_csr_cmd = _RAND_1738[2:0];
  _RAND_1739 = {1{`RANDOM}};
  rob_uop_20_ctrl_is_load = _RAND_1739[0:0];
  _RAND_1740 = {1{`RANDOM}};
  rob_uop_20_ctrl_is_sta = _RAND_1740[0:0];
  _RAND_1741 = {1{`RANDOM}};
  rob_uop_20_ctrl_is_std = _RAND_1741[0:0];
  _RAND_1742 = {1{`RANDOM}};
  rob_uop_20_iw_state = _RAND_1742[1:0];
  _RAND_1743 = {1{`RANDOM}};
  rob_uop_20_iw_p1_poisoned = _RAND_1743[0:0];
  _RAND_1744 = {1{`RANDOM}};
  rob_uop_20_iw_p2_poisoned = _RAND_1744[0:0];
  _RAND_1745 = {1{`RANDOM}};
  rob_uop_20_is_br = _RAND_1745[0:0];
  _RAND_1746 = {1{`RANDOM}};
  rob_uop_20_is_jalr = _RAND_1746[0:0];
  _RAND_1747 = {1{`RANDOM}};
  rob_uop_20_is_jal = _RAND_1747[0:0];
  _RAND_1748 = {1{`RANDOM}};
  rob_uop_20_is_sfb = _RAND_1748[0:0];
  _RAND_1749 = {1{`RANDOM}};
  rob_uop_20_br_mask = _RAND_1749[7:0];
  _RAND_1750 = {1{`RANDOM}};
  rob_uop_20_br_tag = _RAND_1750[2:0];
  _RAND_1751 = {1{`RANDOM}};
  rob_uop_20_ftq_idx = _RAND_1751[3:0];
  _RAND_1752 = {1{`RANDOM}};
  rob_uop_20_edge_inst = _RAND_1752[0:0];
  _RAND_1753 = {1{`RANDOM}};
  rob_uop_20_pc_lob = _RAND_1753[5:0];
  _RAND_1754 = {1{`RANDOM}};
  rob_uop_20_taken = _RAND_1754[0:0];
  _RAND_1755 = {1{`RANDOM}};
  rob_uop_20_imm_packed = _RAND_1755[19:0];
  _RAND_1756 = {1{`RANDOM}};
  rob_uop_20_csr_addr = _RAND_1756[11:0];
  _RAND_1757 = {1{`RANDOM}};
  rob_uop_20_rob_idx = _RAND_1757[4:0];
  _RAND_1758 = {1{`RANDOM}};
  rob_uop_20_ldq_idx = _RAND_1758[2:0];
  _RAND_1759 = {1{`RANDOM}};
  rob_uop_20_stq_idx = _RAND_1759[2:0];
  _RAND_1760 = {1{`RANDOM}};
  rob_uop_20_rxq_idx = _RAND_1760[1:0];
  _RAND_1761 = {1{`RANDOM}};
  rob_uop_20_pdst = _RAND_1761[5:0];
  _RAND_1762 = {1{`RANDOM}};
  rob_uop_20_prs1 = _RAND_1762[5:0];
  _RAND_1763 = {1{`RANDOM}};
  rob_uop_20_prs2 = _RAND_1763[5:0];
  _RAND_1764 = {1{`RANDOM}};
  rob_uop_20_prs3 = _RAND_1764[5:0];
  _RAND_1765 = {1{`RANDOM}};
  rob_uop_20_ppred = _RAND_1765[3:0];
  _RAND_1766 = {1{`RANDOM}};
  rob_uop_20_prs1_busy = _RAND_1766[0:0];
  _RAND_1767 = {1{`RANDOM}};
  rob_uop_20_prs2_busy = _RAND_1767[0:0];
  _RAND_1768 = {1{`RANDOM}};
  rob_uop_20_prs3_busy = _RAND_1768[0:0];
  _RAND_1769 = {1{`RANDOM}};
  rob_uop_20_ppred_busy = _RAND_1769[0:0];
  _RAND_1770 = {1{`RANDOM}};
  rob_uop_20_stale_pdst = _RAND_1770[5:0];
  _RAND_1771 = {1{`RANDOM}};
  rob_uop_20_exception = _RAND_1771[0:0];
  _RAND_1772 = {2{`RANDOM}};
  rob_uop_20_exc_cause = _RAND_1772[63:0];
  _RAND_1773 = {1{`RANDOM}};
  rob_uop_20_bypassable = _RAND_1773[0:0];
  _RAND_1774 = {1{`RANDOM}};
  rob_uop_20_mem_cmd = _RAND_1774[4:0];
  _RAND_1775 = {1{`RANDOM}};
  rob_uop_20_mem_size = _RAND_1775[1:0];
  _RAND_1776 = {1{`RANDOM}};
  rob_uop_20_mem_signed = _RAND_1776[0:0];
  _RAND_1777 = {1{`RANDOM}};
  rob_uop_20_is_fence = _RAND_1777[0:0];
  _RAND_1778 = {1{`RANDOM}};
  rob_uop_20_is_fencei = _RAND_1778[0:0];
  _RAND_1779 = {1{`RANDOM}};
  rob_uop_20_is_amo = _RAND_1779[0:0];
  _RAND_1780 = {1{`RANDOM}};
  rob_uop_20_uses_ldq = _RAND_1780[0:0];
  _RAND_1781 = {1{`RANDOM}};
  rob_uop_20_uses_stq = _RAND_1781[0:0];
  _RAND_1782 = {1{`RANDOM}};
  rob_uop_20_is_sys_pc2epc = _RAND_1782[0:0];
  _RAND_1783 = {1{`RANDOM}};
  rob_uop_20_is_unique = _RAND_1783[0:0];
  _RAND_1784 = {1{`RANDOM}};
  rob_uop_20_flush_on_commit = _RAND_1784[0:0];
  _RAND_1785 = {1{`RANDOM}};
  rob_uop_20_ldst_is_rs1 = _RAND_1785[0:0];
  _RAND_1786 = {1{`RANDOM}};
  rob_uop_20_ldst = _RAND_1786[5:0];
  _RAND_1787 = {1{`RANDOM}};
  rob_uop_20_lrs1 = _RAND_1787[5:0];
  _RAND_1788 = {1{`RANDOM}};
  rob_uop_20_lrs2 = _RAND_1788[5:0];
  _RAND_1789 = {1{`RANDOM}};
  rob_uop_20_lrs3 = _RAND_1789[5:0];
  _RAND_1790 = {1{`RANDOM}};
  rob_uop_20_ldst_val = _RAND_1790[0:0];
  _RAND_1791 = {1{`RANDOM}};
  rob_uop_20_dst_rtype = _RAND_1791[1:0];
  _RAND_1792 = {1{`RANDOM}};
  rob_uop_20_lrs1_rtype = _RAND_1792[1:0];
  _RAND_1793 = {1{`RANDOM}};
  rob_uop_20_lrs2_rtype = _RAND_1793[1:0];
  _RAND_1794 = {1{`RANDOM}};
  rob_uop_20_frs3_en = _RAND_1794[0:0];
  _RAND_1795 = {1{`RANDOM}};
  rob_uop_20_fp_val = _RAND_1795[0:0];
  _RAND_1796 = {1{`RANDOM}};
  rob_uop_20_fp_single = _RAND_1796[0:0];
  _RAND_1797 = {1{`RANDOM}};
  rob_uop_20_xcpt_pf_if = _RAND_1797[0:0];
  _RAND_1798 = {1{`RANDOM}};
  rob_uop_20_xcpt_ae_if = _RAND_1798[0:0];
  _RAND_1799 = {1{`RANDOM}};
  rob_uop_20_xcpt_ma_if = _RAND_1799[0:0];
  _RAND_1800 = {1{`RANDOM}};
  rob_uop_20_bp_debug_if = _RAND_1800[0:0];
  _RAND_1801 = {1{`RANDOM}};
  rob_uop_20_bp_xcpt_if = _RAND_1801[0:0];
  _RAND_1802 = {1{`RANDOM}};
  rob_uop_20_debug_fsrc = _RAND_1802[1:0];
  _RAND_1803 = {1{`RANDOM}};
  rob_uop_20_debug_tsrc = _RAND_1803[1:0];
  _RAND_1804 = {1{`RANDOM}};
  rob_uop_21_uopc = _RAND_1804[6:0];
  _RAND_1805 = {1{`RANDOM}};
  rob_uop_21_inst = _RAND_1805[31:0];
  _RAND_1806 = {1{`RANDOM}};
  rob_uop_21_debug_inst = _RAND_1806[31:0];
  _RAND_1807 = {1{`RANDOM}};
  rob_uop_21_is_rvc = _RAND_1807[0:0];
  _RAND_1808 = {2{`RANDOM}};
  rob_uop_21_debug_pc = _RAND_1808[39:0];
  _RAND_1809 = {1{`RANDOM}};
  rob_uop_21_iq_type = _RAND_1809[2:0];
  _RAND_1810 = {1{`RANDOM}};
  rob_uop_21_fu_code = _RAND_1810[9:0];
  _RAND_1811 = {1{`RANDOM}};
  rob_uop_21_ctrl_br_type = _RAND_1811[3:0];
  _RAND_1812 = {1{`RANDOM}};
  rob_uop_21_ctrl_op1_sel = _RAND_1812[1:0];
  _RAND_1813 = {1{`RANDOM}};
  rob_uop_21_ctrl_op2_sel = _RAND_1813[2:0];
  _RAND_1814 = {1{`RANDOM}};
  rob_uop_21_ctrl_imm_sel = _RAND_1814[2:0];
  _RAND_1815 = {1{`RANDOM}};
  rob_uop_21_ctrl_op_fcn = _RAND_1815[3:0];
  _RAND_1816 = {1{`RANDOM}};
  rob_uop_21_ctrl_fcn_dw = _RAND_1816[0:0];
  _RAND_1817 = {1{`RANDOM}};
  rob_uop_21_ctrl_csr_cmd = _RAND_1817[2:0];
  _RAND_1818 = {1{`RANDOM}};
  rob_uop_21_ctrl_is_load = _RAND_1818[0:0];
  _RAND_1819 = {1{`RANDOM}};
  rob_uop_21_ctrl_is_sta = _RAND_1819[0:0];
  _RAND_1820 = {1{`RANDOM}};
  rob_uop_21_ctrl_is_std = _RAND_1820[0:0];
  _RAND_1821 = {1{`RANDOM}};
  rob_uop_21_iw_state = _RAND_1821[1:0];
  _RAND_1822 = {1{`RANDOM}};
  rob_uop_21_iw_p1_poisoned = _RAND_1822[0:0];
  _RAND_1823 = {1{`RANDOM}};
  rob_uop_21_iw_p2_poisoned = _RAND_1823[0:0];
  _RAND_1824 = {1{`RANDOM}};
  rob_uop_21_is_br = _RAND_1824[0:0];
  _RAND_1825 = {1{`RANDOM}};
  rob_uop_21_is_jalr = _RAND_1825[0:0];
  _RAND_1826 = {1{`RANDOM}};
  rob_uop_21_is_jal = _RAND_1826[0:0];
  _RAND_1827 = {1{`RANDOM}};
  rob_uop_21_is_sfb = _RAND_1827[0:0];
  _RAND_1828 = {1{`RANDOM}};
  rob_uop_21_br_mask = _RAND_1828[7:0];
  _RAND_1829 = {1{`RANDOM}};
  rob_uop_21_br_tag = _RAND_1829[2:0];
  _RAND_1830 = {1{`RANDOM}};
  rob_uop_21_ftq_idx = _RAND_1830[3:0];
  _RAND_1831 = {1{`RANDOM}};
  rob_uop_21_edge_inst = _RAND_1831[0:0];
  _RAND_1832 = {1{`RANDOM}};
  rob_uop_21_pc_lob = _RAND_1832[5:0];
  _RAND_1833 = {1{`RANDOM}};
  rob_uop_21_taken = _RAND_1833[0:0];
  _RAND_1834 = {1{`RANDOM}};
  rob_uop_21_imm_packed = _RAND_1834[19:0];
  _RAND_1835 = {1{`RANDOM}};
  rob_uop_21_csr_addr = _RAND_1835[11:0];
  _RAND_1836 = {1{`RANDOM}};
  rob_uop_21_rob_idx = _RAND_1836[4:0];
  _RAND_1837 = {1{`RANDOM}};
  rob_uop_21_ldq_idx = _RAND_1837[2:0];
  _RAND_1838 = {1{`RANDOM}};
  rob_uop_21_stq_idx = _RAND_1838[2:0];
  _RAND_1839 = {1{`RANDOM}};
  rob_uop_21_rxq_idx = _RAND_1839[1:0];
  _RAND_1840 = {1{`RANDOM}};
  rob_uop_21_pdst = _RAND_1840[5:0];
  _RAND_1841 = {1{`RANDOM}};
  rob_uop_21_prs1 = _RAND_1841[5:0];
  _RAND_1842 = {1{`RANDOM}};
  rob_uop_21_prs2 = _RAND_1842[5:0];
  _RAND_1843 = {1{`RANDOM}};
  rob_uop_21_prs3 = _RAND_1843[5:0];
  _RAND_1844 = {1{`RANDOM}};
  rob_uop_21_ppred = _RAND_1844[3:0];
  _RAND_1845 = {1{`RANDOM}};
  rob_uop_21_prs1_busy = _RAND_1845[0:0];
  _RAND_1846 = {1{`RANDOM}};
  rob_uop_21_prs2_busy = _RAND_1846[0:0];
  _RAND_1847 = {1{`RANDOM}};
  rob_uop_21_prs3_busy = _RAND_1847[0:0];
  _RAND_1848 = {1{`RANDOM}};
  rob_uop_21_ppred_busy = _RAND_1848[0:0];
  _RAND_1849 = {1{`RANDOM}};
  rob_uop_21_stale_pdst = _RAND_1849[5:0];
  _RAND_1850 = {1{`RANDOM}};
  rob_uop_21_exception = _RAND_1850[0:0];
  _RAND_1851 = {2{`RANDOM}};
  rob_uop_21_exc_cause = _RAND_1851[63:0];
  _RAND_1852 = {1{`RANDOM}};
  rob_uop_21_bypassable = _RAND_1852[0:0];
  _RAND_1853 = {1{`RANDOM}};
  rob_uop_21_mem_cmd = _RAND_1853[4:0];
  _RAND_1854 = {1{`RANDOM}};
  rob_uop_21_mem_size = _RAND_1854[1:0];
  _RAND_1855 = {1{`RANDOM}};
  rob_uop_21_mem_signed = _RAND_1855[0:0];
  _RAND_1856 = {1{`RANDOM}};
  rob_uop_21_is_fence = _RAND_1856[0:0];
  _RAND_1857 = {1{`RANDOM}};
  rob_uop_21_is_fencei = _RAND_1857[0:0];
  _RAND_1858 = {1{`RANDOM}};
  rob_uop_21_is_amo = _RAND_1858[0:0];
  _RAND_1859 = {1{`RANDOM}};
  rob_uop_21_uses_ldq = _RAND_1859[0:0];
  _RAND_1860 = {1{`RANDOM}};
  rob_uop_21_uses_stq = _RAND_1860[0:0];
  _RAND_1861 = {1{`RANDOM}};
  rob_uop_21_is_sys_pc2epc = _RAND_1861[0:0];
  _RAND_1862 = {1{`RANDOM}};
  rob_uop_21_is_unique = _RAND_1862[0:0];
  _RAND_1863 = {1{`RANDOM}};
  rob_uop_21_flush_on_commit = _RAND_1863[0:0];
  _RAND_1864 = {1{`RANDOM}};
  rob_uop_21_ldst_is_rs1 = _RAND_1864[0:0];
  _RAND_1865 = {1{`RANDOM}};
  rob_uop_21_ldst = _RAND_1865[5:0];
  _RAND_1866 = {1{`RANDOM}};
  rob_uop_21_lrs1 = _RAND_1866[5:0];
  _RAND_1867 = {1{`RANDOM}};
  rob_uop_21_lrs2 = _RAND_1867[5:0];
  _RAND_1868 = {1{`RANDOM}};
  rob_uop_21_lrs3 = _RAND_1868[5:0];
  _RAND_1869 = {1{`RANDOM}};
  rob_uop_21_ldst_val = _RAND_1869[0:0];
  _RAND_1870 = {1{`RANDOM}};
  rob_uop_21_dst_rtype = _RAND_1870[1:0];
  _RAND_1871 = {1{`RANDOM}};
  rob_uop_21_lrs1_rtype = _RAND_1871[1:0];
  _RAND_1872 = {1{`RANDOM}};
  rob_uop_21_lrs2_rtype = _RAND_1872[1:0];
  _RAND_1873 = {1{`RANDOM}};
  rob_uop_21_frs3_en = _RAND_1873[0:0];
  _RAND_1874 = {1{`RANDOM}};
  rob_uop_21_fp_val = _RAND_1874[0:0];
  _RAND_1875 = {1{`RANDOM}};
  rob_uop_21_fp_single = _RAND_1875[0:0];
  _RAND_1876 = {1{`RANDOM}};
  rob_uop_21_xcpt_pf_if = _RAND_1876[0:0];
  _RAND_1877 = {1{`RANDOM}};
  rob_uop_21_xcpt_ae_if = _RAND_1877[0:0];
  _RAND_1878 = {1{`RANDOM}};
  rob_uop_21_xcpt_ma_if = _RAND_1878[0:0];
  _RAND_1879 = {1{`RANDOM}};
  rob_uop_21_bp_debug_if = _RAND_1879[0:0];
  _RAND_1880 = {1{`RANDOM}};
  rob_uop_21_bp_xcpt_if = _RAND_1880[0:0];
  _RAND_1881 = {1{`RANDOM}};
  rob_uop_21_debug_fsrc = _RAND_1881[1:0];
  _RAND_1882 = {1{`RANDOM}};
  rob_uop_21_debug_tsrc = _RAND_1882[1:0];
  _RAND_1883 = {1{`RANDOM}};
  rob_uop_22_uopc = _RAND_1883[6:0];
  _RAND_1884 = {1{`RANDOM}};
  rob_uop_22_inst = _RAND_1884[31:0];
  _RAND_1885 = {1{`RANDOM}};
  rob_uop_22_debug_inst = _RAND_1885[31:0];
  _RAND_1886 = {1{`RANDOM}};
  rob_uop_22_is_rvc = _RAND_1886[0:0];
  _RAND_1887 = {2{`RANDOM}};
  rob_uop_22_debug_pc = _RAND_1887[39:0];
  _RAND_1888 = {1{`RANDOM}};
  rob_uop_22_iq_type = _RAND_1888[2:0];
  _RAND_1889 = {1{`RANDOM}};
  rob_uop_22_fu_code = _RAND_1889[9:0];
  _RAND_1890 = {1{`RANDOM}};
  rob_uop_22_ctrl_br_type = _RAND_1890[3:0];
  _RAND_1891 = {1{`RANDOM}};
  rob_uop_22_ctrl_op1_sel = _RAND_1891[1:0];
  _RAND_1892 = {1{`RANDOM}};
  rob_uop_22_ctrl_op2_sel = _RAND_1892[2:0];
  _RAND_1893 = {1{`RANDOM}};
  rob_uop_22_ctrl_imm_sel = _RAND_1893[2:0];
  _RAND_1894 = {1{`RANDOM}};
  rob_uop_22_ctrl_op_fcn = _RAND_1894[3:0];
  _RAND_1895 = {1{`RANDOM}};
  rob_uop_22_ctrl_fcn_dw = _RAND_1895[0:0];
  _RAND_1896 = {1{`RANDOM}};
  rob_uop_22_ctrl_csr_cmd = _RAND_1896[2:0];
  _RAND_1897 = {1{`RANDOM}};
  rob_uop_22_ctrl_is_load = _RAND_1897[0:0];
  _RAND_1898 = {1{`RANDOM}};
  rob_uop_22_ctrl_is_sta = _RAND_1898[0:0];
  _RAND_1899 = {1{`RANDOM}};
  rob_uop_22_ctrl_is_std = _RAND_1899[0:0];
  _RAND_1900 = {1{`RANDOM}};
  rob_uop_22_iw_state = _RAND_1900[1:0];
  _RAND_1901 = {1{`RANDOM}};
  rob_uop_22_iw_p1_poisoned = _RAND_1901[0:0];
  _RAND_1902 = {1{`RANDOM}};
  rob_uop_22_iw_p2_poisoned = _RAND_1902[0:0];
  _RAND_1903 = {1{`RANDOM}};
  rob_uop_22_is_br = _RAND_1903[0:0];
  _RAND_1904 = {1{`RANDOM}};
  rob_uop_22_is_jalr = _RAND_1904[0:0];
  _RAND_1905 = {1{`RANDOM}};
  rob_uop_22_is_jal = _RAND_1905[0:0];
  _RAND_1906 = {1{`RANDOM}};
  rob_uop_22_is_sfb = _RAND_1906[0:0];
  _RAND_1907 = {1{`RANDOM}};
  rob_uop_22_br_mask = _RAND_1907[7:0];
  _RAND_1908 = {1{`RANDOM}};
  rob_uop_22_br_tag = _RAND_1908[2:0];
  _RAND_1909 = {1{`RANDOM}};
  rob_uop_22_ftq_idx = _RAND_1909[3:0];
  _RAND_1910 = {1{`RANDOM}};
  rob_uop_22_edge_inst = _RAND_1910[0:0];
  _RAND_1911 = {1{`RANDOM}};
  rob_uop_22_pc_lob = _RAND_1911[5:0];
  _RAND_1912 = {1{`RANDOM}};
  rob_uop_22_taken = _RAND_1912[0:0];
  _RAND_1913 = {1{`RANDOM}};
  rob_uop_22_imm_packed = _RAND_1913[19:0];
  _RAND_1914 = {1{`RANDOM}};
  rob_uop_22_csr_addr = _RAND_1914[11:0];
  _RAND_1915 = {1{`RANDOM}};
  rob_uop_22_rob_idx = _RAND_1915[4:0];
  _RAND_1916 = {1{`RANDOM}};
  rob_uop_22_ldq_idx = _RAND_1916[2:0];
  _RAND_1917 = {1{`RANDOM}};
  rob_uop_22_stq_idx = _RAND_1917[2:0];
  _RAND_1918 = {1{`RANDOM}};
  rob_uop_22_rxq_idx = _RAND_1918[1:0];
  _RAND_1919 = {1{`RANDOM}};
  rob_uop_22_pdst = _RAND_1919[5:0];
  _RAND_1920 = {1{`RANDOM}};
  rob_uop_22_prs1 = _RAND_1920[5:0];
  _RAND_1921 = {1{`RANDOM}};
  rob_uop_22_prs2 = _RAND_1921[5:0];
  _RAND_1922 = {1{`RANDOM}};
  rob_uop_22_prs3 = _RAND_1922[5:0];
  _RAND_1923 = {1{`RANDOM}};
  rob_uop_22_ppred = _RAND_1923[3:0];
  _RAND_1924 = {1{`RANDOM}};
  rob_uop_22_prs1_busy = _RAND_1924[0:0];
  _RAND_1925 = {1{`RANDOM}};
  rob_uop_22_prs2_busy = _RAND_1925[0:0];
  _RAND_1926 = {1{`RANDOM}};
  rob_uop_22_prs3_busy = _RAND_1926[0:0];
  _RAND_1927 = {1{`RANDOM}};
  rob_uop_22_ppred_busy = _RAND_1927[0:0];
  _RAND_1928 = {1{`RANDOM}};
  rob_uop_22_stale_pdst = _RAND_1928[5:0];
  _RAND_1929 = {1{`RANDOM}};
  rob_uop_22_exception = _RAND_1929[0:0];
  _RAND_1930 = {2{`RANDOM}};
  rob_uop_22_exc_cause = _RAND_1930[63:0];
  _RAND_1931 = {1{`RANDOM}};
  rob_uop_22_bypassable = _RAND_1931[0:0];
  _RAND_1932 = {1{`RANDOM}};
  rob_uop_22_mem_cmd = _RAND_1932[4:0];
  _RAND_1933 = {1{`RANDOM}};
  rob_uop_22_mem_size = _RAND_1933[1:0];
  _RAND_1934 = {1{`RANDOM}};
  rob_uop_22_mem_signed = _RAND_1934[0:0];
  _RAND_1935 = {1{`RANDOM}};
  rob_uop_22_is_fence = _RAND_1935[0:0];
  _RAND_1936 = {1{`RANDOM}};
  rob_uop_22_is_fencei = _RAND_1936[0:0];
  _RAND_1937 = {1{`RANDOM}};
  rob_uop_22_is_amo = _RAND_1937[0:0];
  _RAND_1938 = {1{`RANDOM}};
  rob_uop_22_uses_ldq = _RAND_1938[0:0];
  _RAND_1939 = {1{`RANDOM}};
  rob_uop_22_uses_stq = _RAND_1939[0:0];
  _RAND_1940 = {1{`RANDOM}};
  rob_uop_22_is_sys_pc2epc = _RAND_1940[0:0];
  _RAND_1941 = {1{`RANDOM}};
  rob_uop_22_is_unique = _RAND_1941[0:0];
  _RAND_1942 = {1{`RANDOM}};
  rob_uop_22_flush_on_commit = _RAND_1942[0:0];
  _RAND_1943 = {1{`RANDOM}};
  rob_uop_22_ldst_is_rs1 = _RAND_1943[0:0];
  _RAND_1944 = {1{`RANDOM}};
  rob_uop_22_ldst = _RAND_1944[5:0];
  _RAND_1945 = {1{`RANDOM}};
  rob_uop_22_lrs1 = _RAND_1945[5:0];
  _RAND_1946 = {1{`RANDOM}};
  rob_uop_22_lrs2 = _RAND_1946[5:0];
  _RAND_1947 = {1{`RANDOM}};
  rob_uop_22_lrs3 = _RAND_1947[5:0];
  _RAND_1948 = {1{`RANDOM}};
  rob_uop_22_ldst_val = _RAND_1948[0:0];
  _RAND_1949 = {1{`RANDOM}};
  rob_uop_22_dst_rtype = _RAND_1949[1:0];
  _RAND_1950 = {1{`RANDOM}};
  rob_uop_22_lrs1_rtype = _RAND_1950[1:0];
  _RAND_1951 = {1{`RANDOM}};
  rob_uop_22_lrs2_rtype = _RAND_1951[1:0];
  _RAND_1952 = {1{`RANDOM}};
  rob_uop_22_frs3_en = _RAND_1952[0:0];
  _RAND_1953 = {1{`RANDOM}};
  rob_uop_22_fp_val = _RAND_1953[0:0];
  _RAND_1954 = {1{`RANDOM}};
  rob_uop_22_fp_single = _RAND_1954[0:0];
  _RAND_1955 = {1{`RANDOM}};
  rob_uop_22_xcpt_pf_if = _RAND_1955[0:0];
  _RAND_1956 = {1{`RANDOM}};
  rob_uop_22_xcpt_ae_if = _RAND_1956[0:0];
  _RAND_1957 = {1{`RANDOM}};
  rob_uop_22_xcpt_ma_if = _RAND_1957[0:0];
  _RAND_1958 = {1{`RANDOM}};
  rob_uop_22_bp_debug_if = _RAND_1958[0:0];
  _RAND_1959 = {1{`RANDOM}};
  rob_uop_22_bp_xcpt_if = _RAND_1959[0:0];
  _RAND_1960 = {1{`RANDOM}};
  rob_uop_22_debug_fsrc = _RAND_1960[1:0];
  _RAND_1961 = {1{`RANDOM}};
  rob_uop_22_debug_tsrc = _RAND_1961[1:0];
  _RAND_1962 = {1{`RANDOM}};
  rob_uop_23_uopc = _RAND_1962[6:0];
  _RAND_1963 = {1{`RANDOM}};
  rob_uop_23_inst = _RAND_1963[31:0];
  _RAND_1964 = {1{`RANDOM}};
  rob_uop_23_debug_inst = _RAND_1964[31:0];
  _RAND_1965 = {1{`RANDOM}};
  rob_uop_23_is_rvc = _RAND_1965[0:0];
  _RAND_1966 = {2{`RANDOM}};
  rob_uop_23_debug_pc = _RAND_1966[39:0];
  _RAND_1967 = {1{`RANDOM}};
  rob_uop_23_iq_type = _RAND_1967[2:0];
  _RAND_1968 = {1{`RANDOM}};
  rob_uop_23_fu_code = _RAND_1968[9:0];
  _RAND_1969 = {1{`RANDOM}};
  rob_uop_23_ctrl_br_type = _RAND_1969[3:0];
  _RAND_1970 = {1{`RANDOM}};
  rob_uop_23_ctrl_op1_sel = _RAND_1970[1:0];
  _RAND_1971 = {1{`RANDOM}};
  rob_uop_23_ctrl_op2_sel = _RAND_1971[2:0];
  _RAND_1972 = {1{`RANDOM}};
  rob_uop_23_ctrl_imm_sel = _RAND_1972[2:0];
  _RAND_1973 = {1{`RANDOM}};
  rob_uop_23_ctrl_op_fcn = _RAND_1973[3:0];
  _RAND_1974 = {1{`RANDOM}};
  rob_uop_23_ctrl_fcn_dw = _RAND_1974[0:0];
  _RAND_1975 = {1{`RANDOM}};
  rob_uop_23_ctrl_csr_cmd = _RAND_1975[2:0];
  _RAND_1976 = {1{`RANDOM}};
  rob_uop_23_ctrl_is_load = _RAND_1976[0:0];
  _RAND_1977 = {1{`RANDOM}};
  rob_uop_23_ctrl_is_sta = _RAND_1977[0:0];
  _RAND_1978 = {1{`RANDOM}};
  rob_uop_23_ctrl_is_std = _RAND_1978[0:0];
  _RAND_1979 = {1{`RANDOM}};
  rob_uop_23_iw_state = _RAND_1979[1:0];
  _RAND_1980 = {1{`RANDOM}};
  rob_uop_23_iw_p1_poisoned = _RAND_1980[0:0];
  _RAND_1981 = {1{`RANDOM}};
  rob_uop_23_iw_p2_poisoned = _RAND_1981[0:0];
  _RAND_1982 = {1{`RANDOM}};
  rob_uop_23_is_br = _RAND_1982[0:0];
  _RAND_1983 = {1{`RANDOM}};
  rob_uop_23_is_jalr = _RAND_1983[0:0];
  _RAND_1984 = {1{`RANDOM}};
  rob_uop_23_is_jal = _RAND_1984[0:0];
  _RAND_1985 = {1{`RANDOM}};
  rob_uop_23_is_sfb = _RAND_1985[0:0];
  _RAND_1986 = {1{`RANDOM}};
  rob_uop_23_br_mask = _RAND_1986[7:0];
  _RAND_1987 = {1{`RANDOM}};
  rob_uop_23_br_tag = _RAND_1987[2:0];
  _RAND_1988 = {1{`RANDOM}};
  rob_uop_23_ftq_idx = _RAND_1988[3:0];
  _RAND_1989 = {1{`RANDOM}};
  rob_uop_23_edge_inst = _RAND_1989[0:0];
  _RAND_1990 = {1{`RANDOM}};
  rob_uop_23_pc_lob = _RAND_1990[5:0];
  _RAND_1991 = {1{`RANDOM}};
  rob_uop_23_taken = _RAND_1991[0:0];
  _RAND_1992 = {1{`RANDOM}};
  rob_uop_23_imm_packed = _RAND_1992[19:0];
  _RAND_1993 = {1{`RANDOM}};
  rob_uop_23_csr_addr = _RAND_1993[11:0];
  _RAND_1994 = {1{`RANDOM}};
  rob_uop_23_rob_idx = _RAND_1994[4:0];
  _RAND_1995 = {1{`RANDOM}};
  rob_uop_23_ldq_idx = _RAND_1995[2:0];
  _RAND_1996 = {1{`RANDOM}};
  rob_uop_23_stq_idx = _RAND_1996[2:0];
  _RAND_1997 = {1{`RANDOM}};
  rob_uop_23_rxq_idx = _RAND_1997[1:0];
  _RAND_1998 = {1{`RANDOM}};
  rob_uop_23_pdst = _RAND_1998[5:0];
  _RAND_1999 = {1{`RANDOM}};
  rob_uop_23_prs1 = _RAND_1999[5:0];
  _RAND_2000 = {1{`RANDOM}};
  rob_uop_23_prs2 = _RAND_2000[5:0];
  _RAND_2001 = {1{`RANDOM}};
  rob_uop_23_prs3 = _RAND_2001[5:0];
  _RAND_2002 = {1{`RANDOM}};
  rob_uop_23_ppred = _RAND_2002[3:0];
  _RAND_2003 = {1{`RANDOM}};
  rob_uop_23_prs1_busy = _RAND_2003[0:0];
  _RAND_2004 = {1{`RANDOM}};
  rob_uop_23_prs2_busy = _RAND_2004[0:0];
  _RAND_2005 = {1{`RANDOM}};
  rob_uop_23_prs3_busy = _RAND_2005[0:0];
  _RAND_2006 = {1{`RANDOM}};
  rob_uop_23_ppred_busy = _RAND_2006[0:0];
  _RAND_2007 = {1{`RANDOM}};
  rob_uop_23_stale_pdst = _RAND_2007[5:0];
  _RAND_2008 = {1{`RANDOM}};
  rob_uop_23_exception = _RAND_2008[0:0];
  _RAND_2009 = {2{`RANDOM}};
  rob_uop_23_exc_cause = _RAND_2009[63:0];
  _RAND_2010 = {1{`RANDOM}};
  rob_uop_23_bypassable = _RAND_2010[0:0];
  _RAND_2011 = {1{`RANDOM}};
  rob_uop_23_mem_cmd = _RAND_2011[4:0];
  _RAND_2012 = {1{`RANDOM}};
  rob_uop_23_mem_size = _RAND_2012[1:0];
  _RAND_2013 = {1{`RANDOM}};
  rob_uop_23_mem_signed = _RAND_2013[0:0];
  _RAND_2014 = {1{`RANDOM}};
  rob_uop_23_is_fence = _RAND_2014[0:0];
  _RAND_2015 = {1{`RANDOM}};
  rob_uop_23_is_fencei = _RAND_2015[0:0];
  _RAND_2016 = {1{`RANDOM}};
  rob_uop_23_is_amo = _RAND_2016[0:0];
  _RAND_2017 = {1{`RANDOM}};
  rob_uop_23_uses_ldq = _RAND_2017[0:0];
  _RAND_2018 = {1{`RANDOM}};
  rob_uop_23_uses_stq = _RAND_2018[0:0];
  _RAND_2019 = {1{`RANDOM}};
  rob_uop_23_is_sys_pc2epc = _RAND_2019[0:0];
  _RAND_2020 = {1{`RANDOM}};
  rob_uop_23_is_unique = _RAND_2020[0:0];
  _RAND_2021 = {1{`RANDOM}};
  rob_uop_23_flush_on_commit = _RAND_2021[0:0];
  _RAND_2022 = {1{`RANDOM}};
  rob_uop_23_ldst_is_rs1 = _RAND_2022[0:0];
  _RAND_2023 = {1{`RANDOM}};
  rob_uop_23_ldst = _RAND_2023[5:0];
  _RAND_2024 = {1{`RANDOM}};
  rob_uop_23_lrs1 = _RAND_2024[5:0];
  _RAND_2025 = {1{`RANDOM}};
  rob_uop_23_lrs2 = _RAND_2025[5:0];
  _RAND_2026 = {1{`RANDOM}};
  rob_uop_23_lrs3 = _RAND_2026[5:0];
  _RAND_2027 = {1{`RANDOM}};
  rob_uop_23_ldst_val = _RAND_2027[0:0];
  _RAND_2028 = {1{`RANDOM}};
  rob_uop_23_dst_rtype = _RAND_2028[1:0];
  _RAND_2029 = {1{`RANDOM}};
  rob_uop_23_lrs1_rtype = _RAND_2029[1:0];
  _RAND_2030 = {1{`RANDOM}};
  rob_uop_23_lrs2_rtype = _RAND_2030[1:0];
  _RAND_2031 = {1{`RANDOM}};
  rob_uop_23_frs3_en = _RAND_2031[0:0];
  _RAND_2032 = {1{`RANDOM}};
  rob_uop_23_fp_val = _RAND_2032[0:0];
  _RAND_2033 = {1{`RANDOM}};
  rob_uop_23_fp_single = _RAND_2033[0:0];
  _RAND_2034 = {1{`RANDOM}};
  rob_uop_23_xcpt_pf_if = _RAND_2034[0:0];
  _RAND_2035 = {1{`RANDOM}};
  rob_uop_23_xcpt_ae_if = _RAND_2035[0:0];
  _RAND_2036 = {1{`RANDOM}};
  rob_uop_23_xcpt_ma_if = _RAND_2036[0:0];
  _RAND_2037 = {1{`RANDOM}};
  rob_uop_23_bp_debug_if = _RAND_2037[0:0];
  _RAND_2038 = {1{`RANDOM}};
  rob_uop_23_bp_xcpt_if = _RAND_2038[0:0];
  _RAND_2039 = {1{`RANDOM}};
  rob_uop_23_debug_fsrc = _RAND_2039[1:0];
  _RAND_2040 = {1{`RANDOM}};
  rob_uop_23_debug_tsrc = _RAND_2040[1:0];
  _RAND_2041 = {1{`RANDOM}};
  rob_uop_24_uopc = _RAND_2041[6:0];
  _RAND_2042 = {1{`RANDOM}};
  rob_uop_24_inst = _RAND_2042[31:0];
  _RAND_2043 = {1{`RANDOM}};
  rob_uop_24_debug_inst = _RAND_2043[31:0];
  _RAND_2044 = {1{`RANDOM}};
  rob_uop_24_is_rvc = _RAND_2044[0:0];
  _RAND_2045 = {2{`RANDOM}};
  rob_uop_24_debug_pc = _RAND_2045[39:0];
  _RAND_2046 = {1{`RANDOM}};
  rob_uop_24_iq_type = _RAND_2046[2:0];
  _RAND_2047 = {1{`RANDOM}};
  rob_uop_24_fu_code = _RAND_2047[9:0];
  _RAND_2048 = {1{`RANDOM}};
  rob_uop_24_ctrl_br_type = _RAND_2048[3:0];
  _RAND_2049 = {1{`RANDOM}};
  rob_uop_24_ctrl_op1_sel = _RAND_2049[1:0];
  _RAND_2050 = {1{`RANDOM}};
  rob_uop_24_ctrl_op2_sel = _RAND_2050[2:0];
  _RAND_2051 = {1{`RANDOM}};
  rob_uop_24_ctrl_imm_sel = _RAND_2051[2:0];
  _RAND_2052 = {1{`RANDOM}};
  rob_uop_24_ctrl_op_fcn = _RAND_2052[3:0];
  _RAND_2053 = {1{`RANDOM}};
  rob_uop_24_ctrl_fcn_dw = _RAND_2053[0:0];
  _RAND_2054 = {1{`RANDOM}};
  rob_uop_24_ctrl_csr_cmd = _RAND_2054[2:0];
  _RAND_2055 = {1{`RANDOM}};
  rob_uop_24_ctrl_is_load = _RAND_2055[0:0];
  _RAND_2056 = {1{`RANDOM}};
  rob_uop_24_ctrl_is_sta = _RAND_2056[0:0];
  _RAND_2057 = {1{`RANDOM}};
  rob_uop_24_ctrl_is_std = _RAND_2057[0:0];
  _RAND_2058 = {1{`RANDOM}};
  rob_uop_24_iw_state = _RAND_2058[1:0];
  _RAND_2059 = {1{`RANDOM}};
  rob_uop_24_iw_p1_poisoned = _RAND_2059[0:0];
  _RAND_2060 = {1{`RANDOM}};
  rob_uop_24_iw_p2_poisoned = _RAND_2060[0:0];
  _RAND_2061 = {1{`RANDOM}};
  rob_uop_24_is_br = _RAND_2061[0:0];
  _RAND_2062 = {1{`RANDOM}};
  rob_uop_24_is_jalr = _RAND_2062[0:0];
  _RAND_2063 = {1{`RANDOM}};
  rob_uop_24_is_jal = _RAND_2063[0:0];
  _RAND_2064 = {1{`RANDOM}};
  rob_uop_24_is_sfb = _RAND_2064[0:0];
  _RAND_2065 = {1{`RANDOM}};
  rob_uop_24_br_mask = _RAND_2065[7:0];
  _RAND_2066 = {1{`RANDOM}};
  rob_uop_24_br_tag = _RAND_2066[2:0];
  _RAND_2067 = {1{`RANDOM}};
  rob_uop_24_ftq_idx = _RAND_2067[3:0];
  _RAND_2068 = {1{`RANDOM}};
  rob_uop_24_edge_inst = _RAND_2068[0:0];
  _RAND_2069 = {1{`RANDOM}};
  rob_uop_24_pc_lob = _RAND_2069[5:0];
  _RAND_2070 = {1{`RANDOM}};
  rob_uop_24_taken = _RAND_2070[0:0];
  _RAND_2071 = {1{`RANDOM}};
  rob_uop_24_imm_packed = _RAND_2071[19:0];
  _RAND_2072 = {1{`RANDOM}};
  rob_uop_24_csr_addr = _RAND_2072[11:0];
  _RAND_2073 = {1{`RANDOM}};
  rob_uop_24_rob_idx = _RAND_2073[4:0];
  _RAND_2074 = {1{`RANDOM}};
  rob_uop_24_ldq_idx = _RAND_2074[2:0];
  _RAND_2075 = {1{`RANDOM}};
  rob_uop_24_stq_idx = _RAND_2075[2:0];
  _RAND_2076 = {1{`RANDOM}};
  rob_uop_24_rxq_idx = _RAND_2076[1:0];
  _RAND_2077 = {1{`RANDOM}};
  rob_uop_24_pdst = _RAND_2077[5:0];
  _RAND_2078 = {1{`RANDOM}};
  rob_uop_24_prs1 = _RAND_2078[5:0];
  _RAND_2079 = {1{`RANDOM}};
  rob_uop_24_prs2 = _RAND_2079[5:0];
  _RAND_2080 = {1{`RANDOM}};
  rob_uop_24_prs3 = _RAND_2080[5:0];
  _RAND_2081 = {1{`RANDOM}};
  rob_uop_24_ppred = _RAND_2081[3:0];
  _RAND_2082 = {1{`RANDOM}};
  rob_uop_24_prs1_busy = _RAND_2082[0:0];
  _RAND_2083 = {1{`RANDOM}};
  rob_uop_24_prs2_busy = _RAND_2083[0:0];
  _RAND_2084 = {1{`RANDOM}};
  rob_uop_24_prs3_busy = _RAND_2084[0:0];
  _RAND_2085 = {1{`RANDOM}};
  rob_uop_24_ppred_busy = _RAND_2085[0:0];
  _RAND_2086 = {1{`RANDOM}};
  rob_uop_24_stale_pdst = _RAND_2086[5:0];
  _RAND_2087 = {1{`RANDOM}};
  rob_uop_24_exception = _RAND_2087[0:0];
  _RAND_2088 = {2{`RANDOM}};
  rob_uop_24_exc_cause = _RAND_2088[63:0];
  _RAND_2089 = {1{`RANDOM}};
  rob_uop_24_bypassable = _RAND_2089[0:0];
  _RAND_2090 = {1{`RANDOM}};
  rob_uop_24_mem_cmd = _RAND_2090[4:0];
  _RAND_2091 = {1{`RANDOM}};
  rob_uop_24_mem_size = _RAND_2091[1:0];
  _RAND_2092 = {1{`RANDOM}};
  rob_uop_24_mem_signed = _RAND_2092[0:0];
  _RAND_2093 = {1{`RANDOM}};
  rob_uop_24_is_fence = _RAND_2093[0:0];
  _RAND_2094 = {1{`RANDOM}};
  rob_uop_24_is_fencei = _RAND_2094[0:0];
  _RAND_2095 = {1{`RANDOM}};
  rob_uop_24_is_amo = _RAND_2095[0:0];
  _RAND_2096 = {1{`RANDOM}};
  rob_uop_24_uses_ldq = _RAND_2096[0:0];
  _RAND_2097 = {1{`RANDOM}};
  rob_uop_24_uses_stq = _RAND_2097[0:0];
  _RAND_2098 = {1{`RANDOM}};
  rob_uop_24_is_sys_pc2epc = _RAND_2098[0:0];
  _RAND_2099 = {1{`RANDOM}};
  rob_uop_24_is_unique = _RAND_2099[0:0];
  _RAND_2100 = {1{`RANDOM}};
  rob_uop_24_flush_on_commit = _RAND_2100[0:0];
  _RAND_2101 = {1{`RANDOM}};
  rob_uop_24_ldst_is_rs1 = _RAND_2101[0:0];
  _RAND_2102 = {1{`RANDOM}};
  rob_uop_24_ldst = _RAND_2102[5:0];
  _RAND_2103 = {1{`RANDOM}};
  rob_uop_24_lrs1 = _RAND_2103[5:0];
  _RAND_2104 = {1{`RANDOM}};
  rob_uop_24_lrs2 = _RAND_2104[5:0];
  _RAND_2105 = {1{`RANDOM}};
  rob_uop_24_lrs3 = _RAND_2105[5:0];
  _RAND_2106 = {1{`RANDOM}};
  rob_uop_24_ldst_val = _RAND_2106[0:0];
  _RAND_2107 = {1{`RANDOM}};
  rob_uop_24_dst_rtype = _RAND_2107[1:0];
  _RAND_2108 = {1{`RANDOM}};
  rob_uop_24_lrs1_rtype = _RAND_2108[1:0];
  _RAND_2109 = {1{`RANDOM}};
  rob_uop_24_lrs2_rtype = _RAND_2109[1:0];
  _RAND_2110 = {1{`RANDOM}};
  rob_uop_24_frs3_en = _RAND_2110[0:0];
  _RAND_2111 = {1{`RANDOM}};
  rob_uop_24_fp_val = _RAND_2111[0:0];
  _RAND_2112 = {1{`RANDOM}};
  rob_uop_24_fp_single = _RAND_2112[0:0];
  _RAND_2113 = {1{`RANDOM}};
  rob_uop_24_xcpt_pf_if = _RAND_2113[0:0];
  _RAND_2114 = {1{`RANDOM}};
  rob_uop_24_xcpt_ae_if = _RAND_2114[0:0];
  _RAND_2115 = {1{`RANDOM}};
  rob_uop_24_xcpt_ma_if = _RAND_2115[0:0];
  _RAND_2116 = {1{`RANDOM}};
  rob_uop_24_bp_debug_if = _RAND_2116[0:0];
  _RAND_2117 = {1{`RANDOM}};
  rob_uop_24_bp_xcpt_if = _RAND_2117[0:0];
  _RAND_2118 = {1{`RANDOM}};
  rob_uop_24_debug_fsrc = _RAND_2118[1:0];
  _RAND_2119 = {1{`RANDOM}};
  rob_uop_24_debug_tsrc = _RAND_2119[1:0];
  _RAND_2120 = {1{`RANDOM}};
  rob_uop_25_uopc = _RAND_2120[6:0];
  _RAND_2121 = {1{`RANDOM}};
  rob_uop_25_inst = _RAND_2121[31:0];
  _RAND_2122 = {1{`RANDOM}};
  rob_uop_25_debug_inst = _RAND_2122[31:0];
  _RAND_2123 = {1{`RANDOM}};
  rob_uop_25_is_rvc = _RAND_2123[0:0];
  _RAND_2124 = {2{`RANDOM}};
  rob_uop_25_debug_pc = _RAND_2124[39:0];
  _RAND_2125 = {1{`RANDOM}};
  rob_uop_25_iq_type = _RAND_2125[2:0];
  _RAND_2126 = {1{`RANDOM}};
  rob_uop_25_fu_code = _RAND_2126[9:0];
  _RAND_2127 = {1{`RANDOM}};
  rob_uop_25_ctrl_br_type = _RAND_2127[3:0];
  _RAND_2128 = {1{`RANDOM}};
  rob_uop_25_ctrl_op1_sel = _RAND_2128[1:0];
  _RAND_2129 = {1{`RANDOM}};
  rob_uop_25_ctrl_op2_sel = _RAND_2129[2:0];
  _RAND_2130 = {1{`RANDOM}};
  rob_uop_25_ctrl_imm_sel = _RAND_2130[2:0];
  _RAND_2131 = {1{`RANDOM}};
  rob_uop_25_ctrl_op_fcn = _RAND_2131[3:0];
  _RAND_2132 = {1{`RANDOM}};
  rob_uop_25_ctrl_fcn_dw = _RAND_2132[0:0];
  _RAND_2133 = {1{`RANDOM}};
  rob_uop_25_ctrl_csr_cmd = _RAND_2133[2:0];
  _RAND_2134 = {1{`RANDOM}};
  rob_uop_25_ctrl_is_load = _RAND_2134[0:0];
  _RAND_2135 = {1{`RANDOM}};
  rob_uop_25_ctrl_is_sta = _RAND_2135[0:0];
  _RAND_2136 = {1{`RANDOM}};
  rob_uop_25_ctrl_is_std = _RAND_2136[0:0];
  _RAND_2137 = {1{`RANDOM}};
  rob_uop_25_iw_state = _RAND_2137[1:0];
  _RAND_2138 = {1{`RANDOM}};
  rob_uop_25_iw_p1_poisoned = _RAND_2138[0:0];
  _RAND_2139 = {1{`RANDOM}};
  rob_uop_25_iw_p2_poisoned = _RAND_2139[0:0];
  _RAND_2140 = {1{`RANDOM}};
  rob_uop_25_is_br = _RAND_2140[0:0];
  _RAND_2141 = {1{`RANDOM}};
  rob_uop_25_is_jalr = _RAND_2141[0:0];
  _RAND_2142 = {1{`RANDOM}};
  rob_uop_25_is_jal = _RAND_2142[0:0];
  _RAND_2143 = {1{`RANDOM}};
  rob_uop_25_is_sfb = _RAND_2143[0:0];
  _RAND_2144 = {1{`RANDOM}};
  rob_uop_25_br_mask = _RAND_2144[7:0];
  _RAND_2145 = {1{`RANDOM}};
  rob_uop_25_br_tag = _RAND_2145[2:0];
  _RAND_2146 = {1{`RANDOM}};
  rob_uop_25_ftq_idx = _RAND_2146[3:0];
  _RAND_2147 = {1{`RANDOM}};
  rob_uop_25_edge_inst = _RAND_2147[0:0];
  _RAND_2148 = {1{`RANDOM}};
  rob_uop_25_pc_lob = _RAND_2148[5:0];
  _RAND_2149 = {1{`RANDOM}};
  rob_uop_25_taken = _RAND_2149[0:0];
  _RAND_2150 = {1{`RANDOM}};
  rob_uop_25_imm_packed = _RAND_2150[19:0];
  _RAND_2151 = {1{`RANDOM}};
  rob_uop_25_csr_addr = _RAND_2151[11:0];
  _RAND_2152 = {1{`RANDOM}};
  rob_uop_25_rob_idx = _RAND_2152[4:0];
  _RAND_2153 = {1{`RANDOM}};
  rob_uop_25_ldq_idx = _RAND_2153[2:0];
  _RAND_2154 = {1{`RANDOM}};
  rob_uop_25_stq_idx = _RAND_2154[2:0];
  _RAND_2155 = {1{`RANDOM}};
  rob_uop_25_rxq_idx = _RAND_2155[1:0];
  _RAND_2156 = {1{`RANDOM}};
  rob_uop_25_pdst = _RAND_2156[5:0];
  _RAND_2157 = {1{`RANDOM}};
  rob_uop_25_prs1 = _RAND_2157[5:0];
  _RAND_2158 = {1{`RANDOM}};
  rob_uop_25_prs2 = _RAND_2158[5:0];
  _RAND_2159 = {1{`RANDOM}};
  rob_uop_25_prs3 = _RAND_2159[5:0];
  _RAND_2160 = {1{`RANDOM}};
  rob_uop_25_ppred = _RAND_2160[3:0];
  _RAND_2161 = {1{`RANDOM}};
  rob_uop_25_prs1_busy = _RAND_2161[0:0];
  _RAND_2162 = {1{`RANDOM}};
  rob_uop_25_prs2_busy = _RAND_2162[0:0];
  _RAND_2163 = {1{`RANDOM}};
  rob_uop_25_prs3_busy = _RAND_2163[0:0];
  _RAND_2164 = {1{`RANDOM}};
  rob_uop_25_ppred_busy = _RAND_2164[0:0];
  _RAND_2165 = {1{`RANDOM}};
  rob_uop_25_stale_pdst = _RAND_2165[5:0];
  _RAND_2166 = {1{`RANDOM}};
  rob_uop_25_exception = _RAND_2166[0:0];
  _RAND_2167 = {2{`RANDOM}};
  rob_uop_25_exc_cause = _RAND_2167[63:0];
  _RAND_2168 = {1{`RANDOM}};
  rob_uop_25_bypassable = _RAND_2168[0:0];
  _RAND_2169 = {1{`RANDOM}};
  rob_uop_25_mem_cmd = _RAND_2169[4:0];
  _RAND_2170 = {1{`RANDOM}};
  rob_uop_25_mem_size = _RAND_2170[1:0];
  _RAND_2171 = {1{`RANDOM}};
  rob_uop_25_mem_signed = _RAND_2171[0:0];
  _RAND_2172 = {1{`RANDOM}};
  rob_uop_25_is_fence = _RAND_2172[0:0];
  _RAND_2173 = {1{`RANDOM}};
  rob_uop_25_is_fencei = _RAND_2173[0:0];
  _RAND_2174 = {1{`RANDOM}};
  rob_uop_25_is_amo = _RAND_2174[0:0];
  _RAND_2175 = {1{`RANDOM}};
  rob_uop_25_uses_ldq = _RAND_2175[0:0];
  _RAND_2176 = {1{`RANDOM}};
  rob_uop_25_uses_stq = _RAND_2176[0:0];
  _RAND_2177 = {1{`RANDOM}};
  rob_uop_25_is_sys_pc2epc = _RAND_2177[0:0];
  _RAND_2178 = {1{`RANDOM}};
  rob_uop_25_is_unique = _RAND_2178[0:0];
  _RAND_2179 = {1{`RANDOM}};
  rob_uop_25_flush_on_commit = _RAND_2179[0:0];
  _RAND_2180 = {1{`RANDOM}};
  rob_uop_25_ldst_is_rs1 = _RAND_2180[0:0];
  _RAND_2181 = {1{`RANDOM}};
  rob_uop_25_ldst = _RAND_2181[5:0];
  _RAND_2182 = {1{`RANDOM}};
  rob_uop_25_lrs1 = _RAND_2182[5:0];
  _RAND_2183 = {1{`RANDOM}};
  rob_uop_25_lrs2 = _RAND_2183[5:0];
  _RAND_2184 = {1{`RANDOM}};
  rob_uop_25_lrs3 = _RAND_2184[5:0];
  _RAND_2185 = {1{`RANDOM}};
  rob_uop_25_ldst_val = _RAND_2185[0:0];
  _RAND_2186 = {1{`RANDOM}};
  rob_uop_25_dst_rtype = _RAND_2186[1:0];
  _RAND_2187 = {1{`RANDOM}};
  rob_uop_25_lrs1_rtype = _RAND_2187[1:0];
  _RAND_2188 = {1{`RANDOM}};
  rob_uop_25_lrs2_rtype = _RAND_2188[1:0];
  _RAND_2189 = {1{`RANDOM}};
  rob_uop_25_frs3_en = _RAND_2189[0:0];
  _RAND_2190 = {1{`RANDOM}};
  rob_uop_25_fp_val = _RAND_2190[0:0];
  _RAND_2191 = {1{`RANDOM}};
  rob_uop_25_fp_single = _RAND_2191[0:0];
  _RAND_2192 = {1{`RANDOM}};
  rob_uop_25_xcpt_pf_if = _RAND_2192[0:0];
  _RAND_2193 = {1{`RANDOM}};
  rob_uop_25_xcpt_ae_if = _RAND_2193[0:0];
  _RAND_2194 = {1{`RANDOM}};
  rob_uop_25_xcpt_ma_if = _RAND_2194[0:0];
  _RAND_2195 = {1{`RANDOM}};
  rob_uop_25_bp_debug_if = _RAND_2195[0:0];
  _RAND_2196 = {1{`RANDOM}};
  rob_uop_25_bp_xcpt_if = _RAND_2196[0:0];
  _RAND_2197 = {1{`RANDOM}};
  rob_uop_25_debug_fsrc = _RAND_2197[1:0];
  _RAND_2198 = {1{`RANDOM}};
  rob_uop_25_debug_tsrc = _RAND_2198[1:0];
  _RAND_2199 = {1{`RANDOM}};
  rob_uop_26_uopc = _RAND_2199[6:0];
  _RAND_2200 = {1{`RANDOM}};
  rob_uop_26_inst = _RAND_2200[31:0];
  _RAND_2201 = {1{`RANDOM}};
  rob_uop_26_debug_inst = _RAND_2201[31:0];
  _RAND_2202 = {1{`RANDOM}};
  rob_uop_26_is_rvc = _RAND_2202[0:0];
  _RAND_2203 = {2{`RANDOM}};
  rob_uop_26_debug_pc = _RAND_2203[39:0];
  _RAND_2204 = {1{`RANDOM}};
  rob_uop_26_iq_type = _RAND_2204[2:0];
  _RAND_2205 = {1{`RANDOM}};
  rob_uop_26_fu_code = _RAND_2205[9:0];
  _RAND_2206 = {1{`RANDOM}};
  rob_uop_26_ctrl_br_type = _RAND_2206[3:0];
  _RAND_2207 = {1{`RANDOM}};
  rob_uop_26_ctrl_op1_sel = _RAND_2207[1:0];
  _RAND_2208 = {1{`RANDOM}};
  rob_uop_26_ctrl_op2_sel = _RAND_2208[2:0];
  _RAND_2209 = {1{`RANDOM}};
  rob_uop_26_ctrl_imm_sel = _RAND_2209[2:0];
  _RAND_2210 = {1{`RANDOM}};
  rob_uop_26_ctrl_op_fcn = _RAND_2210[3:0];
  _RAND_2211 = {1{`RANDOM}};
  rob_uop_26_ctrl_fcn_dw = _RAND_2211[0:0];
  _RAND_2212 = {1{`RANDOM}};
  rob_uop_26_ctrl_csr_cmd = _RAND_2212[2:0];
  _RAND_2213 = {1{`RANDOM}};
  rob_uop_26_ctrl_is_load = _RAND_2213[0:0];
  _RAND_2214 = {1{`RANDOM}};
  rob_uop_26_ctrl_is_sta = _RAND_2214[0:0];
  _RAND_2215 = {1{`RANDOM}};
  rob_uop_26_ctrl_is_std = _RAND_2215[0:0];
  _RAND_2216 = {1{`RANDOM}};
  rob_uop_26_iw_state = _RAND_2216[1:0];
  _RAND_2217 = {1{`RANDOM}};
  rob_uop_26_iw_p1_poisoned = _RAND_2217[0:0];
  _RAND_2218 = {1{`RANDOM}};
  rob_uop_26_iw_p2_poisoned = _RAND_2218[0:0];
  _RAND_2219 = {1{`RANDOM}};
  rob_uop_26_is_br = _RAND_2219[0:0];
  _RAND_2220 = {1{`RANDOM}};
  rob_uop_26_is_jalr = _RAND_2220[0:0];
  _RAND_2221 = {1{`RANDOM}};
  rob_uop_26_is_jal = _RAND_2221[0:0];
  _RAND_2222 = {1{`RANDOM}};
  rob_uop_26_is_sfb = _RAND_2222[0:0];
  _RAND_2223 = {1{`RANDOM}};
  rob_uop_26_br_mask = _RAND_2223[7:0];
  _RAND_2224 = {1{`RANDOM}};
  rob_uop_26_br_tag = _RAND_2224[2:0];
  _RAND_2225 = {1{`RANDOM}};
  rob_uop_26_ftq_idx = _RAND_2225[3:0];
  _RAND_2226 = {1{`RANDOM}};
  rob_uop_26_edge_inst = _RAND_2226[0:0];
  _RAND_2227 = {1{`RANDOM}};
  rob_uop_26_pc_lob = _RAND_2227[5:0];
  _RAND_2228 = {1{`RANDOM}};
  rob_uop_26_taken = _RAND_2228[0:0];
  _RAND_2229 = {1{`RANDOM}};
  rob_uop_26_imm_packed = _RAND_2229[19:0];
  _RAND_2230 = {1{`RANDOM}};
  rob_uop_26_csr_addr = _RAND_2230[11:0];
  _RAND_2231 = {1{`RANDOM}};
  rob_uop_26_rob_idx = _RAND_2231[4:0];
  _RAND_2232 = {1{`RANDOM}};
  rob_uop_26_ldq_idx = _RAND_2232[2:0];
  _RAND_2233 = {1{`RANDOM}};
  rob_uop_26_stq_idx = _RAND_2233[2:0];
  _RAND_2234 = {1{`RANDOM}};
  rob_uop_26_rxq_idx = _RAND_2234[1:0];
  _RAND_2235 = {1{`RANDOM}};
  rob_uop_26_pdst = _RAND_2235[5:0];
  _RAND_2236 = {1{`RANDOM}};
  rob_uop_26_prs1 = _RAND_2236[5:0];
  _RAND_2237 = {1{`RANDOM}};
  rob_uop_26_prs2 = _RAND_2237[5:0];
  _RAND_2238 = {1{`RANDOM}};
  rob_uop_26_prs3 = _RAND_2238[5:0];
  _RAND_2239 = {1{`RANDOM}};
  rob_uop_26_ppred = _RAND_2239[3:0];
  _RAND_2240 = {1{`RANDOM}};
  rob_uop_26_prs1_busy = _RAND_2240[0:0];
  _RAND_2241 = {1{`RANDOM}};
  rob_uop_26_prs2_busy = _RAND_2241[0:0];
  _RAND_2242 = {1{`RANDOM}};
  rob_uop_26_prs3_busy = _RAND_2242[0:0];
  _RAND_2243 = {1{`RANDOM}};
  rob_uop_26_ppred_busy = _RAND_2243[0:0];
  _RAND_2244 = {1{`RANDOM}};
  rob_uop_26_stale_pdst = _RAND_2244[5:0];
  _RAND_2245 = {1{`RANDOM}};
  rob_uop_26_exception = _RAND_2245[0:0];
  _RAND_2246 = {2{`RANDOM}};
  rob_uop_26_exc_cause = _RAND_2246[63:0];
  _RAND_2247 = {1{`RANDOM}};
  rob_uop_26_bypassable = _RAND_2247[0:0];
  _RAND_2248 = {1{`RANDOM}};
  rob_uop_26_mem_cmd = _RAND_2248[4:0];
  _RAND_2249 = {1{`RANDOM}};
  rob_uop_26_mem_size = _RAND_2249[1:0];
  _RAND_2250 = {1{`RANDOM}};
  rob_uop_26_mem_signed = _RAND_2250[0:0];
  _RAND_2251 = {1{`RANDOM}};
  rob_uop_26_is_fence = _RAND_2251[0:0];
  _RAND_2252 = {1{`RANDOM}};
  rob_uop_26_is_fencei = _RAND_2252[0:0];
  _RAND_2253 = {1{`RANDOM}};
  rob_uop_26_is_amo = _RAND_2253[0:0];
  _RAND_2254 = {1{`RANDOM}};
  rob_uop_26_uses_ldq = _RAND_2254[0:0];
  _RAND_2255 = {1{`RANDOM}};
  rob_uop_26_uses_stq = _RAND_2255[0:0];
  _RAND_2256 = {1{`RANDOM}};
  rob_uop_26_is_sys_pc2epc = _RAND_2256[0:0];
  _RAND_2257 = {1{`RANDOM}};
  rob_uop_26_is_unique = _RAND_2257[0:0];
  _RAND_2258 = {1{`RANDOM}};
  rob_uop_26_flush_on_commit = _RAND_2258[0:0];
  _RAND_2259 = {1{`RANDOM}};
  rob_uop_26_ldst_is_rs1 = _RAND_2259[0:0];
  _RAND_2260 = {1{`RANDOM}};
  rob_uop_26_ldst = _RAND_2260[5:0];
  _RAND_2261 = {1{`RANDOM}};
  rob_uop_26_lrs1 = _RAND_2261[5:0];
  _RAND_2262 = {1{`RANDOM}};
  rob_uop_26_lrs2 = _RAND_2262[5:0];
  _RAND_2263 = {1{`RANDOM}};
  rob_uop_26_lrs3 = _RAND_2263[5:0];
  _RAND_2264 = {1{`RANDOM}};
  rob_uop_26_ldst_val = _RAND_2264[0:0];
  _RAND_2265 = {1{`RANDOM}};
  rob_uop_26_dst_rtype = _RAND_2265[1:0];
  _RAND_2266 = {1{`RANDOM}};
  rob_uop_26_lrs1_rtype = _RAND_2266[1:0];
  _RAND_2267 = {1{`RANDOM}};
  rob_uop_26_lrs2_rtype = _RAND_2267[1:0];
  _RAND_2268 = {1{`RANDOM}};
  rob_uop_26_frs3_en = _RAND_2268[0:0];
  _RAND_2269 = {1{`RANDOM}};
  rob_uop_26_fp_val = _RAND_2269[0:0];
  _RAND_2270 = {1{`RANDOM}};
  rob_uop_26_fp_single = _RAND_2270[0:0];
  _RAND_2271 = {1{`RANDOM}};
  rob_uop_26_xcpt_pf_if = _RAND_2271[0:0];
  _RAND_2272 = {1{`RANDOM}};
  rob_uop_26_xcpt_ae_if = _RAND_2272[0:0];
  _RAND_2273 = {1{`RANDOM}};
  rob_uop_26_xcpt_ma_if = _RAND_2273[0:0];
  _RAND_2274 = {1{`RANDOM}};
  rob_uop_26_bp_debug_if = _RAND_2274[0:0];
  _RAND_2275 = {1{`RANDOM}};
  rob_uop_26_bp_xcpt_if = _RAND_2275[0:0];
  _RAND_2276 = {1{`RANDOM}};
  rob_uop_26_debug_fsrc = _RAND_2276[1:0];
  _RAND_2277 = {1{`RANDOM}};
  rob_uop_26_debug_tsrc = _RAND_2277[1:0];
  _RAND_2278 = {1{`RANDOM}};
  rob_uop_27_uopc = _RAND_2278[6:0];
  _RAND_2279 = {1{`RANDOM}};
  rob_uop_27_inst = _RAND_2279[31:0];
  _RAND_2280 = {1{`RANDOM}};
  rob_uop_27_debug_inst = _RAND_2280[31:0];
  _RAND_2281 = {1{`RANDOM}};
  rob_uop_27_is_rvc = _RAND_2281[0:0];
  _RAND_2282 = {2{`RANDOM}};
  rob_uop_27_debug_pc = _RAND_2282[39:0];
  _RAND_2283 = {1{`RANDOM}};
  rob_uop_27_iq_type = _RAND_2283[2:0];
  _RAND_2284 = {1{`RANDOM}};
  rob_uop_27_fu_code = _RAND_2284[9:0];
  _RAND_2285 = {1{`RANDOM}};
  rob_uop_27_ctrl_br_type = _RAND_2285[3:0];
  _RAND_2286 = {1{`RANDOM}};
  rob_uop_27_ctrl_op1_sel = _RAND_2286[1:0];
  _RAND_2287 = {1{`RANDOM}};
  rob_uop_27_ctrl_op2_sel = _RAND_2287[2:0];
  _RAND_2288 = {1{`RANDOM}};
  rob_uop_27_ctrl_imm_sel = _RAND_2288[2:0];
  _RAND_2289 = {1{`RANDOM}};
  rob_uop_27_ctrl_op_fcn = _RAND_2289[3:0];
  _RAND_2290 = {1{`RANDOM}};
  rob_uop_27_ctrl_fcn_dw = _RAND_2290[0:0];
  _RAND_2291 = {1{`RANDOM}};
  rob_uop_27_ctrl_csr_cmd = _RAND_2291[2:0];
  _RAND_2292 = {1{`RANDOM}};
  rob_uop_27_ctrl_is_load = _RAND_2292[0:0];
  _RAND_2293 = {1{`RANDOM}};
  rob_uop_27_ctrl_is_sta = _RAND_2293[0:0];
  _RAND_2294 = {1{`RANDOM}};
  rob_uop_27_ctrl_is_std = _RAND_2294[0:0];
  _RAND_2295 = {1{`RANDOM}};
  rob_uop_27_iw_state = _RAND_2295[1:0];
  _RAND_2296 = {1{`RANDOM}};
  rob_uop_27_iw_p1_poisoned = _RAND_2296[0:0];
  _RAND_2297 = {1{`RANDOM}};
  rob_uop_27_iw_p2_poisoned = _RAND_2297[0:0];
  _RAND_2298 = {1{`RANDOM}};
  rob_uop_27_is_br = _RAND_2298[0:0];
  _RAND_2299 = {1{`RANDOM}};
  rob_uop_27_is_jalr = _RAND_2299[0:0];
  _RAND_2300 = {1{`RANDOM}};
  rob_uop_27_is_jal = _RAND_2300[0:0];
  _RAND_2301 = {1{`RANDOM}};
  rob_uop_27_is_sfb = _RAND_2301[0:0];
  _RAND_2302 = {1{`RANDOM}};
  rob_uop_27_br_mask = _RAND_2302[7:0];
  _RAND_2303 = {1{`RANDOM}};
  rob_uop_27_br_tag = _RAND_2303[2:0];
  _RAND_2304 = {1{`RANDOM}};
  rob_uop_27_ftq_idx = _RAND_2304[3:0];
  _RAND_2305 = {1{`RANDOM}};
  rob_uop_27_edge_inst = _RAND_2305[0:0];
  _RAND_2306 = {1{`RANDOM}};
  rob_uop_27_pc_lob = _RAND_2306[5:0];
  _RAND_2307 = {1{`RANDOM}};
  rob_uop_27_taken = _RAND_2307[0:0];
  _RAND_2308 = {1{`RANDOM}};
  rob_uop_27_imm_packed = _RAND_2308[19:0];
  _RAND_2309 = {1{`RANDOM}};
  rob_uop_27_csr_addr = _RAND_2309[11:0];
  _RAND_2310 = {1{`RANDOM}};
  rob_uop_27_rob_idx = _RAND_2310[4:0];
  _RAND_2311 = {1{`RANDOM}};
  rob_uop_27_ldq_idx = _RAND_2311[2:0];
  _RAND_2312 = {1{`RANDOM}};
  rob_uop_27_stq_idx = _RAND_2312[2:0];
  _RAND_2313 = {1{`RANDOM}};
  rob_uop_27_rxq_idx = _RAND_2313[1:0];
  _RAND_2314 = {1{`RANDOM}};
  rob_uop_27_pdst = _RAND_2314[5:0];
  _RAND_2315 = {1{`RANDOM}};
  rob_uop_27_prs1 = _RAND_2315[5:0];
  _RAND_2316 = {1{`RANDOM}};
  rob_uop_27_prs2 = _RAND_2316[5:0];
  _RAND_2317 = {1{`RANDOM}};
  rob_uop_27_prs3 = _RAND_2317[5:0];
  _RAND_2318 = {1{`RANDOM}};
  rob_uop_27_ppred = _RAND_2318[3:0];
  _RAND_2319 = {1{`RANDOM}};
  rob_uop_27_prs1_busy = _RAND_2319[0:0];
  _RAND_2320 = {1{`RANDOM}};
  rob_uop_27_prs2_busy = _RAND_2320[0:0];
  _RAND_2321 = {1{`RANDOM}};
  rob_uop_27_prs3_busy = _RAND_2321[0:0];
  _RAND_2322 = {1{`RANDOM}};
  rob_uop_27_ppred_busy = _RAND_2322[0:0];
  _RAND_2323 = {1{`RANDOM}};
  rob_uop_27_stale_pdst = _RAND_2323[5:0];
  _RAND_2324 = {1{`RANDOM}};
  rob_uop_27_exception = _RAND_2324[0:0];
  _RAND_2325 = {2{`RANDOM}};
  rob_uop_27_exc_cause = _RAND_2325[63:0];
  _RAND_2326 = {1{`RANDOM}};
  rob_uop_27_bypassable = _RAND_2326[0:0];
  _RAND_2327 = {1{`RANDOM}};
  rob_uop_27_mem_cmd = _RAND_2327[4:0];
  _RAND_2328 = {1{`RANDOM}};
  rob_uop_27_mem_size = _RAND_2328[1:0];
  _RAND_2329 = {1{`RANDOM}};
  rob_uop_27_mem_signed = _RAND_2329[0:0];
  _RAND_2330 = {1{`RANDOM}};
  rob_uop_27_is_fence = _RAND_2330[0:0];
  _RAND_2331 = {1{`RANDOM}};
  rob_uop_27_is_fencei = _RAND_2331[0:0];
  _RAND_2332 = {1{`RANDOM}};
  rob_uop_27_is_amo = _RAND_2332[0:0];
  _RAND_2333 = {1{`RANDOM}};
  rob_uop_27_uses_ldq = _RAND_2333[0:0];
  _RAND_2334 = {1{`RANDOM}};
  rob_uop_27_uses_stq = _RAND_2334[0:0];
  _RAND_2335 = {1{`RANDOM}};
  rob_uop_27_is_sys_pc2epc = _RAND_2335[0:0];
  _RAND_2336 = {1{`RANDOM}};
  rob_uop_27_is_unique = _RAND_2336[0:0];
  _RAND_2337 = {1{`RANDOM}};
  rob_uop_27_flush_on_commit = _RAND_2337[0:0];
  _RAND_2338 = {1{`RANDOM}};
  rob_uop_27_ldst_is_rs1 = _RAND_2338[0:0];
  _RAND_2339 = {1{`RANDOM}};
  rob_uop_27_ldst = _RAND_2339[5:0];
  _RAND_2340 = {1{`RANDOM}};
  rob_uop_27_lrs1 = _RAND_2340[5:0];
  _RAND_2341 = {1{`RANDOM}};
  rob_uop_27_lrs2 = _RAND_2341[5:0];
  _RAND_2342 = {1{`RANDOM}};
  rob_uop_27_lrs3 = _RAND_2342[5:0];
  _RAND_2343 = {1{`RANDOM}};
  rob_uop_27_ldst_val = _RAND_2343[0:0];
  _RAND_2344 = {1{`RANDOM}};
  rob_uop_27_dst_rtype = _RAND_2344[1:0];
  _RAND_2345 = {1{`RANDOM}};
  rob_uop_27_lrs1_rtype = _RAND_2345[1:0];
  _RAND_2346 = {1{`RANDOM}};
  rob_uop_27_lrs2_rtype = _RAND_2346[1:0];
  _RAND_2347 = {1{`RANDOM}};
  rob_uop_27_frs3_en = _RAND_2347[0:0];
  _RAND_2348 = {1{`RANDOM}};
  rob_uop_27_fp_val = _RAND_2348[0:0];
  _RAND_2349 = {1{`RANDOM}};
  rob_uop_27_fp_single = _RAND_2349[0:0];
  _RAND_2350 = {1{`RANDOM}};
  rob_uop_27_xcpt_pf_if = _RAND_2350[0:0];
  _RAND_2351 = {1{`RANDOM}};
  rob_uop_27_xcpt_ae_if = _RAND_2351[0:0];
  _RAND_2352 = {1{`RANDOM}};
  rob_uop_27_xcpt_ma_if = _RAND_2352[0:0];
  _RAND_2353 = {1{`RANDOM}};
  rob_uop_27_bp_debug_if = _RAND_2353[0:0];
  _RAND_2354 = {1{`RANDOM}};
  rob_uop_27_bp_xcpt_if = _RAND_2354[0:0];
  _RAND_2355 = {1{`RANDOM}};
  rob_uop_27_debug_fsrc = _RAND_2355[1:0];
  _RAND_2356 = {1{`RANDOM}};
  rob_uop_27_debug_tsrc = _RAND_2356[1:0];
  _RAND_2357 = {1{`RANDOM}};
  rob_uop_28_uopc = _RAND_2357[6:0];
  _RAND_2358 = {1{`RANDOM}};
  rob_uop_28_inst = _RAND_2358[31:0];
  _RAND_2359 = {1{`RANDOM}};
  rob_uop_28_debug_inst = _RAND_2359[31:0];
  _RAND_2360 = {1{`RANDOM}};
  rob_uop_28_is_rvc = _RAND_2360[0:0];
  _RAND_2361 = {2{`RANDOM}};
  rob_uop_28_debug_pc = _RAND_2361[39:0];
  _RAND_2362 = {1{`RANDOM}};
  rob_uop_28_iq_type = _RAND_2362[2:0];
  _RAND_2363 = {1{`RANDOM}};
  rob_uop_28_fu_code = _RAND_2363[9:0];
  _RAND_2364 = {1{`RANDOM}};
  rob_uop_28_ctrl_br_type = _RAND_2364[3:0];
  _RAND_2365 = {1{`RANDOM}};
  rob_uop_28_ctrl_op1_sel = _RAND_2365[1:0];
  _RAND_2366 = {1{`RANDOM}};
  rob_uop_28_ctrl_op2_sel = _RAND_2366[2:0];
  _RAND_2367 = {1{`RANDOM}};
  rob_uop_28_ctrl_imm_sel = _RAND_2367[2:0];
  _RAND_2368 = {1{`RANDOM}};
  rob_uop_28_ctrl_op_fcn = _RAND_2368[3:0];
  _RAND_2369 = {1{`RANDOM}};
  rob_uop_28_ctrl_fcn_dw = _RAND_2369[0:0];
  _RAND_2370 = {1{`RANDOM}};
  rob_uop_28_ctrl_csr_cmd = _RAND_2370[2:0];
  _RAND_2371 = {1{`RANDOM}};
  rob_uop_28_ctrl_is_load = _RAND_2371[0:0];
  _RAND_2372 = {1{`RANDOM}};
  rob_uop_28_ctrl_is_sta = _RAND_2372[0:0];
  _RAND_2373 = {1{`RANDOM}};
  rob_uop_28_ctrl_is_std = _RAND_2373[0:0];
  _RAND_2374 = {1{`RANDOM}};
  rob_uop_28_iw_state = _RAND_2374[1:0];
  _RAND_2375 = {1{`RANDOM}};
  rob_uop_28_iw_p1_poisoned = _RAND_2375[0:0];
  _RAND_2376 = {1{`RANDOM}};
  rob_uop_28_iw_p2_poisoned = _RAND_2376[0:0];
  _RAND_2377 = {1{`RANDOM}};
  rob_uop_28_is_br = _RAND_2377[0:0];
  _RAND_2378 = {1{`RANDOM}};
  rob_uop_28_is_jalr = _RAND_2378[0:0];
  _RAND_2379 = {1{`RANDOM}};
  rob_uop_28_is_jal = _RAND_2379[0:0];
  _RAND_2380 = {1{`RANDOM}};
  rob_uop_28_is_sfb = _RAND_2380[0:0];
  _RAND_2381 = {1{`RANDOM}};
  rob_uop_28_br_mask = _RAND_2381[7:0];
  _RAND_2382 = {1{`RANDOM}};
  rob_uop_28_br_tag = _RAND_2382[2:0];
  _RAND_2383 = {1{`RANDOM}};
  rob_uop_28_ftq_idx = _RAND_2383[3:0];
  _RAND_2384 = {1{`RANDOM}};
  rob_uop_28_edge_inst = _RAND_2384[0:0];
  _RAND_2385 = {1{`RANDOM}};
  rob_uop_28_pc_lob = _RAND_2385[5:0];
  _RAND_2386 = {1{`RANDOM}};
  rob_uop_28_taken = _RAND_2386[0:0];
  _RAND_2387 = {1{`RANDOM}};
  rob_uop_28_imm_packed = _RAND_2387[19:0];
  _RAND_2388 = {1{`RANDOM}};
  rob_uop_28_csr_addr = _RAND_2388[11:0];
  _RAND_2389 = {1{`RANDOM}};
  rob_uop_28_rob_idx = _RAND_2389[4:0];
  _RAND_2390 = {1{`RANDOM}};
  rob_uop_28_ldq_idx = _RAND_2390[2:0];
  _RAND_2391 = {1{`RANDOM}};
  rob_uop_28_stq_idx = _RAND_2391[2:0];
  _RAND_2392 = {1{`RANDOM}};
  rob_uop_28_rxq_idx = _RAND_2392[1:0];
  _RAND_2393 = {1{`RANDOM}};
  rob_uop_28_pdst = _RAND_2393[5:0];
  _RAND_2394 = {1{`RANDOM}};
  rob_uop_28_prs1 = _RAND_2394[5:0];
  _RAND_2395 = {1{`RANDOM}};
  rob_uop_28_prs2 = _RAND_2395[5:0];
  _RAND_2396 = {1{`RANDOM}};
  rob_uop_28_prs3 = _RAND_2396[5:0];
  _RAND_2397 = {1{`RANDOM}};
  rob_uop_28_ppred = _RAND_2397[3:0];
  _RAND_2398 = {1{`RANDOM}};
  rob_uop_28_prs1_busy = _RAND_2398[0:0];
  _RAND_2399 = {1{`RANDOM}};
  rob_uop_28_prs2_busy = _RAND_2399[0:0];
  _RAND_2400 = {1{`RANDOM}};
  rob_uop_28_prs3_busy = _RAND_2400[0:0];
  _RAND_2401 = {1{`RANDOM}};
  rob_uop_28_ppred_busy = _RAND_2401[0:0];
  _RAND_2402 = {1{`RANDOM}};
  rob_uop_28_stale_pdst = _RAND_2402[5:0];
  _RAND_2403 = {1{`RANDOM}};
  rob_uop_28_exception = _RAND_2403[0:0];
  _RAND_2404 = {2{`RANDOM}};
  rob_uop_28_exc_cause = _RAND_2404[63:0];
  _RAND_2405 = {1{`RANDOM}};
  rob_uop_28_bypassable = _RAND_2405[0:0];
  _RAND_2406 = {1{`RANDOM}};
  rob_uop_28_mem_cmd = _RAND_2406[4:0];
  _RAND_2407 = {1{`RANDOM}};
  rob_uop_28_mem_size = _RAND_2407[1:0];
  _RAND_2408 = {1{`RANDOM}};
  rob_uop_28_mem_signed = _RAND_2408[0:0];
  _RAND_2409 = {1{`RANDOM}};
  rob_uop_28_is_fence = _RAND_2409[0:0];
  _RAND_2410 = {1{`RANDOM}};
  rob_uop_28_is_fencei = _RAND_2410[0:0];
  _RAND_2411 = {1{`RANDOM}};
  rob_uop_28_is_amo = _RAND_2411[0:0];
  _RAND_2412 = {1{`RANDOM}};
  rob_uop_28_uses_ldq = _RAND_2412[0:0];
  _RAND_2413 = {1{`RANDOM}};
  rob_uop_28_uses_stq = _RAND_2413[0:0];
  _RAND_2414 = {1{`RANDOM}};
  rob_uop_28_is_sys_pc2epc = _RAND_2414[0:0];
  _RAND_2415 = {1{`RANDOM}};
  rob_uop_28_is_unique = _RAND_2415[0:0];
  _RAND_2416 = {1{`RANDOM}};
  rob_uop_28_flush_on_commit = _RAND_2416[0:0];
  _RAND_2417 = {1{`RANDOM}};
  rob_uop_28_ldst_is_rs1 = _RAND_2417[0:0];
  _RAND_2418 = {1{`RANDOM}};
  rob_uop_28_ldst = _RAND_2418[5:0];
  _RAND_2419 = {1{`RANDOM}};
  rob_uop_28_lrs1 = _RAND_2419[5:0];
  _RAND_2420 = {1{`RANDOM}};
  rob_uop_28_lrs2 = _RAND_2420[5:0];
  _RAND_2421 = {1{`RANDOM}};
  rob_uop_28_lrs3 = _RAND_2421[5:0];
  _RAND_2422 = {1{`RANDOM}};
  rob_uop_28_ldst_val = _RAND_2422[0:0];
  _RAND_2423 = {1{`RANDOM}};
  rob_uop_28_dst_rtype = _RAND_2423[1:0];
  _RAND_2424 = {1{`RANDOM}};
  rob_uop_28_lrs1_rtype = _RAND_2424[1:0];
  _RAND_2425 = {1{`RANDOM}};
  rob_uop_28_lrs2_rtype = _RAND_2425[1:0];
  _RAND_2426 = {1{`RANDOM}};
  rob_uop_28_frs3_en = _RAND_2426[0:0];
  _RAND_2427 = {1{`RANDOM}};
  rob_uop_28_fp_val = _RAND_2427[0:0];
  _RAND_2428 = {1{`RANDOM}};
  rob_uop_28_fp_single = _RAND_2428[0:0];
  _RAND_2429 = {1{`RANDOM}};
  rob_uop_28_xcpt_pf_if = _RAND_2429[0:0];
  _RAND_2430 = {1{`RANDOM}};
  rob_uop_28_xcpt_ae_if = _RAND_2430[0:0];
  _RAND_2431 = {1{`RANDOM}};
  rob_uop_28_xcpt_ma_if = _RAND_2431[0:0];
  _RAND_2432 = {1{`RANDOM}};
  rob_uop_28_bp_debug_if = _RAND_2432[0:0];
  _RAND_2433 = {1{`RANDOM}};
  rob_uop_28_bp_xcpt_if = _RAND_2433[0:0];
  _RAND_2434 = {1{`RANDOM}};
  rob_uop_28_debug_fsrc = _RAND_2434[1:0];
  _RAND_2435 = {1{`RANDOM}};
  rob_uop_28_debug_tsrc = _RAND_2435[1:0];
  _RAND_2436 = {1{`RANDOM}};
  rob_uop_29_uopc = _RAND_2436[6:0];
  _RAND_2437 = {1{`RANDOM}};
  rob_uop_29_inst = _RAND_2437[31:0];
  _RAND_2438 = {1{`RANDOM}};
  rob_uop_29_debug_inst = _RAND_2438[31:0];
  _RAND_2439 = {1{`RANDOM}};
  rob_uop_29_is_rvc = _RAND_2439[0:0];
  _RAND_2440 = {2{`RANDOM}};
  rob_uop_29_debug_pc = _RAND_2440[39:0];
  _RAND_2441 = {1{`RANDOM}};
  rob_uop_29_iq_type = _RAND_2441[2:0];
  _RAND_2442 = {1{`RANDOM}};
  rob_uop_29_fu_code = _RAND_2442[9:0];
  _RAND_2443 = {1{`RANDOM}};
  rob_uop_29_ctrl_br_type = _RAND_2443[3:0];
  _RAND_2444 = {1{`RANDOM}};
  rob_uop_29_ctrl_op1_sel = _RAND_2444[1:0];
  _RAND_2445 = {1{`RANDOM}};
  rob_uop_29_ctrl_op2_sel = _RAND_2445[2:0];
  _RAND_2446 = {1{`RANDOM}};
  rob_uop_29_ctrl_imm_sel = _RAND_2446[2:0];
  _RAND_2447 = {1{`RANDOM}};
  rob_uop_29_ctrl_op_fcn = _RAND_2447[3:0];
  _RAND_2448 = {1{`RANDOM}};
  rob_uop_29_ctrl_fcn_dw = _RAND_2448[0:0];
  _RAND_2449 = {1{`RANDOM}};
  rob_uop_29_ctrl_csr_cmd = _RAND_2449[2:0];
  _RAND_2450 = {1{`RANDOM}};
  rob_uop_29_ctrl_is_load = _RAND_2450[0:0];
  _RAND_2451 = {1{`RANDOM}};
  rob_uop_29_ctrl_is_sta = _RAND_2451[0:0];
  _RAND_2452 = {1{`RANDOM}};
  rob_uop_29_ctrl_is_std = _RAND_2452[0:0];
  _RAND_2453 = {1{`RANDOM}};
  rob_uop_29_iw_state = _RAND_2453[1:0];
  _RAND_2454 = {1{`RANDOM}};
  rob_uop_29_iw_p1_poisoned = _RAND_2454[0:0];
  _RAND_2455 = {1{`RANDOM}};
  rob_uop_29_iw_p2_poisoned = _RAND_2455[0:0];
  _RAND_2456 = {1{`RANDOM}};
  rob_uop_29_is_br = _RAND_2456[0:0];
  _RAND_2457 = {1{`RANDOM}};
  rob_uop_29_is_jalr = _RAND_2457[0:0];
  _RAND_2458 = {1{`RANDOM}};
  rob_uop_29_is_jal = _RAND_2458[0:0];
  _RAND_2459 = {1{`RANDOM}};
  rob_uop_29_is_sfb = _RAND_2459[0:0];
  _RAND_2460 = {1{`RANDOM}};
  rob_uop_29_br_mask = _RAND_2460[7:0];
  _RAND_2461 = {1{`RANDOM}};
  rob_uop_29_br_tag = _RAND_2461[2:0];
  _RAND_2462 = {1{`RANDOM}};
  rob_uop_29_ftq_idx = _RAND_2462[3:0];
  _RAND_2463 = {1{`RANDOM}};
  rob_uop_29_edge_inst = _RAND_2463[0:0];
  _RAND_2464 = {1{`RANDOM}};
  rob_uop_29_pc_lob = _RAND_2464[5:0];
  _RAND_2465 = {1{`RANDOM}};
  rob_uop_29_taken = _RAND_2465[0:0];
  _RAND_2466 = {1{`RANDOM}};
  rob_uop_29_imm_packed = _RAND_2466[19:0];
  _RAND_2467 = {1{`RANDOM}};
  rob_uop_29_csr_addr = _RAND_2467[11:0];
  _RAND_2468 = {1{`RANDOM}};
  rob_uop_29_rob_idx = _RAND_2468[4:0];
  _RAND_2469 = {1{`RANDOM}};
  rob_uop_29_ldq_idx = _RAND_2469[2:0];
  _RAND_2470 = {1{`RANDOM}};
  rob_uop_29_stq_idx = _RAND_2470[2:0];
  _RAND_2471 = {1{`RANDOM}};
  rob_uop_29_rxq_idx = _RAND_2471[1:0];
  _RAND_2472 = {1{`RANDOM}};
  rob_uop_29_pdst = _RAND_2472[5:0];
  _RAND_2473 = {1{`RANDOM}};
  rob_uop_29_prs1 = _RAND_2473[5:0];
  _RAND_2474 = {1{`RANDOM}};
  rob_uop_29_prs2 = _RAND_2474[5:0];
  _RAND_2475 = {1{`RANDOM}};
  rob_uop_29_prs3 = _RAND_2475[5:0];
  _RAND_2476 = {1{`RANDOM}};
  rob_uop_29_ppred = _RAND_2476[3:0];
  _RAND_2477 = {1{`RANDOM}};
  rob_uop_29_prs1_busy = _RAND_2477[0:0];
  _RAND_2478 = {1{`RANDOM}};
  rob_uop_29_prs2_busy = _RAND_2478[0:0];
  _RAND_2479 = {1{`RANDOM}};
  rob_uop_29_prs3_busy = _RAND_2479[0:0];
  _RAND_2480 = {1{`RANDOM}};
  rob_uop_29_ppred_busy = _RAND_2480[0:0];
  _RAND_2481 = {1{`RANDOM}};
  rob_uop_29_stale_pdst = _RAND_2481[5:0];
  _RAND_2482 = {1{`RANDOM}};
  rob_uop_29_exception = _RAND_2482[0:0];
  _RAND_2483 = {2{`RANDOM}};
  rob_uop_29_exc_cause = _RAND_2483[63:0];
  _RAND_2484 = {1{`RANDOM}};
  rob_uop_29_bypassable = _RAND_2484[0:0];
  _RAND_2485 = {1{`RANDOM}};
  rob_uop_29_mem_cmd = _RAND_2485[4:0];
  _RAND_2486 = {1{`RANDOM}};
  rob_uop_29_mem_size = _RAND_2486[1:0];
  _RAND_2487 = {1{`RANDOM}};
  rob_uop_29_mem_signed = _RAND_2487[0:0];
  _RAND_2488 = {1{`RANDOM}};
  rob_uop_29_is_fence = _RAND_2488[0:0];
  _RAND_2489 = {1{`RANDOM}};
  rob_uop_29_is_fencei = _RAND_2489[0:0];
  _RAND_2490 = {1{`RANDOM}};
  rob_uop_29_is_amo = _RAND_2490[0:0];
  _RAND_2491 = {1{`RANDOM}};
  rob_uop_29_uses_ldq = _RAND_2491[0:0];
  _RAND_2492 = {1{`RANDOM}};
  rob_uop_29_uses_stq = _RAND_2492[0:0];
  _RAND_2493 = {1{`RANDOM}};
  rob_uop_29_is_sys_pc2epc = _RAND_2493[0:0];
  _RAND_2494 = {1{`RANDOM}};
  rob_uop_29_is_unique = _RAND_2494[0:0];
  _RAND_2495 = {1{`RANDOM}};
  rob_uop_29_flush_on_commit = _RAND_2495[0:0];
  _RAND_2496 = {1{`RANDOM}};
  rob_uop_29_ldst_is_rs1 = _RAND_2496[0:0];
  _RAND_2497 = {1{`RANDOM}};
  rob_uop_29_ldst = _RAND_2497[5:0];
  _RAND_2498 = {1{`RANDOM}};
  rob_uop_29_lrs1 = _RAND_2498[5:0];
  _RAND_2499 = {1{`RANDOM}};
  rob_uop_29_lrs2 = _RAND_2499[5:0];
  _RAND_2500 = {1{`RANDOM}};
  rob_uop_29_lrs3 = _RAND_2500[5:0];
  _RAND_2501 = {1{`RANDOM}};
  rob_uop_29_ldst_val = _RAND_2501[0:0];
  _RAND_2502 = {1{`RANDOM}};
  rob_uop_29_dst_rtype = _RAND_2502[1:0];
  _RAND_2503 = {1{`RANDOM}};
  rob_uop_29_lrs1_rtype = _RAND_2503[1:0];
  _RAND_2504 = {1{`RANDOM}};
  rob_uop_29_lrs2_rtype = _RAND_2504[1:0];
  _RAND_2505 = {1{`RANDOM}};
  rob_uop_29_frs3_en = _RAND_2505[0:0];
  _RAND_2506 = {1{`RANDOM}};
  rob_uop_29_fp_val = _RAND_2506[0:0];
  _RAND_2507 = {1{`RANDOM}};
  rob_uop_29_fp_single = _RAND_2507[0:0];
  _RAND_2508 = {1{`RANDOM}};
  rob_uop_29_xcpt_pf_if = _RAND_2508[0:0];
  _RAND_2509 = {1{`RANDOM}};
  rob_uop_29_xcpt_ae_if = _RAND_2509[0:0];
  _RAND_2510 = {1{`RANDOM}};
  rob_uop_29_xcpt_ma_if = _RAND_2510[0:0];
  _RAND_2511 = {1{`RANDOM}};
  rob_uop_29_bp_debug_if = _RAND_2511[0:0];
  _RAND_2512 = {1{`RANDOM}};
  rob_uop_29_bp_xcpt_if = _RAND_2512[0:0];
  _RAND_2513 = {1{`RANDOM}};
  rob_uop_29_debug_fsrc = _RAND_2513[1:0];
  _RAND_2514 = {1{`RANDOM}};
  rob_uop_29_debug_tsrc = _RAND_2514[1:0];
  _RAND_2515 = {1{`RANDOM}};
  rob_uop_30_uopc = _RAND_2515[6:0];
  _RAND_2516 = {1{`RANDOM}};
  rob_uop_30_inst = _RAND_2516[31:0];
  _RAND_2517 = {1{`RANDOM}};
  rob_uop_30_debug_inst = _RAND_2517[31:0];
  _RAND_2518 = {1{`RANDOM}};
  rob_uop_30_is_rvc = _RAND_2518[0:0];
  _RAND_2519 = {2{`RANDOM}};
  rob_uop_30_debug_pc = _RAND_2519[39:0];
  _RAND_2520 = {1{`RANDOM}};
  rob_uop_30_iq_type = _RAND_2520[2:0];
  _RAND_2521 = {1{`RANDOM}};
  rob_uop_30_fu_code = _RAND_2521[9:0];
  _RAND_2522 = {1{`RANDOM}};
  rob_uop_30_ctrl_br_type = _RAND_2522[3:0];
  _RAND_2523 = {1{`RANDOM}};
  rob_uop_30_ctrl_op1_sel = _RAND_2523[1:0];
  _RAND_2524 = {1{`RANDOM}};
  rob_uop_30_ctrl_op2_sel = _RAND_2524[2:0];
  _RAND_2525 = {1{`RANDOM}};
  rob_uop_30_ctrl_imm_sel = _RAND_2525[2:0];
  _RAND_2526 = {1{`RANDOM}};
  rob_uop_30_ctrl_op_fcn = _RAND_2526[3:0];
  _RAND_2527 = {1{`RANDOM}};
  rob_uop_30_ctrl_fcn_dw = _RAND_2527[0:0];
  _RAND_2528 = {1{`RANDOM}};
  rob_uop_30_ctrl_csr_cmd = _RAND_2528[2:0];
  _RAND_2529 = {1{`RANDOM}};
  rob_uop_30_ctrl_is_load = _RAND_2529[0:0];
  _RAND_2530 = {1{`RANDOM}};
  rob_uop_30_ctrl_is_sta = _RAND_2530[0:0];
  _RAND_2531 = {1{`RANDOM}};
  rob_uop_30_ctrl_is_std = _RAND_2531[0:0];
  _RAND_2532 = {1{`RANDOM}};
  rob_uop_30_iw_state = _RAND_2532[1:0];
  _RAND_2533 = {1{`RANDOM}};
  rob_uop_30_iw_p1_poisoned = _RAND_2533[0:0];
  _RAND_2534 = {1{`RANDOM}};
  rob_uop_30_iw_p2_poisoned = _RAND_2534[0:0];
  _RAND_2535 = {1{`RANDOM}};
  rob_uop_30_is_br = _RAND_2535[0:0];
  _RAND_2536 = {1{`RANDOM}};
  rob_uop_30_is_jalr = _RAND_2536[0:0];
  _RAND_2537 = {1{`RANDOM}};
  rob_uop_30_is_jal = _RAND_2537[0:0];
  _RAND_2538 = {1{`RANDOM}};
  rob_uop_30_is_sfb = _RAND_2538[0:0];
  _RAND_2539 = {1{`RANDOM}};
  rob_uop_30_br_mask = _RAND_2539[7:0];
  _RAND_2540 = {1{`RANDOM}};
  rob_uop_30_br_tag = _RAND_2540[2:0];
  _RAND_2541 = {1{`RANDOM}};
  rob_uop_30_ftq_idx = _RAND_2541[3:0];
  _RAND_2542 = {1{`RANDOM}};
  rob_uop_30_edge_inst = _RAND_2542[0:0];
  _RAND_2543 = {1{`RANDOM}};
  rob_uop_30_pc_lob = _RAND_2543[5:0];
  _RAND_2544 = {1{`RANDOM}};
  rob_uop_30_taken = _RAND_2544[0:0];
  _RAND_2545 = {1{`RANDOM}};
  rob_uop_30_imm_packed = _RAND_2545[19:0];
  _RAND_2546 = {1{`RANDOM}};
  rob_uop_30_csr_addr = _RAND_2546[11:0];
  _RAND_2547 = {1{`RANDOM}};
  rob_uop_30_rob_idx = _RAND_2547[4:0];
  _RAND_2548 = {1{`RANDOM}};
  rob_uop_30_ldq_idx = _RAND_2548[2:0];
  _RAND_2549 = {1{`RANDOM}};
  rob_uop_30_stq_idx = _RAND_2549[2:0];
  _RAND_2550 = {1{`RANDOM}};
  rob_uop_30_rxq_idx = _RAND_2550[1:0];
  _RAND_2551 = {1{`RANDOM}};
  rob_uop_30_pdst = _RAND_2551[5:0];
  _RAND_2552 = {1{`RANDOM}};
  rob_uop_30_prs1 = _RAND_2552[5:0];
  _RAND_2553 = {1{`RANDOM}};
  rob_uop_30_prs2 = _RAND_2553[5:0];
  _RAND_2554 = {1{`RANDOM}};
  rob_uop_30_prs3 = _RAND_2554[5:0];
  _RAND_2555 = {1{`RANDOM}};
  rob_uop_30_ppred = _RAND_2555[3:0];
  _RAND_2556 = {1{`RANDOM}};
  rob_uop_30_prs1_busy = _RAND_2556[0:0];
  _RAND_2557 = {1{`RANDOM}};
  rob_uop_30_prs2_busy = _RAND_2557[0:0];
  _RAND_2558 = {1{`RANDOM}};
  rob_uop_30_prs3_busy = _RAND_2558[0:0];
  _RAND_2559 = {1{`RANDOM}};
  rob_uop_30_ppred_busy = _RAND_2559[0:0];
  _RAND_2560 = {1{`RANDOM}};
  rob_uop_30_stale_pdst = _RAND_2560[5:0];
  _RAND_2561 = {1{`RANDOM}};
  rob_uop_30_exception = _RAND_2561[0:0];
  _RAND_2562 = {2{`RANDOM}};
  rob_uop_30_exc_cause = _RAND_2562[63:0];
  _RAND_2563 = {1{`RANDOM}};
  rob_uop_30_bypassable = _RAND_2563[0:0];
  _RAND_2564 = {1{`RANDOM}};
  rob_uop_30_mem_cmd = _RAND_2564[4:0];
  _RAND_2565 = {1{`RANDOM}};
  rob_uop_30_mem_size = _RAND_2565[1:0];
  _RAND_2566 = {1{`RANDOM}};
  rob_uop_30_mem_signed = _RAND_2566[0:0];
  _RAND_2567 = {1{`RANDOM}};
  rob_uop_30_is_fence = _RAND_2567[0:0];
  _RAND_2568 = {1{`RANDOM}};
  rob_uop_30_is_fencei = _RAND_2568[0:0];
  _RAND_2569 = {1{`RANDOM}};
  rob_uop_30_is_amo = _RAND_2569[0:0];
  _RAND_2570 = {1{`RANDOM}};
  rob_uop_30_uses_ldq = _RAND_2570[0:0];
  _RAND_2571 = {1{`RANDOM}};
  rob_uop_30_uses_stq = _RAND_2571[0:0];
  _RAND_2572 = {1{`RANDOM}};
  rob_uop_30_is_sys_pc2epc = _RAND_2572[0:0];
  _RAND_2573 = {1{`RANDOM}};
  rob_uop_30_is_unique = _RAND_2573[0:0];
  _RAND_2574 = {1{`RANDOM}};
  rob_uop_30_flush_on_commit = _RAND_2574[0:0];
  _RAND_2575 = {1{`RANDOM}};
  rob_uop_30_ldst_is_rs1 = _RAND_2575[0:0];
  _RAND_2576 = {1{`RANDOM}};
  rob_uop_30_ldst = _RAND_2576[5:0];
  _RAND_2577 = {1{`RANDOM}};
  rob_uop_30_lrs1 = _RAND_2577[5:0];
  _RAND_2578 = {1{`RANDOM}};
  rob_uop_30_lrs2 = _RAND_2578[5:0];
  _RAND_2579 = {1{`RANDOM}};
  rob_uop_30_lrs3 = _RAND_2579[5:0];
  _RAND_2580 = {1{`RANDOM}};
  rob_uop_30_ldst_val = _RAND_2580[0:0];
  _RAND_2581 = {1{`RANDOM}};
  rob_uop_30_dst_rtype = _RAND_2581[1:0];
  _RAND_2582 = {1{`RANDOM}};
  rob_uop_30_lrs1_rtype = _RAND_2582[1:0];
  _RAND_2583 = {1{`RANDOM}};
  rob_uop_30_lrs2_rtype = _RAND_2583[1:0];
  _RAND_2584 = {1{`RANDOM}};
  rob_uop_30_frs3_en = _RAND_2584[0:0];
  _RAND_2585 = {1{`RANDOM}};
  rob_uop_30_fp_val = _RAND_2585[0:0];
  _RAND_2586 = {1{`RANDOM}};
  rob_uop_30_fp_single = _RAND_2586[0:0];
  _RAND_2587 = {1{`RANDOM}};
  rob_uop_30_xcpt_pf_if = _RAND_2587[0:0];
  _RAND_2588 = {1{`RANDOM}};
  rob_uop_30_xcpt_ae_if = _RAND_2588[0:0];
  _RAND_2589 = {1{`RANDOM}};
  rob_uop_30_xcpt_ma_if = _RAND_2589[0:0];
  _RAND_2590 = {1{`RANDOM}};
  rob_uop_30_bp_debug_if = _RAND_2590[0:0];
  _RAND_2591 = {1{`RANDOM}};
  rob_uop_30_bp_xcpt_if = _RAND_2591[0:0];
  _RAND_2592 = {1{`RANDOM}};
  rob_uop_30_debug_fsrc = _RAND_2592[1:0];
  _RAND_2593 = {1{`RANDOM}};
  rob_uop_30_debug_tsrc = _RAND_2593[1:0];
  _RAND_2594 = {1{`RANDOM}};
  rob_uop_31_uopc = _RAND_2594[6:0];
  _RAND_2595 = {1{`RANDOM}};
  rob_uop_31_inst = _RAND_2595[31:0];
  _RAND_2596 = {1{`RANDOM}};
  rob_uop_31_debug_inst = _RAND_2596[31:0];
  _RAND_2597 = {1{`RANDOM}};
  rob_uop_31_is_rvc = _RAND_2597[0:0];
  _RAND_2598 = {2{`RANDOM}};
  rob_uop_31_debug_pc = _RAND_2598[39:0];
  _RAND_2599 = {1{`RANDOM}};
  rob_uop_31_iq_type = _RAND_2599[2:0];
  _RAND_2600 = {1{`RANDOM}};
  rob_uop_31_fu_code = _RAND_2600[9:0];
  _RAND_2601 = {1{`RANDOM}};
  rob_uop_31_ctrl_br_type = _RAND_2601[3:0];
  _RAND_2602 = {1{`RANDOM}};
  rob_uop_31_ctrl_op1_sel = _RAND_2602[1:0];
  _RAND_2603 = {1{`RANDOM}};
  rob_uop_31_ctrl_op2_sel = _RAND_2603[2:0];
  _RAND_2604 = {1{`RANDOM}};
  rob_uop_31_ctrl_imm_sel = _RAND_2604[2:0];
  _RAND_2605 = {1{`RANDOM}};
  rob_uop_31_ctrl_op_fcn = _RAND_2605[3:0];
  _RAND_2606 = {1{`RANDOM}};
  rob_uop_31_ctrl_fcn_dw = _RAND_2606[0:0];
  _RAND_2607 = {1{`RANDOM}};
  rob_uop_31_ctrl_csr_cmd = _RAND_2607[2:0];
  _RAND_2608 = {1{`RANDOM}};
  rob_uop_31_ctrl_is_load = _RAND_2608[0:0];
  _RAND_2609 = {1{`RANDOM}};
  rob_uop_31_ctrl_is_sta = _RAND_2609[0:0];
  _RAND_2610 = {1{`RANDOM}};
  rob_uop_31_ctrl_is_std = _RAND_2610[0:0];
  _RAND_2611 = {1{`RANDOM}};
  rob_uop_31_iw_state = _RAND_2611[1:0];
  _RAND_2612 = {1{`RANDOM}};
  rob_uop_31_iw_p1_poisoned = _RAND_2612[0:0];
  _RAND_2613 = {1{`RANDOM}};
  rob_uop_31_iw_p2_poisoned = _RAND_2613[0:0];
  _RAND_2614 = {1{`RANDOM}};
  rob_uop_31_is_br = _RAND_2614[0:0];
  _RAND_2615 = {1{`RANDOM}};
  rob_uop_31_is_jalr = _RAND_2615[0:0];
  _RAND_2616 = {1{`RANDOM}};
  rob_uop_31_is_jal = _RAND_2616[0:0];
  _RAND_2617 = {1{`RANDOM}};
  rob_uop_31_is_sfb = _RAND_2617[0:0];
  _RAND_2618 = {1{`RANDOM}};
  rob_uop_31_br_mask = _RAND_2618[7:0];
  _RAND_2619 = {1{`RANDOM}};
  rob_uop_31_br_tag = _RAND_2619[2:0];
  _RAND_2620 = {1{`RANDOM}};
  rob_uop_31_ftq_idx = _RAND_2620[3:0];
  _RAND_2621 = {1{`RANDOM}};
  rob_uop_31_edge_inst = _RAND_2621[0:0];
  _RAND_2622 = {1{`RANDOM}};
  rob_uop_31_pc_lob = _RAND_2622[5:0];
  _RAND_2623 = {1{`RANDOM}};
  rob_uop_31_taken = _RAND_2623[0:0];
  _RAND_2624 = {1{`RANDOM}};
  rob_uop_31_imm_packed = _RAND_2624[19:0];
  _RAND_2625 = {1{`RANDOM}};
  rob_uop_31_csr_addr = _RAND_2625[11:0];
  _RAND_2626 = {1{`RANDOM}};
  rob_uop_31_rob_idx = _RAND_2626[4:0];
  _RAND_2627 = {1{`RANDOM}};
  rob_uop_31_ldq_idx = _RAND_2627[2:0];
  _RAND_2628 = {1{`RANDOM}};
  rob_uop_31_stq_idx = _RAND_2628[2:0];
  _RAND_2629 = {1{`RANDOM}};
  rob_uop_31_rxq_idx = _RAND_2629[1:0];
  _RAND_2630 = {1{`RANDOM}};
  rob_uop_31_pdst = _RAND_2630[5:0];
  _RAND_2631 = {1{`RANDOM}};
  rob_uop_31_prs1 = _RAND_2631[5:0];
  _RAND_2632 = {1{`RANDOM}};
  rob_uop_31_prs2 = _RAND_2632[5:0];
  _RAND_2633 = {1{`RANDOM}};
  rob_uop_31_prs3 = _RAND_2633[5:0];
  _RAND_2634 = {1{`RANDOM}};
  rob_uop_31_ppred = _RAND_2634[3:0];
  _RAND_2635 = {1{`RANDOM}};
  rob_uop_31_prs1_busy = _RAND_2635[0:0];
  _RAND_2636 = {1{`RANDOM}};
  rob_uop_31_prs2_busy = _RAND_2636[0:0];
  _RAND_2637 = {1{`RANDOM}};
  rob_uop_31_prs3_busy = _RAND_2637[0:0];
  _RAND_2638 = {1{`RANDOM}};
  rob_uop_31_ppred_busy = _RAND_2638[0:0];
  _RAND_2639 = {1{`RANDOM}};
  rob_uop_31_stale_pdst = _RAND_2639[5:0];
  _RAND_2640 = {1{`RANDOM}};
  rob_uop_31_exception = _RAND_2640[0:0];
  _RAND_2641 = {2{`RANDOM}};
  rob_uop_31_exc_cause = _RAND_2641[63:0];
  _RAND_2642 = {1{`RANDOM}};
  rob_uop_31_bypassable = _RAND_2642[0:0];
  _RAND_2643 = {1{`RANDOM}};
  rob_uop_31_mem_cmd = _RAND_2643[4:0];
  _RAND_2644 = {1{`RANDOM}};
  rob_uop_31_mem_size = _RAND_2644[1:0];
  _RAND_2645 = {1{`RANDOM}};
  rob_uop_31_mem_signed = _RAND_2645[0:0];
  _RAND_2646 = {1{`RANDOM}};
  rob_uop_31_is_fence = _RAND_2646[0:0];
  _RAND_2647 = {1{`RANDOM}};
  rob_uop_31_is_fencei = _RAND_2647[0:0];
  _RAND_2648 = {1{`RANDOM}};
  rob_uop_31_is_amo = _RAND_2648[0:0];
  _RAND_2649 = {1{`RANDOM}};
  rob_uop_31_uses_ldq = _RAND_2649[0:0];
  _RAND_2650 = {1{`RANDOM}};
  rob_uop_31_uses_stq = _RAND_2650[0:0];
  _RAND_2651 = {1{`RANDOM}};
  rob_uop_31_is_sys_pc2epc = _RAND_2651[0:0];
  _RAND_2652 = {1{`RANDOM}};
  rob_uop_31_is_unique = _RAND_2652[0:0];
  _RAND_2653 = {1{`RANDOM}};
  rob_uop_31_flush_on_commit = _RAND_2653[0:0];
  _RAND_2654 = {1{`RANDOM}};
  rob_uop_31_ldst_is_rs1 = _RAND_2654[0:0];
  _RAND_2655 = {1{`RANDOM}};
  rob_uop_31_ldst = _RAND_2655[5:0];
  _RAND_2656 = {1{`RANDOM}};
  rob_uop_31_lrs1 = _RAND_2656[5:0];
  _RAND_2657 = {1{`RANDOM}};
  rob_uop_31_lrs2 = _RAND_2657[5:0];
  _RAND_2658 = {1{`RANDOM}};
  rob_uop_31_lrs3 = _RAND_2658[5:0];
  _RAND_2659 = {1{`RANDOM}};
  rob_uop_31_ldst_val = _RAND_2659[0:0];
  _RAND_2660 = {1{`RANDOM}};
  rob_uop_31_dst_rtype = _RAND_2660[1:0];
  _RAND_2661 = {1{`RANDOM}};
  rob_uop_31_lrs1_rtype = _RAND_2661[1:0];
  _RAND_2662 = {1{`RANDOM}};
  rob_uop_31_lrs2_rtype = _RAND_2662[1:0];
  _RAND_2663 = {1{`RANDOM}};
  rob_uop_31_frs3_en = _RAND_2663[0:0];
  _RAND_2664 = {1{`RANDOM}};
  rob_uop_31_fp_val = _RAND_2664[0:0];
  _RAND_2665 = {1{`RANDOM}};
  rob_uop_31_fp_single = _RAND_2665[0:0];
  _RAND_2666 = {1{`RANDOM}};
  rob_uop_31_xcpt_pf_if = _RAND_2666[0:0];
  _RAND_2667 = {1{`RANDOM}};
  rob_uop_31_xcpt_ae_if = _RAND_2667[0:0];
  _RAND_2668 = {1{`RANDOM}};
  rob_uop_31_xcpt_ma_if = _RAND_2668[0:0];
  _RAND_2669 = {1{`RANDOM}};
  rob_uop_31_bp_debug_if = _RAND_2669[0:0];
  _RAND_2670 = {1{`RANDOM}};
  rob_uop_31_bp_xcpt_if = _RAND_2670[0:0];
  _RAND_2671 = {1{`RANDOM}};
  rob_uop_31_debug_fsrc = _RAND_2671[1:0];
  _RAND_2672 = {1{`RANDOM}};
  rob_uop_31_debug_tsrc = _RAND_2672[1:0];
  _RAND_2673 = {1{`RANDOM}};
  rob_predicated_0 = _RAND_2673[0:0];
  _RAND_2674 = {1{`RANDOM}};
  rob_predicated_1 = _RAND_2674[0:0];
  _RAND_2675 = {1{`RANDOM}};
  rob_predicated_2 = _RAND_2675[0:0];
  _RAND_2676 = {1{`RANDOM}};
  rob_predicated_3 = _RAND_2676[0:0];
  _RAND_2677 = {1{`RANDOM}};
  rob_predicated_4 = _RAND_2677[0:0];
  _RAND_2678 = {1{`RANDOM}};
  rob_predicated_5 = _RAND_2678[0:0];
  _RAND_2679 = {1{`RANDOM}};
  rob_predicated_6 = _RAND_2679[0:0];
  _RAND_2680 = {1{`RANDOM}};
  rob_predicated_7 = _RAND_2680[0:0];
  _RAND_2681 = {1{`RANDOM}};
  rob_predicated_8 = _RAND_2681[0:0];
  _RAND_2682 = {1{`RANDOM}};
  rob_predicated_9 = _RAND_2682[0:0];
  _RAND_2683 = {1{`RANDOM}};
  rob_predicated_10 = _RAND_2683[0:0];
  _RAND_2684 = {1{`RANDOM}};
  rob_predicated_11 = _RAND_2684[0:0];
  _RAND_2685 = {1{`RANDOM}};
  rob_predicated_12 = _RAND_2685[0:0];
  _RAND_2686 = {1{`RANDOM}};
  rob_predicated_13 = _RAND_2686[0:0];
  _RAND_2687 = {1{`RANDOM}};
  rob_predicated_14 = _RAND_2687[0:0];
  _RAND_2688 = {1{`RANDOM}};
  rob_predicated_15 = _RAND_2688[0:0];
  _RAND_2689 = {1{`RANDOM}};
  rob_predicated_16 = _RAND_2689[0:0];
  _RAND_2690 = {1{`RANDOM}};
  rob_predicated_17 = _RAND_2690[0:0];
  _RAND_2691 = {1{`RANDOM}};
  rob_predicated_18 = _RAND_2691[0:0];
  _RAND_2692 = {1{`RANDOM}};
  rob_predicated_19 = _RAND_2692[0:0];
  _RAND_2693 = {1{`RANDOM}};
  rob_predicated_20 = _RAND_2693[0:0];
  _RAND_2694 = {1{`RANDOM}};
  rob_predicated_21 = _RAND_2694[0:0];
  _RAND_2695 = {1{`RANDOM}};
  rob_predicated_22 = _RAND_2695[0:0];
  _RAND_2696 = {1{`RANDOM}};
  rob_predicated_23 = _RAND_2696[0:0];
  _RAND_2697 = {1{`RANDOM}};
  rob_predicated_24 = _RAND_2697[0:0];
  _RAND_2698 = {1{`RANDOM}};
  rob_predicated_25 = _RAND_2698[0:0];
  _RAND_2699 = {1{`RANDOM}};
  rob_predicated_26 = _RAND_2699[0:0];
  _RAND_2700 = {1{`RANDOM}};
  rob_predicated_27 = _RAND_2700[0:0];
  _RAND_2701 = {1{`RANDOM}};
  rob_predicated_28 = _RAND_2701[0:0];
  _RAND_2702 = {1{`RANDOM}};
  rob_predicated_29 = _RAND_2702[0:0];
  _RAND_2703 = {1{`RANDOM}};
  rob_predicated_30 = _RAND_2703[0:0];
  _RAND_2704 = {1{`RANDOM}};
  rob_predicated_31 = _RAND_2704[0:0];
  _RAND_2705 = {1{`RANDOM}};
  _T_406 = _RAND_2705[0:0];
  _RAND_2706 = {1{`RANDOM}};
  r_partial_row = _RAND_2706[0:0];
  _RAND_2707 = {1{`RANDOM}};
  pnr_maybe_at_tail = _RAND_2707[0:0];
  _RAND_2708 = {1{`RANDOM}};
  _T_609 = _RAND_2708[0:0];
  _RAND_2709 = {1{`RANDOM}};
  _T_610 = _RAND_2709[0:0];
  _RAND_2710 = {1{`RANDOM}};
  _T_614 = _RAND_2710[0:0];
  _RAND_2711 = {1{`RANDOM}};
  _T_618 = _RAND_2711[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
