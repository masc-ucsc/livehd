module hier_tuple2 (
  output [3:0] out,
);

assign out  = 4'd12;

endmodule 
