module scalar_tuple (
  output [1:0] out,
  output [1:0] out2
);

assign out = 2'd3;
assign out2 = 2'd3;

endmodule
