module FlipSimple3(
  output  io_in_ab,
  input   io_out_ab
);
  assign io_in_ab = io_out_ab;
endmodule
