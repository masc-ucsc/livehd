module trivial( input [3:0] a, input [3:0] b, output [3:0] c, output [3:0] d);
assign c = a + b;
assign d = a - b;
endmodule

