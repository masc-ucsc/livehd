module hier_tuple (
  output [1:0] out,
  output [2:0] out2,
  output [2:0] out3
);

assign out  = 2'd3;
assign out2 = 3'd5;
assign out3 = 3'd6;

endmodule 
