module tuple_nested1(
   output reg signed [5:0] out
);
always @(*) begin
  out = 25;
end
endmodule
