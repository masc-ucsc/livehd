module sum1( input [1:0] a, output [3:0] c);
assign c = a + 1'b1;
endmodule

