module attr_set (
  output [1:0] out
);

assign out = 2'd2;

endmodule 
