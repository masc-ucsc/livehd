module trivialx( input a, input [1:0] b, output c);
assign c = a & b;
endmodule

