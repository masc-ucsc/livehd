module funcall4 (
  output [4:0] out
);

assign out = 5'd15;

endmodule
