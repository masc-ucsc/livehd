module tup_out2 (
  output [1:0] out_a
);

  assign out_a = 2'h1;

endmodule
