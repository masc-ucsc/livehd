module sum1( input a, output [2:0] c);
assign c = a + 1'b1;
endmodule

