module capricious_bits (
  output [3:0] out
);

assign out = 4'd9;

endmodule
