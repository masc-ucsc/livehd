

module blackbox(input a, input b, output c);

  undefined_potato potato1(.a(a), .b(b), .c(c));

endmodule

