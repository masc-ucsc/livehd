module bits_rhs (
  output [6:0] out
);

assign out = {4'd8,3'd5};

endmodule 
