module testing;
  input a, b;
  output unsigned c, d;
  inout unsigned [LENGTH-1:0] e, f;
  input [WIDTH-1:0] g, h;
  output reg signed i, j;
  inout unsigned tri k, l;
  input unsigned wire [BREADTH-1:0] m, n;
  output reg [NUMBER-1:0] o, p;


  wire aa;
  wire signed [WORD-1:0][ANOTHER:23] bb, cc;
  reg [DIM1:99] [DIM2:234857] dd [DIM3:0][DIM4:0], ee[DIM5:0];
endmodule
