module capricious_bits4 (
  output [4:0] out,
  output [4:0] out2,
);

  assign out = 5'h17;
  assign out2 = 15;

endmodule
