module tuple_empty_attr (
  output out,
  output [2:0] out2
);

assign out = 1'd0;
assign out2 = 3'd3;

endmodule
