VERSION 5.8 ;

BUSBITCHARS "[]" ;

DIVIDERCHAR "/" ;

UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.000500 ;

CLEARANCEMEASURE EUCLIDEAN ;
USEMINSPACING OBS ON ;

SITE CoreSite
    CLASS CORE ;
    SIZE 0.200000 BY 1.710000 ; 
END CoreSite

LAYER Metal1
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    MINWIDTH 0.060000 ;
    AREA 0.020000 ;
    WIDTH 0.060000 ;
    SPACING 0.060000 ;
    SPACING 0.090000 ENDOFLINE 0.090000 WITHIN 0.025000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.060000
      WIDTH  0.100000  0.100000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.190000 0.190000 ;
END Metal1

LAYER Via1
    TYPE CUT ;
    SPACING 0.070000 ;
    WIDTH 0.06 ;
END Via1

LAYER Metal2
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    MINWIDTH 0.070000 ;
    AREA 0.020000 ;
    WIDTH 0.070000 ;
    SPACING 0.070000 ;
    SPACING 0.100000 ENDOFLINE 0.100000 WITHIN 0.035000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.070000
      WIDTH  0.100000  0.150000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.200000 0.200000 ;
END Metal2

LAYER Via2
    TYPE CUT ;
    SPACING 0.070000 ;
    WIDTH 0.07 ;
END Via2

LAYER Metal3
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    MINWIDTH 0.070000 ;
    AREA 0.020000 ;
    WIDTH 0.070000 ;
    SPACING 0.070000 ;
    SPACING 0.100000 ENDOFLINE 0.100000 WITHIN 0.035000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.070000
      WIDTH  0.100000  0.150000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.200000 0.200000 ;
END Metal3

LAYER Via3
    TYPE CUT ;
    SPACING 0.070000 ;
    WIDTH 0.07 ;
END Via3

LAYER Metal4
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    MINWIDTH 0.070000 ;
    AREA 0.020000 ;
    WIDTH 0.070000 ;
    SPACING 0.070000 ;
    SPACING 0.100000 ENDOFLINE 0.100000 WITHIN 0.035000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.070000
      WIDTH  0.100000  0.150000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.200000 0.200000 ;
END Metal4

LAYER Via4
    TYPE CUT ;
    SPACING 0.070000 ;
    WIDTH 0.07 ;
END Via4

LAYER Metal5
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    MINWIDTH 0.070000 ;
    AREA 0.020000 ;
    WIDTH 0.070000 ;
    SPACING 0.070000 ;
    SPACING 0.100000 ENDOFLINE 0.100000 WITHIN 0.035000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.070000
      WIDTH  0.100000  0.150000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.200000 0.200000 ;
END Metal5

LAYER Via5
    TYPE CUT ;
    SPACING 0.070000 ;
    WIDTH 0.07 ;
END Via5

LAYER Metal6
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    MINWIDTH 0.070000 ;
    AREA 0.020000 ;
    WIDTH 0.070000 ;
    SPACING 0.070000 ;
    SPACING 0.100000 ENDOFLINE 0.100000 WITHIN 0.035000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.070000
      WIDTH  0.100000  0.150000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.200000 0.200000 ;
END Metal6

LAYER Via6
    TYPE CUT ;
    SPACING 0.070000 ;
    WIDTH 0.07 ;
END Via6

LAYER Metal7
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    MINWIDTH 0.070000 ;
    AREA 0.020000 ;
    WIDTH 0.070000 ;
    SPACING 0.070000 ;
    SPACING 0.100000 ENDOFLINE 0.100000 WITHIN 0.035000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.070000
      WIDTH  0.100000  0.150000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.200000 0.200000 ;
END Metal7

LAYER Via7
    TYPE CUT ;
    SPACING 0.070000 ;
    WIDTH 0.07 ;
END Via7

LAYER Metal8
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    MINWIDTH 0.070000 ;
    AREA 0.020000 ;
    WIDTH 0.070000 ;
    SPACING 0.070000 ;
    SPACING 0.100000 ENDOFLINE 0.100000 WITHIN 0.035000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.070000
      WIDTH  0.100000  0.150000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.200000 0.200000 ;
END Metal8

LAYER Via8
    TYPE CUT ;
    SPACING 0.070000 ;
    WIDTH 0.07 ;
END Via8

LAYER Metal9
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    MINWIDTH 0.070000 ;
    AREA 0.020000 ;
    WIDTH 0.070000 ;
    SPACING 0.070000 ;
    SPACING 0.100000 ENDOFLINE 0.100000 WITHIN 0.035000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.070000
      WIDTH  0.100000  0.150000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.330000 0.330000 ;
END Metal9

LAYER OVERLAP
    TYPE OVERLAP ;
END OVERLAP

VIA VIA12_1C DEFAULT 
    LAYER Metal1 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via1 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal2 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA12_1C

VIA VIA12_1C_H DEFAULT 
    LAYER Metal1 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via1 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal2 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA12_1C_H

VIA VIA12_1C_V DEFAULT 
    LAYER Metal1 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via1 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal2 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA12_1C_V

VIA VIA23_1C DEFAULT 
    LAYER Metal2 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA23_1C

VIA VIA23_1C_H DEFAULT 
    LAYER Metal2 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA23_1C_H

VIA VIA23_1C_V DEFAULT 
    LAYER Metal2 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal3 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA23_1C_V

VIA VIA23_1ST_N DEFAULT 
    LAYER Metal2 ;
        RECT -0.035000 -0.065000 0.035000 0.325000 ;
    LAYER Via2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA23_1ST_N

VIA VIA23_1ST_S DEFAULT 
    LAYER Metal2 ;
        RECT -0.035000 -0.325000 0.035000 0.065000 ;
    LAYER Via2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA23_1ST_S

VIA VIA34_1C DEFAULT 
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA34_1C

VIA VIA34_1C_H DEFAULT 
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal4 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA34_1C_H

VIA VIA34_1C_V DEFAULT 
    LAYER Metal3 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA34_1C_V

VIA VIA34_1ST_E DEFAULT 
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.325000 0.035000 ;
    LAYER Via3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA34_1ST_E

VIA VIA34_1ST_W DEFAULT 
    LAYER Metal3 ;
        RECT -0.325000 -0.035000 0.065000 0.035000 ;
    LAYER Via3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA34_1ST_W

VIA VIA45_1C DEFAULT 
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal5 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA45_1C

VIA VIA45_1C_H DEFAULT 
    LAYER Metal4 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal5 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA45_1C_H

VIA VIA45_1C_V DEFAULT 
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal5 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA45_1C_V

VIA VIA45_1ST_N DEFAULT 
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.325000 ;
    LAYER Via4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal5 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA45_1ST_N

VIA VIA45_1ST_S DEFAULT 
    LAYER Metal4 ;
        RECT -0.035000 -0.325000 0.035000 0.065000 ;
    LAYER Via4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal5 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA45_1ST_S

VIA VIA5_0_VH DEFAULT 
    LAYER Metal5 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via5 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal6 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA5_0_VH

VIA VIA6_0_HV DEFAULT 
    LAYER Metal6 ;
        RECT -0.260000 -0.200000 0.260000 0.200000 ;
    LAYER Via6 ;
        RECT -0.180000 -0.180000 0.180000 0.180000 ;
    LAYER Metal7 ;
        RECT -0.200000 -0.260000 0.200000 0.260000 ;
END VIA6_0_HV

VIA VIA7_0_VH DEFAULT 
    LAYER Metal7 ;
        RECT -0.200000 -0.260000 0.200000 0.260000 ;
    LAYER Via7 ;
        RECT -0.180000 -0.180000 0.180000 0.180000 ;
    LAYER Metal8 ;
        RECT -0.260000 -0.200000 0.260000 0.200000 ;
END VIA7_0_VH

VIA VIA8_0_VH DEFAULT 
    LAYER Metal8 ;
        RECT -0.200000 -0.260000 0.200000 0.260000 ;
    LAYER Via8 ;
        RECT -0.180000 -0.180000 0.180000 0.180000 ;
    LAYER Metal9 ;
        RECT -0.260000 -0.200000 0.260000 0.200000 ;
END VIA8_0_VH


MACRO AOI221X2
    CLASS CORE ;
    FOREIGN AOI221X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.600000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.235000 0.625000 0.365000 0.715000 ;
        RECT 0.285000 0.610000 0.960000 0.690000 ;
        RECT 0.285000 0.610000 0.365000 0.715000 ;
        RECT 0.235000 0.625000 0.960000 0.690000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.660000 0.765000 0.740000 1.065000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.635000 0.625000 1.765000 0.715000 ;
        RECT 1.240000 0.635000 1.935000 0.715000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.435000 0.815000 1.935000 0.895000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.065000 0.815000 2.565000 0.895000 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 2.600000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 2.600000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.060000 0.790000 1.140000 0.920000 ;
        RECT 2.220000 0.995000 2.280000 1.135000 ;
        RECT 1.080000 0.995000 2.280000 1.055000 ;
        RECT 1.080000 0.450000 1.140000 1.055000 ;
        RECT 0.605000 0.450000 2.170000 0.510000 ;
        END
    END Y
END AOI221X2

MACRO NAND3X2
    CLASS CORE ;
    FOREIGN NAND3X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.260000 0.600000 0.370000 0.735000 ;
        RECT 1.240000 0.495000 1.300000 0.735000 ;
        RECT 0.310000 0.495000 1.300000 0.555000 ;
        RECT 0.310000 0.495000 0.370000 0.735000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.060000 0.655000 1.140000 0.920000 ;
        RECT 0.470000 0.655000 1.140000 0.715000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.520000 0.815000 0.765000 0.955000 ;
        RECT 0.520000 0.815000 0.960000 0.895000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 1.600000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 1.600000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.435000 1.005000 1.565000 1.115000 ;
        RECT 0.360000 1.055000 0.430000 1.335000 ;
        RECT 1.505000 0.335000 1.565000 1.115000 ;
        RECT 1.190000 1.055000 1.250000 1.335000 ;
        RECT 0.795000 0.335000 1.565000 0.395000 ;
        RECT 0.780000 1.055000 0.840000 1.335000 ;
        RECT 0.360000 1.055000 1.565000 1.115000 ;
        END
    END Y
END NAND3X2

MACRO AOI222X1
    CLASS CORE ;
    FOREIGN AOI222X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.260000 0.490000 0.340000 0.990000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.460000 0.220000 0.545000 0.715000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.880000 0.860000 1.095000 1.100000 ;
        RECT 0.860000 0.755000 0.940000 0.920000 ;
        RECT 0.880000 0.755000 0.940000 1.100000 ;
        RECT 0.860000 0.860000 1.095000 0.920000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.660000 0.620000 0.760000 0.920000 ;
        RECT 0.680000 0.620000 0.760000 1.100000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.195000 0.790000 1.340000 0.920000 ;
        RECT 1.195000 0.790000 1.275000 1.225000 ;
        END
    END C0
    PIN C1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.440000 0.620000 1.540000 1.100000 ;
        END
    END C1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 1.800000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 1.800000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.450000 0.410000 1.720000 0.520000 ;
        RECT 1.660000 0.980000 1.740000 1.260000 ;
        RECT 1.660000 0.410000 1.720000 1.260000 ;
        RECT 1.375000 1.200000 1.740000 1.260000 ;
        RECT 1.375000 1.200000 1.435000 1.320000 ;
        RECT 0.760000 0.460000 1.720000 0.520000 ;
        RECT 0.760000 0.380000 0.820000 0.520000 ;
        END
    END Y
END AOI222X1

MACRO NOR4X4
    CLASS CORE ;
    FOREIGN NOR4X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 3.800000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.860000 0.755000 0.940000 0.950000 ;
        RECT 0.350000 0.870000 0.940000 0.950000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.725000 0.755000 1.805000 0.895000 ;
        RECT 1.240000 0.815000 1.805000 0.895000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.435000 0.775000 2.570000 0.895000 ;
        RECT 2.110000 0.815000 2.570000 0.895000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 3.105000 0.775000 3.185000 0.895000 ;
        RECT 2.835000 0.815000 3.420000 0.895000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 3.800000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 3.800000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.060000 0.790000 1.140000 0.920000 ;
        RECT 3.460000 0.515000 3.520000 0.655000 ;
        RECT 3.405000 0.995000 3.465000 1.135000 ;
        RECT 3.050000 0.515000 3.110000 0.655000 ;
        RECT 2.995000 0.995000 3.055000 1.135000 ;
        RECT 2.640000 0.515000 2.700000 0.655000 ;
        RECT 2.230000 0.515000 2.290000 0.655000 ;
        RECT 1.820000 0.515000 1.880000 0.655000 ;
        RECT 1.410000 0.515000 1.470000 0.655000 ;
        RECT 1.080000 0.995000 3.465000 1.055000 ;
        RECT 1.080000 0.595000 1.140000 1.055000 ;
        RECT 1.000000 0.515000 1.060000 0.655000 ;
        RECT 0.590000 0.595000 3.520000 0.655000 ;
        RECT 0.590000 0.515000 0.650000 0.655000 ;
        END
    END Y
END NOR4X4

MACRO NOR4X2
    CLASS CORE ;
    FOREIGN NOR4X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.660000 0.980000 1.740000 1.185000 ;
        RECT 1.680000 0.820000 1.740000 1.185000 ;
        RECT 0.260000 1.125000 1.740000 1.185000 ;
        RECT 0.260000 0.820000 0.320000 1.185000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.460000 0.790000 0.540000 0.920000 ;
        RECT 1.435000 0.845000 1.495000 1.025000 ;
        RECT 0.480000 0.965000 1.495000 1.025000 ;
        RECT 0.480000 0.790000 0.540000 1.025000 ;
        RECT 0.420000 0.835000 0.540000 0.895000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.275000 0.625000 1.565000 0.705000 ;
        RECT 1.275000 0.625000 1.335000 0.865000 ;
        RECT 0.640000 0.805000 1.335000 0.865000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.640000 0.625000 1.140000 0.705000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 2.000000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 2.000000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.860000 1.170000 1.940000 1.345000 ;
        RECT 1.595000 0.445000 1.715000 0.525000 ;
        RECT 1.155000 0.445000 1.275000 0.525000 ;
        RECT 0.715000 0.445000 0.835000 0.525000 ;
        RECT 1.880000 0.465000 1.940000 1.345000 ;
        RECT 1.010000 1.285000 1.940000 1.345000 ;
        RECT 0.345000 0.465000 1.940000 0.525000 ;
        RECT 0.275000 0.445000 0.395000 0.505000 ;
        END
    END Y
END NOR4X2

MACRO NAND4X2
    CLASS CORE ;
    FOREIGN NAND4X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.200000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.860000 0.820000 1.940000 1.185000 ;
        RECT 0.260000 1.125000 1.940000 1.185000 ;
        RECT 0.260000 0.820000 0.320000 1.185000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.460000 0.790000 0.540000 0.920000 ;
        RECT 1.600000 0.845000 1.660000 1.025000 ;
        RECT 0.480000 0.965000 1.660000 1.025000 ;
        RECT 0.480000 0.790000 0.540000 1.025000 ;
        RECT 0.420000 0.835000 0.540000 0.895000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.235000 0.625000 1.395000 0.705000 ;
        RECT 1.335000 0.625000 1.395000 0.865000 ;
        RECT 0.685000 0.805000 1.395000 0.865000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.860000 0.625000 1.135000 0.705000 ;
        RECT 0.860000 0.400000 0.940000 0.705000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 2.200000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 2.200000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.060000 1.170000 2.140000 1.345000 ;
        RECT 2.060000 0.465000 2.120000 1.345000 ;
        RECT 1.730000 1.285000 1.790000 1.405000 ;
        RECT 1.260000 1.285000 1.320000 1.405000 ;
        RECT 1.185000 0.465000 2.120000 0.525000 ;
        RECT 1.070000 0.445000 1.235000 0.505000 ;
        RECT 0.790000 1.285000 0.850000 1.405000 ;
        RECT 0.320000 1.285000 2.140000 1.345000 ;
        RECT 0.320000 1.285000 0.380000 1.405000 ;
        END
    END Y
END NAND4X2

MACRO BUFX3
    CLASS CORE ;
    FOREIGN BUFX3 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.200000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.860000 0.720000 0.940000 1.220000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 1.200000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 1.200000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.260000 0.980000 0.340000 1.110000 ;
        RECT 0.625000 1.050000 0.685000 1.440000 ;
        RECT 0.585000 0.345000 0.645000 0.465000 ;
        RECT 0.540000 0.405000 0.645000 0.465000 ;
        RECT 0.540000 0.405000 0.600000 0.620000 ;
        RECT 0.260000 0.560000 0.320000 1.110000 ;
        RECT 0.215000 1.050000 0.685000 1.110000 ;
        RECT 0.215000 1.050000 0.275000 1.440000 ;
        RECT 0.175000 0.560000 0.600000 0.620000 ;
        RECT 0.175000 0.480000 0.235000 0.620000 ;
        END
    END Y
END BUFX3

MACRO AOI22X2
    CLASS CORE ;
    FOREIGN AOI22X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.200000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.840000 0.635000 1.065000 0.715000 ;
        RECT 0.840000 0.575000 0.920000 0.715000 ;
        RECT 0.480000 0.575000 0.920000 0.655000 ;
        RECT 0.480000 0.575000 0.560000 0.705000 ;
        RECT 0.235000 0.625000 0.560000 0.705000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.655000 0.715000 0.745000 0.960000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.840000 0.580000 1.960000 0.895000 ;
        RECT 1.840000 0.815000 2.165000 0.895000 ;
        RECT 1.500000 0.580000 1.960000 0.640000 ;
        RECT 1.500000 0.580000 1.560000 0.715000 ;
        RECT 1.325000 0.655000 1.560000 0.715000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.660000 0.740000 1.740000 1.030000 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 2.200000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 2.200000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.035000 0.815000 1.225000 0.895000 ;
        RECT 1.840000 0.995000 1.900000 1.165000 ;
        RECT 1.430000 1.105000 1.900000 1.165000 ;
        RECT 1.430000 0.835000 1.490000 1.165000 ;
        RECT 1.165000 0.415000 1.225000 0.895000 ;
        RECT 1.035000 0.835000 1.490000 0.895000 ;
        RECT 0.710000 0.415000 1.685000 0.475000 ;
        END
    END Y
END AOI22X2

MACRO OR4X1
    CLASS CORE ;
    FOREIGN OR4X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.060000 0.475000 1.140000 0.765000 ;
        RECT 0.850000 0.685000 1.140000 0.765000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.460000 0.980000 0.590000 1.070000 ;
        RECT 0.510000 0.660000 0.590000 1.070000 ;
        RECT 0.460000 0.980000 0.540000 1.110000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.330000 0.590000 0.410000 0.870000 ;
        RECT 0.260000 0.790000 0.410000 0.870000 ;
        RECT 0.260000 0.790000 0.340000 1.020000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.060000 0.590000 0.160000 0.795000 ;
        RECT 0.030000 0.735000 0.120000 1.040000 ;
        RECT 0.060000 0.590000 0.120000 1.040000 ;
        RECT 0.030000 0.735000 0.160000 0.795000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 1.400000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 1.400000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.240000 0.410000 1.340000 0.540000 ;
        RECT 1.240000 0.395000 1.300000 1.385000 ;
        END
    END Y
END OR4X1

MACRO NAND3X1
    CLASS CORE ;
    FOREIGN NAND3X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.000000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.260000 0.600000 0.340000 1.100000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.480000 0.480000 0.560000 0.890000 ;
        RECT 0.460000 0.410000 0.540000 0.540000 ;
        RECT 0.480000 0.410000 0.540000 0.890000 ;
        RECT 0.460000 0.480000 0.560000 0.540000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.660000 0.600000 0.740000 1.100000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 1.000000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 1.000000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.860000 1.200000 0.940000 1.490000 ;
        RECT 0.860000 0.440000 0.920000 1.490000 ;
        RECT 0.745000 0.440000 0.920000 0.500000 ;
        RECT 0.745000 0.380000 0.805000 0.500000 ;
        RECT 0.425000 1.200000 0.940000 1.260000 ;
        RECT 0.425000 1.200000 0.485000 1.480000 ;
        END
    END Y
END NAND3X1

MACRO NOR2X1
    CLASS CORE ;
    FOREIGN NOR2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.800000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.260000 0.570000 0.340000 1.070000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.460000 0.980000 0.560000 1.085000 ;
        RECT 0.480000 0.730000 0.560000 1.085000 ;
        RECT 0.460000 0.980000 0.540000 1.210000 ;
        RECT 0.480000 0.730000 0.540000 1.210000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 0.800000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 0.800000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.660000 0.600000 0.740000 0.730000 ;
        RECT 0.660000 0.570000 0.720000 1.290000 ;
        RECT 0.460000 0.570000 0.720000 0.630000 ;
        RECT 0.460000 0.490000 0.520000 0.630000 ;
        END
    END Y
END NOR2X1

MACRO AOI221X1
    CLASS CORE ;
    FOREIGN AOI221X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.260000 0.450000 0.340000 0.950000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.460000 0.220000 0.540000 0.720000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.060000 0.580000 1.140000 1.080000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.860000 0.580000 0.940000 1.080000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.260000 0.650000 1.380000 0.730000 ;
        RECT 1.260000 0.580000 1.340000 1.040000 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 1.800000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 1.800000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.460000 0.220000 1.540000 0.480000 ;
        RECT 1.480000 0.220000 1.540000 1.460000 ;
        RECT 0.870000 0.420000 1.540000 0.480000 ;
        RECT 0.800000 0.400000 0.920000 0.460000 ;
        END
    END Y
END AOI221X1

MACRO NAND4X1
    CLASS CORE ;
    FOREIGN NAND4X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.200000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.230000 0.650000 0.340000 0.920000 ;
        RECT 0.030000 0.840000 0.340000 0.920000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.480000 0.460000 0.560000 0.890000 ;
        RECT 0.460000 0.460000 0.560000 0.540000 ;
        RECT 0.460000 0.410000 0.540000 0.540000 ;
        RECT 0.480000 0.410000 0.540000 0.890000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.660000 0.220000 0.740000 0.830000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.860000 0.410000 0.940000 0.910000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 1.200000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 1.200000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.040000 0.790000 1.140000 1.080000 ;
        RECT 1.040000 0.540000 1.100000 1.080000 ;
        RECT 0.790000 1.020000 0.850000 1.300000 ;
        RECT 0.370000 1.020000 1.140000 1.080000 ;
        RECT 0.370000 1.020000 0.430000 1.300000 ;
        END
    END Y
END NAND4X1

MACRO AOI22X1
    CLASS CORE ;
    FOREIGN AOI22X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.260000 0.600000 0.340000 1.100000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.480000 0.270000 0.560000 0.700000 ;
        RECT 0.460000 0.270000 0.560000 0.350000 ;
        RECT 0.460000 0.220000 0.540000 0.350000 ;
        RECT 0.480000 0.220000 0.540000 0.700000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.060000 0.450000 1.140000 0.950000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.860000 0.410000 0.940000 0.910000 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 1.400000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 1.400000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.660000 0.980000 0.740000 1.110000 ;
        RECT 0.935000 1.050000 0.995000 1.190000 ;
        RECT 0.680000 0.370000 0.740000 1.110000 ;
        RECT 0.660000 1.050000 0.995000 1.110000 ;
        END
    END Y
END AOI22X1

MACRO BUFX6
    CLASS CORE ;
    FOREIGN BUFX6 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.460000 0.570000 1.540000 1.070000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 1.800000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 1.800000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.060000 0.790000 0.140000 0.975000 ;
        RECT 0.060000 0.350000 0.130000 1.370000 ;
        RECT 0.890000 0.915000 0.950000 1.370000 ;
        RECT 0.890000 0.350000 0.950000 0.655000 ;
        RECT 0.480000 0.915000 0.540000 1.370000 ;
        RECT 0.480000 0.350000 0.540000 0.655000 ;
        RECT 0.060000 0.915000 0.950000 0.975000 ;
        RECT 0.060000 0.595000 0.950000 0.655000 ;
        END
    END Y
END BUFX6

MACRO AO22XL
    CLASS CORE ;
    FOREIGN AO22XL 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.260000 0.600000 0.340000 1.100000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.460000 0.230000 0.540000 0.730000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.060000 0.790000 1.140000 1.230000 ;
        RECT 1.000000 0.790000 1.140000 0.870000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.660000 0.595000 0.740000 1.095000 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 1.600000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 1.600000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.260000 0.910000 1.510000 0.990000 ;
        RECT 1.260000 0.600000 1.340000 0.990000 ;
        RECT 1.250000 0.600000 1.340000 0.680000 ;
        RECT 1.250000 0.405000 1.330000 0.680000 ;
        RECT 1.260000 0.405000 1.330000 0.990000 ;
        END
    END Y
END AO22XL

MACRO MEM
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN MEM 0 0 ;
  SIZE 6.965 BY 6.80 ;
  SYMMETRY X Y R90 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 6.000 0.87 6.660 1.07 ;
      LAYER Metal6 ;
        RECT 6.000 0.87 6.660 1.07 ;
      LAYER Metal3 ;
        RECT 6.000 0.87 6.660 1.07 ;
      LAYER Metal4 ;
        RECT 6.000 0.87 6.660 1.07 ;
    END
  END A
  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 6.000 1.68 6.660 1.88 ;
      LAYER Metal6 ;
        RECT 6.000 1.68 6.660 1.88 ;
      LAYER Metal3 ;
        RECT 6.000 1.68 6.660 1.88 ;
      LAYER Metal4 ;
        RECT 6.000 1.68 6.660 1.88 ;
    END
  END CE
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal5 ;
        RECT 6.000 2.49 6.660 2.69 ;
      LAYER Metal6 ;
        RECT 6.000 2.49 6.660 2.69 ;
      LAYER Metal3 ;
        RECT 6.000 2.49 6.660 2.69 ;
      LAYER Metal4 ;
        RECT 6.000 2.49 6.660 2.69 ;
    END
  END CK
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 6.000 3.3 6.660 3.5 ;
      LAYER Metal6 ;
        RECT 6.000 3.3 6.660 3.5 ;
      LAYER Metal3 ;
        RECT 6.000 3.3 6.660 3.5 ;
      LAYER Metal4 ;
        RECT 6.000 3.3 6.660 3.5 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 6.000 4.11 6.660 4.31 ;
      LAYER Metal6 ;
        RECT 6.000 4.11 6.660 4.31 ;
      LAYER Metal3 ;
        RECT 6.000 4.11 6.660 4.31 ;
      LAYER Metal4 ;
        RECT 6.000 4.11 6.660 4.31 ;
    END
  END D[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 6.000 4.92 6.660 5.12 ;
      LAYER Metal6 ;
        RECT 6.000 4.92 6.660 5.12 ;
      LAYER Metal3 ;
        RECT 6.000 4.92 6.660 5.12 ;
      LAYER Metal4 ;
        RECT 6.000 4.92 6.660 5.12 ;
    END
  END Q[0]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 6.000 5.73 6.660 5.93 ;
      LAYER Metal6 ;
        RECT 6.000 5.73 6.660 5.93 ;
      LAYER Metal3 ;
        RECT 6.000 5.73 6.660 5.93 ;
      LAYER Metal4 ;
        RECT 6.000 5.73 6.660 5.93 ;
    END
  END Q[1]
  OBS
    LAYER Metal1 ;
      RECT 1 1 6 6 ;
    LAYER Metal2 ;
      RECT 1 1 6 6 ;
    LAYER Metal3 ;
      RECT 1 1 6 6 ;
    LAYER Metal4 ;
      RECT 1 1 6 6 ;
    LAYER Metal5 ;
      RECT 1 1 6 6 ;
    LAYER Metal6 ;
      RECT 1 1 6 6 ;
  END
END MEM

END LIBRARY
