module div( input [3:0] a, output [3:0] b);
assign b = a / 4'b0011;
endmodule

