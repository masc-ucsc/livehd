module trivial_assign( input a, output c);
assign c = a;
endmodule

