module tuple_nested2(
   output reg signed [5:0] out
);
always @(*) begin
  out = 3;
end
endmodule
