module scalar_tuple (
  output [2:0] out1,
  output [3:0] out2,
  output [3:0] out3,
  output [3:0] out4,
  output [2:0] out5,
  output [2:0] out6,
  output [1:0] out7,
  output [1:0] out8,
  /* output [2:0] out9, */
  output [2:0] out10
);

assign out1  = 3'd7;
assign out2  = 4'd8;
assign out3  = 4'd9;
assign out4  = 4'd10;
assign out5  = 3'd7;
assign out6  = 3'd6;
assign out7  = 2'd3;
assign out8  = 2'd3;
/* assign out9  = 3'd7; */
assign out10 = 3'd5;

endmodule
