module tuple_copy (
  output [2:0] out
);

assign out = 3'd5;

endmodule
