module xor_100000(
    input a,
    input b,
    output wire z
    );

    wire t0 = a ^ b;
    wire t1 = t0 ^ t0;
    wire t2 = t1 ^ t1;
    wire t3 = t2 ^ t2;
    wire t4 = t3 ^ t3;
    wire t5 = t4 ^ t4;
    wire t6 = t5 ^ t5;
    wire t7 = t6 ^ t6;
    wire t8 = t7 ^ t7;
    wire t9 = t8 ^ t8;
    wire t10 = t9 ^ t9;
    wire t11 = t10 ^ t10;
    wire t12 = t11 ^ t11;
    wire t13 = t12 ^ t12;
    wire t14 = t13 ^ t13;
    wire t15 = t14 ^ t14;
    wire t16 = t15 ^ t15;
    wire t17 = t16 ^ t16;
    wire t18 = t17 ^ t17;
    wire t19 = t18 ^ t18;
    wire t20 = t19 ^ t19;
    wire t21 = t20 ^ t20;
    wire t22 = t21 ^ t21;
    wire t23 = t22 ^ t22;
    wire t24 = t23 ^ t23;
    wire t25 = t24 ^ t24;
    wire t26 = t25 ^ t25;
    wire t27 = t26 ^ t26;
    wire t28 = t27 ^ t27;
    wire t29 = t28 ^ t28;
    wire t30 = t29 ^ t29;
    wire t31 = t30 ^ t30;
    wire t32 = t31 ^ t31;
    wire t33 = t32 ^ t32;
    wire t34 = t33 ^ t33;
    wire t35 = t34 ^ t34;
    wire t36 = t35 ^ t35;
    wire t37 = t36 ^ t36;
    wire t38 = t37 ^ t37;
    wire t39 = t38 ^ t38;
    wire t40 = t39 ^ t39;
    wire t41 = t40 ^ t40;
    wire t42 = t41 ^ t41;
    wire t43 = t42 ^ t42;
    wire t44 = t43 ^ t43;
    wire t45 = t44 ^ t44;
    wire t46 = t45 ^ t45;
    wire t47 = t46 ^ t46;
    wire t48 = t47 ^ t47;
    wire t49 = t48 ^ t48;
    wire t50 = t49 ^ t49;
    wire t51 = t50 ^ t50;
    wire t52 = t51 ^ t51;
    wire t53 = t52 ^ t52;
    wire t54 = t53 ^ t53;
    wire t55 = t54 ^ t54;
    wire t56 = t55 ^ t55;
    wire t57 = t56 ^ t56;
    wire t58 = t57 ^ t57;
    wire t59 = t58 ^ t58;
    wire t60 = t59 ^ t59;
    wire t61 = t60 ^ t60;
    wire t62 = t61 ^ t61;
    wire t63 = t62 ^ t62;
    wire t64 = t63 ^ t63;
    wire t65 = t64 ^ t64;
    wire t66 = t65 ^ t65;
    wire t67 = t66 ^ t66;
    wire t68 = t67 ^ t67;
    wire t69 = t68 ^ t68;
    wire t70 = t69 ^ t69;
    wire t71 = t70 ^ t70;
    wire t72 = t71 ^ t71;
    wire t73 = t72 ^ t72;
    wire t74 = t73 ^ t73;
    wire t75 = t74 ^ t74;
    wire t76 = t75 ^ t75;
    wire t77 = t76 ^ t76;
    wire t78 = t77 ^ t77;
    wire t79 = t78 ^ t78;
    wire t80 = t79 ^ t79;
    wire t81 = t80 ^ t80;
    wire t82 = t81 ^ t81;
    wire t83 = t82 ^ t82;
    wire t84 = t83 ^ t83;
    wire t85 = t84 ^ t84;
    wire t86 = t85 ^ t85;
    wire t87 = t86 ^ t86;
    wire t88 = t87 ^ t87;
    wire t89 = t88 ^ t88;
    wire t90 = t89 ^ t89;
    wire t91 = t90 ^ t90;
    wire t92 = t91 ^ t91;
    wire t93 = t92 ^ t92;
    wire t94 = t93 ^ t93;
    wire t95 = t94 ^ t94;
    wire t96 = t95 ^ t95;
    wire t97 = t96 ^ t96;
    wire t98 = t97 ^ t97;
    wire t99 = t98 ^ t98;
    wire t100 = t99 ^ t99;
    wire t101 = t100 ^ t100;
    wire t102 = t101 ^ t101;
    wire t103 = t102 ^ t102;
    wire t104 = t103 ^ t103;
    wire t105 = t104 ^ t104;
    wire t106 = t105 ^ t105;
    wire t107 = t106 ^ t106;
    wire t108 = t107 ^ t107;
    wire t109 = t108 ^ t108;
    wire t110 = t109 ^ t109;
    wire t111 = t110 ^ t110;
    wire t112 = t111 ^ t111;
    wire t113 = t112 ^ t112;
    wire t114 = t113 ^ t113;
    wire t115 = t114 ^ t114;
    wire t116 = t115 ^ t115;
    wire t117 = t116 ^ t116;
    wire t118 = t117 ^ t117;
    wire t119 = t118 ^ t118;
    wire t120 = t119 ^ t119;
    wire t121 = t120 ^ t120;
    wire t122 = t121 ^ t121;
    wire t123 = t122 ^ t122;
    wire t124 = t123 ^ t123;
    wire t125 = t124 ^ t124;
    wire t126 = t125 ^ t125;
    wire t127 = t126 ^ t126;
    wire t128 = t127 ^ t127;
    wire t129 = t128 ^ t128;
    wire t130 = t129 ^ t129;
    wire t131 = t130 ^ t130;
    wire t132 = t131 ^ t131;
    wire t133 = t132 ^ t132;
    wire t134 = t133 ^ t133;
    wire t135 = t134 ^ t134;
    wire t136 = t135 ^ t135;
    wire t137 = t136 ^ t136;
    wire t138 = t137 ^ t137;
    wire t139 = t138 ^ t138;
    wire t140 = t139 ^ t139;
    wire t141 = t140 ^ t140;
    wire t142 = t141 ^ t141;
    wire t143 = t142 ^ t142;
    wire t144 = t143 ^ t143;
    wire t145 = t144 ^ t144;
    wire t146 = t145 ^ t145;
    wire t147 = t146 ^ t146;
    wire t148 = t147 ^ t147;
    wire t149 = t148 ^ t148;
    wire t150 = t149 ^ t149;
    wire t151 = t150 ^ t150;
    wire t152 = t151 ^ t151;
    wire t153 = t152 ^ t152;
    wire t154 = t153 ^ t153;
    wire t155 = t154 ^ t154;
    wire t156 = t155 ^ t155;
    wire t157 = t156 ^ t156;
    wire t158 = t157 ^ t157;
    wire t159 = t158 ^ t158;
    wire t160 = t159 ^ t159;
    wire t161 = t160 ^ t160;
    wire t162 = t161 ^ t161;
    wire t163 = t162 ^ t162;
    wire t164 = t163 ^ t163;
    wire t165 = t164 ^ t164;
    wire t166 = t165 ^ t165;
    wire t167 = t166 ^ t166;
    wire t168 = t167 ^ t167;
    wire t169 = t168 ^ t168;
    wire t170 = t169 ^ t169;
    wire t171 = t170 ^ t170;
    wire t172 = t171 ^ t171;
    wire t173 = t172 ^ t172;
    wire t174 = t173 ^ t173;
    wire t175 = t174 ^ t174;
    wire t176 = t175 ^ t175;
    wire t177 = t176 ^ t176;
    wire t178 = t177 ^ t177;
    wire t179 = t178 ^ t178;
    wire t180 = t179 ^ t179;
    wire t181 = t180 ^ t180;
    wire t182 = t181 ^ t181;
    wire t183 = t182 ^ t182;
    wire t184 = t183 ^ t183;
    wire t185 = t184 ^ t184;
    wire t186 = t185 ^ t185;
    wire t187 = t186 ^ t186;
    wire t188 = t187 ^ t187;
    wire t189 = t188 ^ t188;
    wire t190 = t189 ^ t189;
    wire t191 = t190 ^ t190;
    wire t192 = t191 ^ t191;
    wire t193 = t192 ^ t192;
    wire t194 = t193 ^ t193;
    wire t195 = t194 ^ t194;
    wire t196 = t195 ^ t195;
    wire t197 = t196 ^ t196;
    wire t198 = t197 ^ t197;
    wire t199 = t198 ^ t198;
    wire t200 = t199 ^ t199;
    wire t201 = t200 ^ t200;
    wire t202 = t201 ^ t201;
    wire t203 = t202 ^ t202;
    wire t204 = t203 ^ t203;
    wire t205 = t204 ^ t204;
    wire t206 = t205 ^ t205;
    wire t207 = t206 ^ t206;
    wire t208 = t207 ^ t207;
    wire t209 = t208 ^ t208;
    wire t210 = t209 ^ t209;
    wire t211 = t210 ^ t210;
    wire t212 = t211 ^ t211;
    wire t213 = t212 ^ t212;
    wire t214 = t213 ^ t213;
    wire t215 = t214 ^ t214;
    wire t216 = t215 ^ t215;
    wire t217 = t216 ^ t216;
    wire t218 = t217 ^ t217;
    wire t219 = t218 ^ t218;
    wire t220 = t219 ^ t219;
    wire t221 = t220 ^ t220;
    wire t222 = t221 ^ t221;
    wire t223 = t222 ^ t222;
    wire t224 = t223 ^ t223;
    wire t225 = t224 ^ t224;
    wire t226 = t225 ^ t225;
    wire t227 = t226 ^ t226;
    wire t228 = t227 ^ t227;
    wire t229 = t228 ^ t228;
    wire t230 = t229 ^ t229;
    wire t231 = t230 ^ t230;
    wire t232 = t231 ^ t231;
    wire t233 = t232 ^ t232;
    wire t234 = t233 ^ t233;
    wire t235 = t234 ^ t234;
    wire t236 = t235 ^ t235;
    wire t237 = t236 ^ t236;
    wire t238 = t237 ^ t237;
    wire t239 = t238 ^ t238;
    wire t240 = t239 ^ t239;
    wire t241 = t240 ^ t240;
    wire t242 = t241 ^ t241;
    wire t243 = t242 ^ t242;
    wire t244 = t243 ^ t243;
    wire t245 = t244 ^ t244;
    wire t246 = t245 ^ t245;
    wire t247 = t246 ^ t246;
    wire t248 = t247 ^ t247;
    wire t249 = t248 ^ t248;
    wire t250 = t249 ^ t249;
    wire t251 = t250 ^ t250;
    wire t252 = t251 ^ t251;
    wire t253 = t252 ^ t252;
    wire t254 = t253 ^ t253;
    wire t255 = t254 ^ t254;
    wire t256 = t255 ^ t255;
    wire t257 = t256 ^ t256;
    wire t258 = t257 ^ t257;
    wire t259 = t258 ^ t258;
    wire t260 = t259 ^ t259;
    wire t261 = t260 ^ t260;
    wire t262 = t261 ^ t261;
    wire t263 = t262 ^ t262;
    wire t264 = t263 ^ t263;
    wire t265 = t264 ^ t264;
    wire t266 = t265 ^ t265;
    wire t267 = t266 ^ t266;
    wire t268 = t267 ^ t267;
    wire t269 = t268 ^ t268;
    wire t270 = t269 ^ t269;
    wire t271 = t270 ^ t270;
    wire t272 = t271 ^ t271;
    wire t273 = t272 ^ t272;
    wire t274 = t273 ^ t273;
    wire t275 = t274 ^ t274;
    wire t276 = t275 ^ t275;
    wire t277 = t276 ^ t276;
    wire t278 = t277 ^ t277;
    wire t279 = t278 ^ t278;
    wire t280 = t279 ^ t279;
    wire t281 = t280 ^ t280;
    wire t282 = t281 ^ t281;
    wire t283 = t282 ^ t282;
    wire t284 = t283 ^ t283;
    wire t285 = t284 ^ t284;
    wire t286 = t285 ^ t285;
    wire t287 = t286 ^ t286;
    wire t288 = t287 ^ t287;
    wire t289 = t288 ^ t288;
    wire t290 = t289 ^ t289;
    wire t291 = t290 ^ t290;
    wire t292 = t291 ^ t291;
    wire t293 = t292 ^ t292;
    wire t294 = t293 ^ t293;
    wire t295 = t294 ^ t294;
    wire t296 = t295 ^ t295;
    wire t297 = t296 ^ t296;
    wire t298 = t297 ^ t297;
    wire t299 = t298 ^ t298;
    wire t300 = t299 ^ t299;
    wire t301 = t300 ^ t300;
    wire t302 = t301 ^ t301;
    wire t303 = t302 ^ t302;
    wire t304 = t303 ^ t303;
    wire t305 = t304 ^ t304;
    wire t306 = t305 ^ t305;
    wire t307 = t306 ^ t306;
    wire t308 = t307 ^ t307;
    wire t309 = t308 ^ t308;
    wire t310 = t309 ^ t309;
    wire t311 = t310 ^ t310;
    wire t312 = t311 ^ t311;
    wire t313 = t312 ^ t312;
    wire t314 = t313 ^ t313;
    wire t315 = t314 ^ t314;
    wire t316 = t315 ^ t315;
    wire t317 = t316 ^ t316;
    wire t318 = t317 ^ t317;
    wire t319 = t318 ^ t318;
    wire t320 = t319 ^ t319;
    wire t321 = t320 ^ t320;
    wire t322 = t321 ^ t321;
    wire t323 = t322 ^ t322;
    wire t324 = t323 ^ t323;
    wire t325 = t324 ^ t324;
    wire t326 = t325 ^ t325;
    wire t327 = t326 ^ t326;
    wire t328 = t327 ^ t327;
    wire t329 = t328 ^ t328;
    wire t330 = t329 ^ t329;
    wire t331 = t330 ^ t330;
    wire t332 = t331 ^ t331;
    wire t333 = t332 ^ t332;
    wire t334 = t333 ^ t333;
    wire t335 = t334 ^ t334;
    wire t336 = t335 ^ t335;
    wire t337 = t336 ^ t336;
    wire t338 = t337 ^ t337;
    wire t339 = t338 ^ t338;
    wire t340 = t339 ^ t339;
    wire t341 = t340 ^ t340;
    wire t342 = t341 ^ t341;
    wire t343 = t342 ^ t342;
    wire t344 = t343 ^ t343;
    wire t345 = t344 ^ t344;
    wire t346 = t345 ^ t345;
    wire t347 = t346 ^ t346;
    wire t348 = t347 ^ t347;
    wire t349 = t348 ^ t348;
    wire t350 = t349 ^ t349;
    wire t351 = t350 ^ t350;
    wire t352 = t351 ^ t351;
    wire t353 = t352 ^ t352;
    wire t354 = t353 ^ t353;
    wire t355 = t354 ^ t354;
    wire t356 = t355 ^ t355;
    wire t357 = t356 ^ t356;
    wire t358 = t357 ^ t357;
    wire t359 = t358 ^ t358;
    wire t360 = t359 ^ t359;
    wire t361 = t360 ^ t360;
    wire t362 = t361 ^ t361;
    wire t363 = t362 ^ t362;
    wire t364 = t363 ^ t363;
    wire t365 = t364 ^ t364;
    wire t366 = t365 ^ t365;
    wire t367 = t366 ^ t366;
    wire t368 = t367 ^ t367;
    wire t369 = t368 ^ t368;
    wire t370 = t369 ^ t369;
    wire t371 = t370 ^ t370;
    wire t372 = t371 ^ t371;
    wire t373 = t372 ^ t372;
    wire t374 = t373 ^ t373;
    wire t375 = t374 ^ t374;
    wire t376 = t375 ^ t375;
    wire t377 = t376 ^ t376;
    wire t378 = t377 ^ t377;
    wire t379 = t378 ^ t378;
    wire t380 = t379 ^ t379;
    wire t381 = t380 ^ t380;
    wire t382 = t381 ^ t381;
    wire t383 = t382 ^ t382;
    wire t384 = t383 ^ t383;
    wire t385 = t384 ^ t384;
    wire t386 = t385 ^ t385;
    wire t387 = t386 ^ t386;
    wire t388 = t387 ^ t387;
    wire t389 = t388 ^ t388;
    wire t390 = t389 ^ t389;
    wire t391 = t390 ^ t390;
    wire t392 = t391 ^ t391;
    wire t393 = t392 ^ t392;
    wire t394 = t393 ^ t393;
    wire t395 = t394 ^ t394;
    wire t396 = t395 ^ t395;
    wire t397 = t396 ^ t396;
    wire t398 = t397 ^ t397;
    wire t399 = t398 ^ t398;
    wire t400 = t399 ^ t399;
    wire t401 = t400 ^ t400;
    wire t402 = t401 ^ t401;
    wire t403 = t402 ^ t402;
    wire t404 = t403 ^ t403;
    wire t405 = t404 ^ t404;
    wire t406 = t405 ^ t405;
    wire t407 = t406 ^ t406;
    wire t408 = t407 ^ t407;
    wire t409 = t408 ^ t408;
    wire t410 = t409 ^ t409;
    wire t411 = t410 ^ t410;
    wire t412 = t411 ^ t411;
    wire t413 = t412 ^ t412;
    wire t414 = t413 ^ t413;
    wire t415 = t414 ^ t414;
    wire t416 = t415 ^ t415;
    wire t417 = t416 ^ t416;
    wire t418 = t417 ^ t417;
    wire t419 = t418 ^ t418;
    wire t420 = t419 ^ t419;
    wire t421 = t420 ^ t420;
    wire t422 = t421 ^ t421;
    wire t423 = t422 ^ t422;
    wire t424 = t423 ^ t423;
    wire t425 = t424 ^ t424;
    wire t426 = t425 ^ t425;
    wire t427 = t426 ^ t426;
    wire t428 = t427 ^ t427;
    wire t429 = t428 ^ t428;
    wire t430 = t429 ^ t429;
    wire t431 = t430 ^ t430;
    wire t432 = t431 ^ t431;
    wire t433 = t432 ^ t432;
    wire t434 = t433 ^ t433;
    wire t435 = t434 ^ t434;
    wire t436 = t435 ^ t435;
    wire t437 = t436 ^ t436;
    wire t438 = t437 ^ t437;
    wire t439 = t438 ^ t438;
    wire t440 = t439 ^ t439;
    wire t441 = t440 ^ t440;
    wire t442 = t441 ^ t441;
    wire t443 = t442 ^ t442;
    wire t444 = t443 ^ t443;
    wire t445 = t444 ^ t444;
    wire t446 = t445 ^ t445;
    wire t447 = t446 ^ t446;
    wire t448 = t447 ^ t447;
    wire t449 = t448 ^ t448;
    wire t450 = t449 ^ t449;
    wire t451 = t450 ^ t450;
    wire t452 = t451 ^ t451;
    wire t453 = t452 ^ t452;
    wire t454 = t453 ^ t453;
    wire t455 = t454 ^ t454;
    wire t456 = t455 ^ t455;
    wire t457 = t456 ^ t456;
    wire t458 = t457 ^ t457;
    wire t459 = t458 ^ t458;
    wire t460 = t459 ^ t459;
    wire t461 = t460 ^ t460;
    wire t462 = t461 ^ t461;
    wire t463 = t462 ^ t462;
    wire t464 = t463 ^ t463;
    wire t465 = t464 ^ t464;
    wire t466 = t465 ^ t465;
    wire t467 = t466 ^ t466;
    wire t468 = t467 ^ t467;
    wire t469 = t468 ^ t468;
    wire t470 = t469 ^ t469;
    wire t471 = t470 ^ t470;
    wire t472 = t471 ^ t471;
    wire t473 = t472 ^ t472;
    wire t474 = t473 ^ t473;
    wire t475 = t474 ^ t474;
    wire t476 = t475 ^ t475;
    wire t477 = t476 ^ t476;
    wire t478 = t477 ^ t477;
    wire t479 = t478 ^ t478;
    wire t480 = t479 ^ t479;
    wire t481 = t480 ^ t480;
    wire t482 = t481 ^ t481;
    wire t483 = t482 ^ t482;
    wire t484 = t483 ^ t483;
    wire t485 = t484 ^ t484;
    wire t486 = t485 ^ t485;
    wire t487 = t486 ^ t486;
    wire t488 = t487 ^ t487;
    wire t489 = t488 ^ t488;
    wire t490 = t489 ^ t489;
    wire t491 = t490 ^ t490;
    wire t492 = t491 ^ t491;
    wire t493 = t492 ^ t492;
    wire t494 = t493 ^ t493;
    wire t495 = t494 ^ t494;
    wire t496 = t495 ^ t495;
    wire t497 = t496 ^ t496;
    wire t498 = t497 ^ t497;
    wire t499 = t498 ^ t498;
    wire t500 = t499 ^ t499;
    wire t501 = t500 ^ t500;
    wire t502 = t501 ^ t501;
    wire t503 = t502 ^ t502;
    wire t504 = t503 ^ t503;
    wire t505 = t504 ^ t504;
    wire t506 = t505 ^ t505;
    wire t507 = t506 ^ t506;
    wire t508 = t507 ^ t507;
    wire t509 = t508 ^ t508;
    wire t510 = t509 ^ t509;
    wire t511 = t510 ^ t510;
    wire t512 = t511 ^ t511;
    wire t513 = t512 ^ t512;
    wire t514 = t513 ^ t513;
    wire t515 = t514 ^ t514;
    wire t516 = t515 ^ t515;
    wire t517 = t516 ^ t516;
    wire t518 = t517 ^ t517;
    wire t519 = t518 ^ t518;
    wire t520 = t519 ^ t519;
    wire t521 = t520 ^ t520;
    wire t522 = t521 ^ t521;
    wire t523 = t522 ^ t522;
    wire t524 = t523 ^ t523;
    wire t525 = t524 ^ t524;
    wire t526 = t525 ^ t525;
    wire t527 = t526 ^ t526;
    wire t528 = t527 ^ t527;
    wire t529 = t528 ^ t528;
    wire t530 = t529 ^ t529;
    wire t531 = t530 ^ t530;
    wire t532 = t531 ^ t531;
    wire t533 = t532 ^ t532;
    wire t534 = t533 ^ t533;
    wire t535 = t534 ^ t534;
    wire t536 = t535 ^ t535;
    wire t537 = t536 ^ t536;
    wire t538 = t537 ^ t537;
    wire t539 = t538 ^ t538;
    wire t540 = t539 ^ t539;
    wire t541 = t540 ^ t540;
    wire t542 = t541 ^ t541;
    wire t543 = t542 ^ t542;
    wire t544 = t543 ^ t543;
    wire t545 = t544 ^ t544;
    wire t546 = t545 ^ t545;
    wire t547 = t546 ^ t546;
    wire t548 = t547 ^ t547;
    wire t549 = t548 ^ t548;
    wire t550 = t549 ^ t549;
    wire t551 = t550 ^ t550;
    wire t552 = t551 ^ t551;
    wire t553 = t552 ^ t552;
    wire t554 = t553 ^ t553;
    wire t555 = t554 ^ t554;
    wire t556 = t555 ^ t555;
    wire t557 = t556 ^ t556;
    wire t558 = t557 ^ t557;
    wire t559 = t558 ^ t558;
    wire t560 = t559 ^ t559;
    wire t561 = t560 ^ t560;
    wire t562 = t561 ^ t561;
    wire t563 = t562 ^ t562;
    wire t564 = t563 ^ t563;
    wire t565 = t564 ^ t564;
    wire t566 = t565 ^ t565;
    wire t567 = t566 ^ t566;
    wire t568 = t567 ^ t567;
    wire t569 = t568 ^ t568;
    wire t570 = t569 ^ t569;
    wire t571 = t570 ^ t570;
    wire t572 = t571 ^ t571;
    wire t573 = t572 ^ t572;
    wire t574 = t573 ^ t573;
    wire t575 = t574 ^ t574;
    wire t576 = t575 ^ t575;
    wire t577 = t576 ^ t576;
    wire t578 = t577 ^ t577;
    wire t579 = t578 ^ t578;
    wire t580 = t579 ^ t579;
    wire t581 = t580 ^ t580;
    wire t582 = t581 ^ t581;
    wire t583 = t582 ^ t582;
    wire t584 = t583 ^ t583;
    wire t585 = t584 ^ t584;
    wire t586 = t585 ^ t585;
    wire t587 = t586 ^ t586;
    wire t588 = t587 ^ t587;
    wire t589 = t588 ^ t588;
    wire t590 = t589 ^ t589;
    wire t591 = t590 ^ t590;
    wire t592 = t591 ^ t591;
    wire t593 = t592 ^ t592;
    wire t594 = t593 ^ t593;
    wire t595 = t594 ^ t594;
    wire t596 = t595 ^ t595;
    wire t597 = t596 ^ t596;
    wire t598 = t597 ^ t597;
    wire t599 = t598 ^ t598;
    wire t600 = t599 ^ t599;
    wire t601 = t600 ^ t600;
    wire t602 = t601 ^ t601;
    wire t603 = t602 ^ t602;
    wire t604 = t603 ^ t603;
    wire t605 = t604 ^ t604;
    wire t606 = t605 ^ t605;
    wire t607 = t606 ^ t606;
    wire t608 = t607 ^ t607;
    wire t609 = t608 ^ t608;
    wire t610 = t609 ^ t609;
    wire t611 = t610 ^ t610;
    wire t612 = t611 ^ t611;
    wire t613 = t612 ^ t612;
    wire t614 = t613 ^ t613;
    wire t615 = t614 ^ t614;
    wire t616 = t615 ^ t615;
    wire t617 = t616 ^ t616;
    wire t618 = t617 ^ t617;
    wire t619 = t618 ^ t618;
    wire t620 = t619 ^ t619;
    wire t621 = t620 ^ t620;
    wire t622 = t621 ^ t621;
    wire t623 = t622 ^ t622;
    wire t624 = t623 ^ t623;
    wire t625 = t624 ^ t624;
    wire t626 = t625 ^ t625;
    wire t627 = t626 ^ t626;
    wire t628 = t627 ^ t627;
    wire t629 = t628 ^ t628;
    wire t630 = t629 ^ t629;
    wire t631 = t630 ^ t630;
    wire t632 = t631 ^ t631;
    wire t633 = t632 ^ t632;
    wire t634 = t633 ^ t633;
    wire t635 = t634 ^ t634;
    wire t636 = t635 ^ t635;
    wire t637 = t636 ^ t636;
    wire t638 = t637 ^ t637;
    wire t639 = t638 ^ t638;
    wire t640 = t639 ^ t639;
    wire t641 = t640 ^ t640;
    wire t642 = t641 ^ t641;
    wire t643 = t642 ^ t642;
    wire t644 = t643 ^ t643;
    wire t645 = t644 ^ t644;
    wire t646 = t645 ^ t645;
    wire t647 = t646 ^ t646;
    wire t648 = t647 ^ t647;
    wire t649 = t648 ^ t648;
    wire t650 = t649 ^ t649;
    wire t651 = t650 ^ t650;
    wire t652 = t651 ^ t651;
    wire t653 = t652 ^ t652;
    wire t654 = t653 ^ t653;
    wire t655 = t654 ^ t654;
    wire t656 = t655 ^ t655;
    wire t657 = t656 ^ t656;
    wire t658 = t657 ^ t657;
    wire t659 = t658 ^ t658;
    wire t660 = t659 ^ t659;
    wire t661 = t660 ^ t660;
    wire t662 = t661 ^ t661;
    wire t663 = t662 ^ t662;
    wire t664 = t663 ^ t663;
    wire t665 = t664 ^ t664;
    wire t666 = t665 ^ t665;
    wire t667 = t666 ^ t666;
    wire t668 = t667 ^ t667;
    wire t669 = t668 ^ t668;
    wire t670 = t669 ^ t669;
    wire t671 = t670 ^ t670;
    wire t672 = t671 ^ t671;
    wire t673 = t672 ^ t672;
    wire t674 = t673 ^ t673;
    wire t675 = t674 ^ t674;
    wire t676 = t675 ^ t675;
    wire t677 = t676 ^ t676;
    wire t678 = t677 ^ t677;
    wire t679 = t678 ^ t678;
    wire t680 = t679 ^ t679;
    wire t681 = t680 ^ t680;
    wire t682 = t681 ^ t681;
    wire t683 = t682 ^ t682;
    wire t684 = t683 ^ t683;
    wire t685 = t684 ^ t684;
    wire t686 = t685 ^ t685;
    wire t687 = t686 ^ t686;
    wire t688 = t687 ^ t687;
    wire t689 = t688 ^ t688;
    wire t690 = t689 ^ t689;
    wire t691 = t690 ^ t690;
    wire t692 = t691 ^ t691;
    wire t693 = t692 ^ t692;
    wire t694 = t693 ^ t693;
    wire t695 = t694 ^ t694;
    wire t696 = t695 ^ t695;
    wire t697 = t696 ^ t696;
    wire t698 = t697 ^ t697;
    wire t699 = t698 ^ t698;
    wire t700 = t699 ^ t699;
    wire t701 = t700 ^ t700;
    wire t702 = t701 ^ t701;
    wire t703 = t702 ^ t702;
    wire t704 = t703 ^ t703;
    wire t705 = t704 ^ t704;
    wire t706 = t705 ^ t705;
    wire t707 = t706 ^ t706;
    wire t708 = t707 ^ t707;
    wire t709 = t708 ^ t708;
    wire t710 = t709 ^ t709;
    wire t711 = t710 ^ t710;
    wire t712 = t711 ^ t711;
    wire t713 = t712 ^ t712;
    wire t714 = t713 ^ t713;
    wire t715 = t714 ^ t714;
    wire t716 = t715 ^ t715;
    wire t717 = t716 ^ t716;
    wire t718 = t717 ^ t717;
    wire t719 = t718 ^ t718;
    wire t720 = t719 ^ t719;
    wire t721 = t720 ^ t720;
    wire t722 = t721 ^ t721;
    wire t723 = t722 ^ t722;
    wire t724 = t723 ^ t723;
    wire t725 = t724 ^ t724;
    wire t726 = t725 ^ t725;
    wire t727 = t726 ^ t726;
    wire t728 = t727 ^ t727;
    wire t729 = t728 ^ t728;
    wire t730 = t729 ^ t729;
    wire t731 = t730 ^ t730;
    wire t732 = t731 ^ t731;
    wire t733 = t732 ^ t732;
    wire t734 = t733 ^ t733;
    wire t735 = t734 ^ t734;
    wire t736 = t735 ^ t735;
    wire t737 = t736 ^ t736;
    wire t738 = t737 ^ t737;
    wire t739 = t738 ^ t738;
    wire t740 = t739 ^ t739;
    wire t741 = t740 ^ t740;
    wire t742 = t741 ^ t741;
    wire t743 = t742 ^ t742;
    wire t744 = t743 ^ t743;
    wire t745 = t744 ^ t744;
    wire t746 = t745 ^ t745;
    wire t747 = t746 ^ t746;
    wire t748 = t747 ^ t747;
    wire t749 = t748 ^ t748;
    wire t750 = t749 ^ t749;
    wire t751 = t750 ^ t750;
    wire t752 = t751 ^ t751;
    wire t753 = t752 ^ t752;
    wire t754 = t753 ^ t753;
    wire t755 = t754 ^ t754;
    wire t756 = t755 ^ t755;
    wire t757 = t756 ^ t756;
    wire t758 = t757 ^ t757;
    wire t759 = t758 ^ t758;
    wire t760 = t759 ^ t759;
    wire t761 = t760 ^ t760;
    wire t762 = t761 ^ t761;
    wire t763 = t762 ^ t762;
    wire t764 = t763 ^ t763;
    wire t765 = t764 ^ t764;
    wire t766 = t765 ^ t765;
    wire t767 = t766 ^ t766;
    wire t768 = t767 ^ t767;
    wire t769 = t768 ^ t768;
    wire t770 = t769 ^ t769;
    wire t771 = t770 ^ t770;
    wire t772 = t771 ^ t771;
    wire t773 = t772 ^ t772;
    wire t774 = t773 ^ t773;
    wire t775 = t774 ^ t774;
    wire t776 = t775 ^ t775;
    wire t777 = t776 ^ t776;
    wire t778 = t777 ^ t777;
    wire t779 = t778 ^ t778;
    wire t780 = t779 ^ t779;
    wire t781 = t780 ^ t780;
    wire t782 = t781 ^ t781;
    wire t783 = t782 ^ t782;
    wire t784 = t783 ^ t783;
    wire t785 = t784 ^ t784;
    wire t786 = t785 ^ t785;
    wire t787 = t786 ^ t786;
    wire t788 = t787 ^ t787;
    wire t789 = t788 ^ t788;
    wire t790 = t789 ^ t789;
    wire t791 = t790 ^ t790;
    wire t792 = t791 ^ t791;
    wire t793 = t792 ^ t792;
    wire t794 = t793 ^ t793;
    wire t795 = t794 ^ t794;
    wire t796 = t795 ^ t795;
    wire t797 = t796 ^ t796;
    wire t798 = t797 ^ t797;
    wire t799 = t798 ^ t798;
    wire t800 = t799 ^ t799;
    wire t801 = t800 ^ t800;
    wire t802 = t801 ^ t801;
    wire t803 = t802 ^ t802;
    wire t804 = t803 ^ t803;
    wire t805 = t804 ^ t804;
    wire t806 = t805 ^ t805;
    wire t807 = t806 ^ t806;
    wire t808 = t807 ^ t807;
    wire t809 = t808 ^ t808;
    wire t810 = t809 ^ t809;
    wire t811 = t810 ^ t810;
    wire t812 = t811 ^ t811;
    wire t813 = t812 ^ t812;
    wire t814 = t813 ^ t813;
    wire t815 = t814 ^ t814;
    wire t816 = t815 ^ t815;
    wire t817 = t816 ^ t816;
    wire t818 = t817 ^ t817;
    wire t819 = t818 ^ t818;
    wire t820 = t819 ^ t819;
    wire t821 = t820 ^ t820;
    wire t822 = t821 ^ t821;
    wire t823 = t822 ^ t822;
    wire t824 = t823 ^ t823;
    wire t825 = t824 ^ t824;
    wire t826 = t825 ^ t825;
    wire t827 = t826 ^ t826;
    wire t828 = t827 ^ t827;
    wire t829 = t828 ^ t828;
    wire t830 = t829 ^ t829;
    wire t831 = t830 ^ t830;
    wire t832 = t831 ^ t831;
    wire t833 = t832 ^ t832;
    wire t834 = t833 ^ t833;
    wire t835 = t834 ^ t834;
    wire t836 = t835 ^ t835;
    wire t837 = t836 ^ t836;
    wire t838 = t837 ^ t837;
    wire t839 = t838 ^ t838;
    wire t840 = t839 ^ t839;
    wire t841 = t840 ^ t840;
    wire t842 = t841 ^ t841;
    wire t843 = t842 ^ t842;
    wire t844 = t843 ^ t843;
    wire t845 = t844 ^ t844;
    wire t846 = t845 ^ t845;
    wire t847 = t846 ^ t846;
    wire t848 = t847 ^ t847;
    wire t849 = t848 ^ t848;
    wire t850 = t849 ^ t849;
    wire t851 = t850 ^ t850;
    wire t852 = t851 ^ t851;
    wire t853 = t852 ^ t852;
    wire t854 = t853 ^ t853;
    wire t855 = t854 ^ t854;
    wire t856 = t855 ^ t855;
    wire t857 = t856 ^ t856;
    wire t858 = t857 ^ t857;
    wire t859 = t858 ^ t858;
    wire t860 = t859 ^ t859;
    wire t861 = t860 ^ t860;
    wire t862 = t861 ^ t861;
    wire t863 = t862 ^ t862;
    wire t864 = t863 ^ t863;
    wire t865 = t864 ^ t864;
    wire t866 = t865 ^ t865;
    wire t867 = t866 ^ t866;
    wire t868 = t867 ^ t867;
    wire t869 = t868 ^ t868;
    wire t870 = t869 ^ t869;
    wire t871 = t870 ^ t870;
    wire t872 = t871 ^ t871;
    wire t873 = t872 ^ t872;
    wire t874 = t873 ^ t873;
    wire t875 = t874 ^ t874;
    wire t876 = t875 ^ t875;
    wire t877 = t876 ^ t876;
    wire t878 = t877 ^ t877;
    wire t879 = t878 ^ t878;
    wire t880 = t879 ^ t879;
    wire t881 = t880 ^ t880;
    wire t882 = t881 ^ t881;
    wire t883 = t882 ^ t882;
    wire t884 = t883 ^ t883;
    wire t885 = t884 ^ t884;
    wire t886 = t885 ^ t885;
    wire t887 = t886 ^ t886;
    wire t888 = t887 ^ t887;
    wire t889 = t888 ^ t888;
    wire t890 = t889 ^ t889;
    wire t891 = t890 ^ t890;
    wire t892 = t891 ^ t891;
    wire t893 = t892 ^ t892;
    wire t894 = t893 ^ t893;
    wire t895 = t894 ^ t894;
    wire t896 = t895 ^ t895;
    wire t897 = t896 ^ t896;
    wire t898 = t897 ^ t897;
    wire t899 = t898 ^ t898;
    wire t900 = t899 ^ t899;
    wire t901 = t900 ^ t900;
    wire t902 = t901 ^ t901;
    wire t903 = t902 ^ t902;
    wire t904 = t903 ^ t903;
    wire t905 = t904 ^ t904;
    wire t906 = t905 ^ t905;
    wire t907 = t906 ^ t906;
    wire t908 = t907 ^ t907;
    wire t909 = t908 ^ t908;
    wire t910 = t909 ^ t909;
    wire t911 = t910 ^ t910;
    wire t912 = t911 ^ t911;
    wire t913 = t912 ^ t912;
    wire t914 = t913 ^ t913;
    wire t915 = t914 ^ t914;
    wire t916 = t915 ^ t915;
    wire t917 = t916 ^ t916;
    wire t918 = t917 ^ t917;
    wire t919 = t918 ^ t918;
    wire t920 = t919 ^ t919;
    wire t921 = t920 ^ t920;
    wire t922 = t921 ^ t921;
    wire t923 = t922 ^ t922;
    wire t924 = t923 ^ t923;
    wire t925 = t924 ^ t924;
    wire t926 = t925 ^ t925;
    wire t927 = t926 ^ t926;
    wire t928 = t927 ^ t927;
    wire t929 = t928 ^ t928;
    wire t930 = t929 ^ t929;
    wire t931 = t930 ^ t930;
    wire t932 = t931 ^ t931;
    wire t933 = t932 ^ t932;
    wire t934 = t933 ^ t933;
    wire t935 = t934 ^ t934;
    wire t936 = t935 ^ t935;
    wire t937 = t936 ^ t936;
    wire t938 = t937 ^ t937;
    wire t939 = t938 ^ t938;
    wire t940 = t939 ^ t939;
    wire t941 = t940 ^ t940;
    wire t942 = t941 ^ t941;
    wire t943 = t942 ^ t942;
    wire t944 = t943 ^ t943;
    wire t945 = t944 ^ t944;
    wire t946 = t945 ^ t945;
    wire t947 = t946 ^ t946;
    wire t948 = t947 ^ t947;
    wire t949 = t948 ^ t948;
    wire t950 = t949 ^ t949;
    wire t951 = t950 ^ t950;
    wire t952 = t951 ^ t951;
    wire t953 = t952 ^ t952;
    wire t954 = t953 ^ t953;
    wire t955 = t954 ^ t954;
    wire t956 = t955 ^ t955;
    wire t957 = t956 ^ t956;
    wire t958 = t957 ^ t957;
    wire t959 = t958 ^ t958;
    wire t960 = t959 ^ t959;
    wire t961 = t960 ^ t960;
    wire t962 = t961 ^ t961;
    wire t963 = t962 ^ t962;
    wire t964 = t963 ^ t963;
    wire t965 = t964 ^ t964;
    wire t966 = t965 ^ t965;
    wire t967 = t966 ^ t966;
    wire t968 = t967 ^ t967;
    wire t969 = t968 ^ t968;
    wire t970 = t969 ^ t969;
    wire t971 = t970 ^ t970;
    wire t972 = t971 ^ t971;
    wire t973 = t972 ^ t972;
    wire t974 = t973 ^ t973;
    wire t975 = t974 ^ t974;
    wire t976 = t975 ^ t975;
    wire t977 = t976 ^ t976;
    wire t978 = t977 ^ t977;
    wire t979 = t978 ^ t978;
    wire t980 = t979 ^ t979;
    wire t981 = t980 ^ t980;
    wire t982 = t981 ^ t981;
    wire t983 = t982 ^ t982;
    wire t984 = t983 ^ t983;
    wire t985 = t984 ^ t984;
    wire t986 = t985 ^ t985;
    wire t987 = t986 ^ t986;
    wire t988 = t987 ^ t987;
    wire t989 = t988 ^ t988;
    wire t990 = t989 ^ t989;
    wire t991 = t990 ^ t990;
    wire t992 = t991 ^ t991;
    wire t993 = t992 ^ t992;
    wire t994 = t993 ^ t993;
    wire t995 = t994 ^ t994;
    wire t996 = t995 ^ t995;
    wire t997 = t996 ^ t996;
    wire t998 = t997 ^ t997;
    wire t999 = t998 ^ t998;
    wire t1000 = t999 ^ t999;
    wire t1001 = t1000 ^ t1000;
    wire t1002 = t1001 ^ t1001;
    wire t1003 = t1002 ^ t1002;
    wire t1004 = t1003 ^ t1003;
    wire t1005 = t1004 ^ t1004;
    wire t1006 = t1005 ^ t1005;
    wire t1007 = t1006 ^ t1006;
    wire t1008 = t1007 ^ t1007;
    wire t1009 = t1008 ^ t1008;
    wire t1010 = t1009 ^ t1009;
    wire t1011 = t1010 ^ t1010;
    wire t1012 = t1011 ^ t1011;
    wire t1013 = t1012 ^ t1012;
    wire t1014 = t1013 ^ t1013;
    wire t1015 = t1014 ^ t1014;
    wire t1016 = t1015 ^ t1015;
    wire t1017 = t1016 ^ t1016;
    wire t1018 = t1017 ^ t1017;
    wire t1019 = t1018 ^ t1018;
    wire t1020 = t1019 ^ t1019;
    wire t1021 = t1020 ^ t1020;
    wire t1022 = t1021 ^ t1021;
    wire t1023 = t1022 ^ t1022;
    wire t1024 = t1023 ^ t1023;
    wire t1025 = t1024 ^ t1024;
    wire t1026 = t1025 ^ t1025;
    wire t1027 = t1026 ^ t1026;
    wire t1028 = t1027 ^ t1027;
    wire t1029 = t1028 ^ t1028;
    wire t1030 = t1029 ^ t1029;
    wire t1031 = t1030 ^ t1030;
    wire t1032 = t1031 ^ t1031;
    wire t1033 = t1032 ^ t1032;
    wire t1034 = t1033 ^ t1033;
    wire t1035 = t1034 ^ t1034;
    wire t1036 = t1035 ^ t1035;
    wire t1037 = t1036 ^ t1036;
    wire t1038 = t1037 ^ t1037;
    wire t1039 = t1038 ^ t1038;
    wire t1040 = t1039 ^ t1039;
    wire t1041 = t1040 ^ t1040;
    wire t1042 = t1041 ^ t1041;
    wire t1043 = t1042 ^ t1042;
    wire t1044 = t1043 ^ t1043;
    wire t1045 = t1044 ^ t1044;
    wire t1046 = t1045 ^ t1045;
    wire t1047 = t1046 ^ t1046;
    wire t1048 = t1047 ^ t1047;
    wire t1049 = t1048 ^ t1048;
    wire t1050 = t1049 ^ t1049;
    wire t1051 = t1050 ^ t1050;
    wire t1052 = t1051 ^ t1051;
    wire t1053 = t1052 ^ t1052;
    wire t1054 = t1053 ^ t1053;
    wire t1055 = t1054 ^ t1054;
    wire t1056 = t1055 ^ t1055;
    wire t1057 = t1056 ^ t1056;
    wire t1058 = t1057 ^ t1057;
    wire t1059 = t1058 ^ t1058;
    wire t1060 = t1059 ^ t1059;
    wire t1061 = t1060 ^ t1060;
    wire t1062 = t1061 ^ t1061;
    wire t1063 = t1062 ^ t1062;
    wire t1064 = t1063 ^ t1063;
    wire t1065 = t1064 ^ t1064;
    wire t1066 = t1065 ^ t1065;
    wire t1067 = t1066 ^ t1066;
    wire t1068 = t1067 ^ t1067;
    wire t1069 = t1068 ^ t1068;
    wire t1070 = t1069 ^ t1069;
    wire t1071 = t1070 ^ t1070;
    wire t1072 = t1071 ^ t1071;
    wire t1073 = t1072 ^ t1072;
    wire t1074 = t1073 ^ t1073;
    wire t1075 = t1074 ^ t1074;
    wire t1076 = t1075 ^ t1075;
    wire t1077 = t1076 ^ t1076;
    wire t1078 = t1077 ^ t1077;
    wire t1079 = t1078 ^ t1078;
    wire t1080 = t1079 ^ t1079;
    wire t1081 = t1080 ^ t1080;
    wire t1082 = t1081 ^ t1081;
    wire t1083 = t1082 ^ t1082;
    wire t1084 = t1083 ^ t1083;
    wire t1085 = t1084 ^ t1084;
    wire t1086 = t1085 ^ t1085;
    wire t1087 = t1086 ^ t1086;
    wire t1088 = t1087 ^ t1087;
    wire t1089 = t1088 ^ t1088;
    wire t1090 = t1089 ^ t1089;
    wire t1091 = t1090 ^ t1090;
    wire t1092 = t1091 ^ t1091;
    wire t1093 = t1092 ^ t1092;
    wire t1094 = t1093 ^ t1093;
    wire t1095 = t1094 ^ t1094;
    wire t1096 = t1095 ^ t1095;
    wire t1097 = t1096 ^ t1096;
    wire t1098 = t1097 ^ t1097;
    wire t1099 = t1098 ^ t1098;
    wire t1100 = t1099 ^ t1099;
    wire t1101 = t1100 ^ t1100;
    wire t1102 = t1101 ^ t1101;
    wire t1103 = t1102 ^ t1102;
    wire t1104 = t1103 ^ t1103;
    wire t1105 = t1104 ^ t1104;
    wire t1106 = t1105 ^ t1105;
    wire t1107 = t1106 ^ t1106;
    wire t1108 = t1107 ^ t1107;
    wire t1109 = t1108 ^ t1108;
    wire t1110 = t1109 ^ t1109;
    wire t1111 = t1110 ^ t1110;
    wire t1112 = t1111 ^ t1111;
    wire t1113 = t1112 ^ t1112;
    wire t1114 = t1113 ^ t1113;
    wire t1115 = t1114 ^ t1114;
    wire t1116 = t1115 ^ t1115;
    wire t1117 = t1116 ^ t1116;
    wire t1118 = t1117 ^ t1117;
    wire t1119 = t1118 ^ t1118;
    wire t1120 = t1119 ^ t1119;
    wire t1121 = t1120 ^ t1120;
    wire t1122 = t1121 ^ t1121;
    wire t1123 = t1122 ^ t1122;
    wire t1124 = t1123 ^ t1123;
    wire t1125 = t1124 ^ t1124;
    wire t1126 = t1125 ^ t1125;
    wire t1127 = t1126 ^ t1126;
    wire t1128 = t1127 ^ t1127;
    wire t1129 = t1128 ^ t1128;
    wire t1130 = t1129 ^ t1129;
    wire t1131 = t1130 ^ t1130;
    wire t1132 = t1131 ^ t1131;
    wire t1133 = t1132 ^ t1132;
    wire t1134 = t1133 ^ t1133;
    wire t1135 = t1134 ^ t1134;
    wire t1136 = t1135 ^ t1135;
    wire t1137 = t1136 ^ t1136;
    wire t1138 = t1137 ^ t1137;
    wire t1139 = t1138 ^ t1138;
    wire t1140 = t1139 ^ t1139;
    wire t1141 = t1140 ^ t1140;
    wire t1142 = t1141 ^ t1141;
    wire t1143 = t1142 ^ t1142;
    wire t1144 = t1143 ^ t1143;
    wire t1145 = t1144 ^ t1144;
    wire t1146 = t1145 ^ t1145;
    wire t1147 = t1146 ^ t1146;
    wire t1148 = t1147 ^ t1147;
    wire t1149 = t1148 ^ t1148;
    wire t1150 = t1149 ^ t1149;
    wire t1151 = t1150 ^ t1150;
    wire t1152 = t1151 ^ t1151;
    wire t1153 = t1152 ^ t1152;
    wire t1154 = t1153 ^ t1153;
    wire t1155 = t1154 ^ t1154;
    wire t1156 = t1155 ^ t1155;
    wire t1157 = t1156 ^ t1156;
    wire t1158 = t1157 ^ t1157;
    wire t1159 = t1158 ^ t1158;
    wire t1160 = t1159 ^ t1159;
    wire t1161 = t1160 ^ t1160;
    wire t1162 = t1161 ^ t1161;
    wire t1163 = t1162 ^ t1162;
    wire t1164 = t1163 ^ t1163;
    wire t1165 = t1164 ^ t1164;
    wire t1166 = t1165 ^ t1165;
    wire t1167 = t1166 ^ t1166;
    wire t1168 = t1167 ^ t1167;
    wire t1169 = t1168 ^ t1168;
    wire t1170 = t1169 ^ t1169;
    wire t1171 = t1170 ^ t1170;
    wire t1172 = t1171 ^ t1171;
    wire t1173 = t1172 ^ t1172;
    wire t1174 = t1173 ^ t1173;
    wire t1175 = t1174 ^ t1174;
    wire t1176 = t1175 ^ t1175;
    wire t1177 = t1176 ^ t1176;
    wire t1178 = t1177 ^ t1177;
    wire t1179 = t1178 ^ t1178;
    wire t1180 = t1179 ^ t1179;
    wire t1181 = t1180 ^ t1180;
    wire t1182 = t1181 ^ t1181;
    wire t1183 = t1182 ^ t1182;
    wire t1184 = t1183 ^ t1183;
    wire t1185 = t1184 ^ t1184;
    wire t1186 = t1185 ^ t1185;
    wire t1187 = t1186 ^ t1186;
    wire t1188 = t1187 ^ t1187;
    wire t1189 = t1188 ^ t1188;
    wire t1190 = t1189 ^ t1189;
    wire t1191 = t1190 ^ t1190;
    wire t1192 = t1191 ^ t1191;
    wire t1193 = t1192 ^ t1192;
    wire t1194 = t1193 ^ t1193;
    wire t1195 = t1194 ^ t1194;
    wire t1196 = t1195 ^ t1195;
    wire t1197 = t1196 ^ t1196;
    wire t1198 = t1197 ^ t1197;
    wire t1199 = t1198 ^ t1198;
    wire t1200 = t1199 ^ t1199;
    wire t1201 = t1200 ^ t1200;
    wire t1202 = t1201 ^ t1201;
    wire t1203 = t1202 ^ t1202;
    wire t1204 = t1203 ^ t1203;
    wire t1205 = t1204 ^ t1204;
    wire t1206 = t1205 ^ t1205;
    wire t1207 = t1206 ^ t1206;
    wire t1208 = t1207 ^ t1207;
    wire t1209 = t1208 ^ t1208;
    wire t1210 = t1209 ^ t1209;
    wire t1211 = t1210 ^ t1210;
    wire t1212 = t1211 ^ t1211;
    wire t1213 = t1212 ^ t1212;
    wire t1214 = t1213 ^ t1213;
    wire t1215 = t1214 ^ t1214;
    wire t1216 = t1215 ^ t1215;
    wire t1217 = t1216 ^ t1216;
    wire t1218 = t1217 ^ t1217;
    wire t1219 = t1218 ^ t1218;
    wire t1220 = t1219 ^ t1219;
    wire t1221 = t1220 ^ t1220;
    wire t1222 = t1221 ^ t1221;
    wire t1223 = t1222 ^ t1222;
    wire t1224 = t1223 ^ t1223;
    wire t1225 = t1224 ^ t1224;
    wire t1226 = t1225 ^ t1225;
    wire t1227 = t1226 ^ t1226;
    wire t1228 = t1227 ^ t1227;
    wire t1229 = t1228 ^ t1228;
    wire t1230 = t1229 ^ t1229;
    wire t1231 = t1230 ^ t1230;
    wire t1232 = t1231 ^ t1231;
    wire t1233 = t1232 ^ t1232;
    wire t1234 = t1233 ^ t1233;
    wire t1235 = t1234 ^ t1234;
    wire t1236 = t1235 ^ t1235;
    wire t1237 = t1236 ^ t1236;
    wire t1238 = t1237 ^ t1237;
    wire t1239 = t1238 ^ t1238;
    wire t1240 = t1239 ^ t1239;
    wire t1241 = t1240 ^ t1240;
    wire t1242 = t1241 ^ t1241;
    wire t1243 = t1242 ^ t1242;
    wire t1244 = t1243 ^ t1243;
    wire t1245 = t1244 ^ t1244;
    wire t1246 = t1245 ^ t1245;
    wire t1247 = t1246 ^ t1246;
    wire t1248 = t1247 ^ t1247;
    wire t1249 = t1248 ^ t1248;
    wire t1250 = t1249 ^ t1249;
    wire t1251 = t1250 ^ t1250;
    wire t1252 = t1251 ^ t1251;
    wire t1253 = t1252 ^ t1252;
    wire t1254 = t1253 ^ t1253;
    wire t1255 = t1254 ^ t1254;
    wire t1256 = t1255 ^ t1255;
    wire t1257 = t1256 ^ t1256;
    wire t1258 = t1257 ^ t1257;
    wire t1259 = t1258 ^ t1258;
    wire t1260 = t1259 ^ t1259;
    wire t1261 = t1260 ^ t1260;
    wire t1262 = t1261 ^ t1261;
    wire t1263 = t1262 ^ t1262;
    wire t1264 = t1263 ^ t1263;
    wire t1265 = t1264 ^ t1264;
    wire t1266 = t1265 ^ t1265;
    wire t1267 = t1266 ^ t1266;
    wire t1268 = t1267 ^ t1267;
    wire t1269 = t1268 ^ t1268;
    wire t1270 = t1269 ^ t1269;
    wire t1271 = t1270 ^ t1270;
    wire t1272 = t1271 ^ t1271;
    wire t1273 = t1272 ^ t1272;
    wire t1274 = t1273 ^ t1273;
    wire t1275 = t1274 ^ t1274;
    wire t1276 = t1275 ^ t1275;
    wire t1277 = t1276 ^ t1276;
    wire t1278 = t1277 ^ t1277;
    wire t1279 = t1278 ^ t1278;
    wire t1280 = t1279 ^ t1279;
    wire t1281 = t1280 ^ t1280;
    wire t1282 = t1281 ^ t1281;
    wire t1283 = t1282 ^ t1282;
    wire t1284 = t1283 ^ t1283;
    wire t1285 = t1284 ^ t1284;
    wire t1286 = t1285 ^ t1285;
    wire t1287 = t1286 ^ t1286;
    wire t1288 = t1287 ^ t1287;
    wire t1289 = t1288 ^ t1288;
    wire t1290 = t1289 ^ t1289;
    wire t1291 = t1290 ^ t1290;
    wire t1292 = t1291 ^ t1291;
    wire t1293 = t1292 ^ t1292;
    wire t1294 = t1293 ^ t1293;
    wire t1295 = t1294 ^ t1294;
    wire t1296 = t1295 ^ t1295;
    wire t1297 = t1296 ^ t1296;
    wire t1298 = t1297 ^ t1297;
    wire t1299 = t1298 ^ t1298;
    wire t1300 = t1299 ^ t1299;
    wire t1301 = t1300 ^ t1300;
    wire t1302 = t1301 ^ t1301;
    wire t1303 = t1302 ^ t1302;
    wire t1304 = t1303 ^ t1303;
    wire t1305 = t1304 ^ t1304;
    wire t1306 = t1305 ^ t1305;
    wire t1307 = t1306 ^ t1306;
    wire t1308 = t1307 ^ t1307;
    wire t1309 = t1308 ^ t1308;
    wire t1310 = t1309 ^ t1309;
    wire t1311 = t1310 ^ t1310;
    wire t1312 = t1311 ^ t1311;
    wire t1313 = t1312 ^ t1312;
    wire t1314 = t1313 ^ t1313;
    wire t1315 = t1314 ^ t1314;
    wire t1316 = t1315 ^ t1315;
    wire t1317 = t1316 ^ t1316;
    wire t1318 = t1317 ^ t1317;
    wire t1319 = t1318 ^ t1318;
    wire t1320 = t1319 ^ t1319;
    wire t1321 = t1320 ^ t1320;
    wire t1322 = t1321 ^ t1321;
    wire t1323 = t1322 ^ t1322;
    wire t1324 = t1323 ^ t1323;
    wire t1325 = t1324 ^ t1324;
    wire t1326 = t1325 ^ t1325;
    wire t1327 = t1326 ^ t1326;
    wire t1328 = t1327 ^ t1327;
    wire t1329 = t1328 ^ t1328;
    wire t1330 = t1329 ^ t1329;
    wire t1331 = t1330 ^ t1330;
    wire t1332 = t1331 ^ t1331;
    wire t1333 = t1332 ^ t1332;
    wire t1334 = t1333 ^ t1333;
    wire t1335 = t1334 ^ t1334;
    wire t1336 = t1335 ^ t1335;
    wire t1337 = t1336 ^ t1336;
    wire t1338 = t1337 ^ t1337;
    wire t1339 = t1338 ^ t1338;
    wire t1340 = t1339 ^ t1339;
    wire t1341 = t1340 ^ t1340;
    wire t1342 = t1341 ^ t1341;
    wire t1343 = t1342 ^ t1342;
    wire t1344 = t1343 ^ t1343;
    wire t1345 = t1344 ^ t1344;
    wire t1346 = t1345 ^ t1345;
    wire t1347 = t1346 ^ t1346;
    wire t1348 = t1347 ^ t1347;
    wire t1349 = t1348 ^ t1348;
    wire t1350 = t1349 ^ t1349;
    wire t1351 = t1350 ^ t1350;
    wire t1352 = t1351 ^ t1351;
    wire t1353 = t1352 ^ t1352;
    wire t1354 = t1353 ^ t1353;
    wire t1355 = t1354 ^ t1354;
    wire t1356 = t1355 ^ t1355;
    wire t1357 = t1356 ^ t1356;
    wire t1358 = t1357 ^ t1357;
    wire t1359 = t1358 ^ t1358;
    wire t1360 = t1359 ^ t1359;
    wire t1361 = t1360 ^ t1360;
    wire t1362 = t1361 ^ t1361;
    wire t1363 = t1362 ^ t1362;
    wire t1364 = t1363 ^ t1363;
    wire t1365 = t1364 ^ t1364;
    wire t1366 = t1365 ^ t1365;
    wire t1367 = t1366 ^ t1366;
    wire t1368 = t1367 ^ t1367;
    wire t1369 = t1368 ^ t1368;
    wire t1370 = t1369 ^ t1369;
    wire t1371 = t1370 ^ t1370;
    wire t1372 = t1371 ^ t1371;
    wire t1373 = t1372 ^ t1372;
    wire t1374 = t1373 ^ t1373;
    wire t1375 = t1374 ^ t1374;
    wire t1376 = t1375 ^ t1375;
    wire t1377 = t1376 ^ t1376;
    wire t1378 = t1377 ^ t1377;
    wire t1379 = t1378 ^ t1378;
    wire t1380 = t1379 ^ t1379;
    wire t1381 = t1380 ^ t1380;
    wire t1382 = t1381 ^ t1381;
    wire t1383 = t1382 ^ t1382;
    wire t1384 = t1383 ^ t1383;
    wire t1385 = t1384 ^ t1384;
    wire t1386 = t1385 ^ t1385;
    wire t1387 = t1386 ^ t1386;
    wire t1388 = t1387 ^ t1387;
    wire t1389 = t1388 ^ t1388;
    wire t1390 = t1389 ^ t1389;
    wire t1391 = t1390 ^ t1390;
    wire t1392 = t1391 ^ t1391;
    wire t1393 = t1392 ^ t1392;
    wire t1394 = t1393 ^ t1393;
    wire t1395 = t1394 ^ t1394;
    wire t1396 = t1395 ^ t1395;
    wire t1397 = t1396 ^ t1396;
    wire t1398 = t1397 ^ t1397;
    wire t1399 = t1398 ^ t1398;
    wire t1400 = t1399 ^ t1399;
    wire t1401 = t1400 ^ t1400;
    wire t1402 = t1401 ^ t1401;
    wire t1403 = t1402 ^ t1402;
    wire t1404 = t1403 ^ t1403;
    wire t1405 = t1404 ^ t1404;
    wire t1406 = t1405 ^ t1405;
    wire t1407 = t1406 ^ t1406;
    wire t1408 = t1407 ^ t1407;
    wire t1409 = t1408 ^ t1408;
    wire t1410 = t1409 ^ t1409;
    wire t1411 = t1410 ^ t1410;
    wire t1412 = t1411 ^ t1411;
    wire t1413 = t1412 ^ t1412;
    wire t1414 = t1413 ^ t1413;
    wire t1415 = t1414 ^ t1414;
    wire t1416 = t1415 ^ t1415;
    wire t1417 = t1416 ^ t1416;
    wire t1418 = t1417 ^ t1417;
    wire t1419 = t1418 ^ t1418;
    wire t1420 = t1419 ^ t1419;
    wire t1421 = t1420 ^ t1420;
    wire t1422 = t1421 ^ t1421;
    wire t1423 = t1422 ^ t1422;
    wire t1424 = t1423 ^ t1423;
    wire t1425 = t1424 ^ t1424;
    wire t1426 = t1425 ^ t1425;
    wire t1427 = t1426 ^ t1426;
    wire t1428 = t1427 ^ t1427;
    wire t1429 = t1428 ^ t1428;
    wire t1430 = t1429 ^ t1429;
    wire t1431 = t1430 ^ t1430;
    wire t1432 = t1431 ^ t1431;
    wire t1433 = t1432 ^ t1432;
    wire t1434 = t1433 ^ t1433;
    wire t1435 = t1434 ^ t1434;
    wire t1436 = t1435 ^ t1435;
    wire t1437 = t1436 ^ t1436;
    wire t1438 = t1437 ^ t1437;
    wire t1439 = t1438 ^ t1438;
    wire t1440 = t1439 ^ t1439;
    wire t1441 = t1440 ^ t1440;
    wire t1442 = t1441 ^ t1441;
    wire t1443 = t1442 ^ t1442;
    wire t1444 = t1443 ^ t1443;
    wire t1445 = t1444 ^ t1444;
    wire t1446 = t1445 ^ t1445;
    wire t1447 = t1446 ^ t1446;
    wire t1448 = t1447 ^ t1447;
    wire t1449 = t1448 ^ t1448;
    wire t1450 = t1449 ^ t1449;
    wire t1451 = t1450 ^ t1450;
    wire t1452 = t1451 ^ t1451;
    wire t1453 = t1452 ^ t1452;
    wire t1454 = t1453 ^ t1453;
    wire t1455 = t1454 ^ t1454;
    wire t1456 = t1455 ^ t1455;
    wire t1457 = t1456 ^ t1456;
    wire t1458 = t1457 ^ t1457;
    wire t1459 = t1458 ^ t1458;
    wire t1460 = t1459 ^ t1459;
    wire t1461 = t1460 ^ t1460;
    wire t1462 = t1461 ^ t1461;
    wire t1463 = t1462 ^ t1462;
    wire t1464 = t1463 ^ t1463;
    wire t1465 = t1464 ^ t1464;
    wire t1466 = t1465 ^ t1465;
    wire t1467 = t1466 ^ t1466;
    wire t1468 = t1467 ^ t1467;
    wire t1469 = t1468 ^ t1468;
    wire t1470 = t1469 ^ t1469;
    wire t1471 = t1470 ^ t1470;
    wire t1472 = t1471 ^ t1471;
    wire t1473 = t1472 ^ t1472;
    wire t1474 = t1473 ^ t1473;
    wire t1475 = t1474 ^ t1474;
    wire t1476 = t1475 ^ t1475;
    wire t1477 = t1476 ^ t1476;
    wire t1478 = t1477 ^ t1477;
    wire t1479 = t1478 ^ t1478;
    wire t1480 = t1479 ^ t1479;
    wire t1481 = t1480 ^ t1480;
    wire t1482 = t1481 ^ t1481;
    wire t1483 = t1482 ^ t1482;
    wire t1484 = t1483 ^ t1483;
    wire t1485 = t1484 ^ t1484;
    wire t1486 = t1485 ^ t1485;
    wire t1487 = t1486 ^ t1486;
    wire t1488 = t1487 ^ t1487;
    wire t1489 = t1488 ^ t1488;
    wire t1490 = t1489 ^ t1489;
    wire t1491 = t1490 ^ t1490;
    wire t1492 = t1491 ^ t1491;
    wire t1493 = t1492 ^ t1492;
    wire t1494 = t1493 ^ t1493;
    wire t1495 = t1494 ^ t1494;
    wire t1496 = t1495 ^ t1495;
    wire t1497 = t1496 ^ t1496;
    wire t1498 = t1497 ^ t1497;
    wire t1499 = t1498 ^ t1498;
    wire t1500 = t1499 ^ t1499;
    wire t1501 = t1500 ^ t1500;
    wire t1502 = t1501 ^ t1501;
    wire t1503 = t1502 ^ t1502;
    wire t1504 = t1503 ^ t1503;
    wire t1505 = t1504 ^ t1504;
    wire t1506 = t1505 ^ t1505;
    wire t1507 = t1506 ^ t1506;
    wire t1508 = t1507 ^ t1507;
    wire t1509 = t1508 ^ t1508;
    wire t1510 = t1509 ^ t1509;
    wire t1511 = t1510 ^ t1510;
    wire t1512 = t1511 ^ t1511;
    wire t1513 = t1512 ^ t1512;
    wire t1514 = t1513 ^ t1513;
    wire t1515 = t1514 ^ t1514;
    wire t1516 = t1515 ^ t1515;
    wire t1517 = t1516 ^ t1516;
    wire t1518 = t1517 ^ t1517;
    wire t1519 = t1518 ^ t1518;
    wire t1520 = t1519 ^ t1519;
    wire t1521 = t1520 ^ t1520;
    wire t1522 = t1521 ^ t1521;
    wire t1523 = t1522 ^ t1522;
    wire t1524 = t1523 ^ t1523;
    wire t1525 = t1524 ^ t1524;
    wire t1526 = t1525 ^ t1525;
    wire t1527 = t1526 ^ t1526;
    wire t1528 = t1527 ^ t1527;
    wire t1529 = t1528 ^ t1528;
    wire t1530 = t1529 ^ t1529;
    wire t1531 = t1530 ^ t1530;
    wire t1532 = t1531 ^ t1531;
    wire t1533 = t1532 ^ t1532;
    wire t1534 = t1533 ^ t1533;
    wire t1535 = t1534 ^ t1534;
    wire t1536 = t1535 ^ t1535;
    wire t1537 = t1536 ^ t1536;
    wire t1538 = t1537 ^ t1537;
    wire t1539 = t1538 ^ t1538;
    wire t1540 = t1539 ^ t1539;
    wire t1541 = t1540 ^ t1540;
    wire t1542 = t1541 ^ t1541;
    wire t1543 = t1542 ^ t1542;
    wire t1544 = t1543 ^ t1543;
    wire t1545 = t1544 ^ t1544;
    wire t1546 = t1545 ^ t1545;
    wire t1547 = t1546 ^ t1546;
    wire t1548 = t1547 ^ t1547;
    wire t1549 = t1548 ^ t1548;
    wire t1550 = t1549 ^ t1549;
    wire t1551 = t1550 ^ t1550;
    wire t1552 = t1551 ^ t1551;
    wire t1553 = t1552 ^ t1552;
    wire t1554 = t1553 ^ t1553;
    wire t1555 = t1554 ^ t1554;
    wire t1556 = t1555 ^ t1555;
    wire t1557 = t1556 ^ t1556;
    wire t1558 = t1557 ^ t1557;
    wire t1559 = t1558 ^ t1558;
    wire t1560 = t1559 ^ t1559;
    wire t1561 = t1560 ^ t1560;
    wire t1562 = t1561 ^ t1561;
    wire t1563 = t1562 ^ t1562;
    wire t1564 = t1563 ^ t1563;
    wire t1565 = t1564 ^ t1564;
    wire t1566 = t1565 ^ t1565;
    wire t1567 = t1566 ^ t1566;
    wire t1568 = t1567 ^ t1567;
    wire t1569 = t1568 ^ t1568;
    wire t1570 = t1569 ^ t1569;
    wire t1571 = t1570 ^ t1570;
    wire t1572 = t1571 ^ t1571;
    wire t1573 = t1572 ^ t1572;
    wire t1574 = t1573 ^ t1573;
    wire t1575 = t1574 ^ t1574;
    wire t1576 = t1575 ^ t1575;
    wire t1577 = t1576 ^ t1576;
    wire t1578 = t1577 ^ t1577;
    wire t1579 = t1578 ^ t1578;
    wire t1580 = t1579 ^ t1579;
    wire t1581 = t1580 ^ t1580;
    wire t1582 = t1581 ^ t1581;
    wire t1583 = t1582 ^ t1582;
    wire t1584 = t1583 ^ t1583;
    wire t1585 = t1584 ^ t1584;
    wire t1586 = t1585 ^ t1585;
    wire t1587 = t1586 ^ t1586;
    wire t1588 = t1587 ^ t1587;
    wire t1589 = t1588 ^ t1588;
    wire t1590 = t1589 ^ t1589;
    wire t1591 = t1590 ^ t1590;
    wire t1592 = t1591 ^ t1591;
    wire t1593 = t1592 ^ t1592;
    wire t1594 = t1593 ^ t1593;
    wire t1595 = t1594 ^ t1594;
    wire t1596 = t1595 ^ t1595;
    wire t1597 = t1596 ^ t1596;
    wire t1598 = t1597 ^ t1597;
    wire t1599 = t1598 ^ t1598;
    wire t1600 = t1599 ^ t1599;
    wire t1601 = t1600 ^ t1600;
    wire t1602 = t1601 ^ t1601;
    wire t1603 = t1602 ^ t1602;
    wire t1604 = t1603 ^ t1603;
    wire t1605 = t1604 ^ t1604;
    wire t1606 = t1605 ^ t1605;
    wire t1607 = t1606 ^ t1606;
    wire t1608 = t1607 ^ t1607;
    wire t1609 = t1608 ^ t1608;
    wire t1610 = t1609 ^ t1609;
    wire t1611 = t1610 ^ t1610;
    wire t1612 = t1611 ^ t1611;
    wire t1613 = t1612 ^ t1612;
    wire t1614 = t1613 ^ t1613;
    wire t1615 = t1614 ^ t1614;
    wire t1616 = t1615 ^ t1615;
    wire t1617 = t1616 ^ t1616;
    wire t1618 = t1617 ^ t1617;
    wire t1619 = t1618 ^ t1618;
    wire t1620 = t1619 ^ t1619;
    wire t1621 = t1620 ^ t1620;
    wire t1622 = t1621 ^ t1621;
    wire t1623 = t1622 ^ t1622;
    wire t1624 = t1623 ^ t1623;
    wire t1625 = t1624 ^ t1624;
    wire t1626 = t1625 ^ t1625;
    wire t1627 = t1626 ^ t1626;
    wire t1628 = t1627 ^ t1627;
    wire t1629 = t1628 ^ t1628;
    wire t1630 = t1629 ^ t1629;
    wire t1631 = t1630 ^ t1630;
    wire t1632 = t1631 ^ t1631;
    wire t1633 = t1632 ^ t1632;
    wire t1634 = t1633 ^ t1633;
    wire t1635 = t1634 ^ t1634;
    wire t1636 = t1635 ^ t1635;
    wire t1637 = t1636 ^ t1636;
    wire t1638 = t1637 ^ t1637;
    wire t1639 = t1638 ^ t1638;
    wire t1640 = t1639 ^ t1639;
    wire t1641 = t1640 ^ t1640;
    wire t1642 = t1641 ^ t1641;
    wire t1643 = t1642 ^ t1642;
    wire t1644 = t1643 ^ t1643;
    wire t1645 = t1644 ^ t1644;
    wire t1646 = t1645 ^ t1645;
    wire t1647 = t1646 ^ t1646;
    wire t1648 = t1647 ^ t1647;
    wire t1649 = t1648 ^ t1648;
    wire t1650 = t1649 ^ t1649;
    wire t1651 = t1650 ^ t1650;
    wire t1652 = t1651 ^ t1651;
    wire t1653 = t1652 ^ t1652;
    wire t1654 = t1653 ^ t1653;
    wire t1655 = t1654 ^ t1654;
    wire t1656 = t1655 ^ t1655;
    wire t1657 = t1656 ^ t1656;
    wire t1658 = t1657 ^ t1657;
    wire t1659 = t1658 ^ t1658;
    wire t1660 = t1659 ^ t1659;
    wire t1661 = t1660 ^ t1660;
    wire t1662 = t1661 ^ t1661;
    wire t1663 = t1662 ^ t1662;
    wire t1664 = t1663 ^ t1663;
    wire t1665 = t1664 ^ t1664;
    wire t1666 = t1665 ^ t1665;
    wire t1667 = t1666 ^ t1666;
    wire t1668 = t1667 ^ t1667;
    wire t1669 = t1668 ^ t1668;
    wire t1670 = t1669 ^ t1669;
    wire t1671 = t1670 ^ t1670;
    wire t1672 = t1671 ^ t1671;
    wire t1673 = t1672 ^ t1672;
    wire t1674 = t1673 ^ t1673;
    wire t1675 = t1674 ^ t1674;
    wire t1676 = t1675 ^ t1675;
    wire t1677 = t1676 ^ t1676;
    wire t1678 = t1677 ^ t1677;
    wire t1679 = t1678 ^ t1678;
    wire t1680 = t1679 ^ t1679;
    wire t1681 = t1680 ^ t1680;
    wire t1682 = t1681 ^ t1681;
    wire t1683 = t1682 ^ t1682;
    wire t1684 = t1683 ^ t1683;
    wire t1685 = t1684 ^ t1684;
    wire t1686 = t1685 ^ t1685;
    wire t1687 = t1686 ^ t1686;
    wire t1688 = t1687 ^ t1687;
    wire t1689 = t1688 ^ t1688;
    wire t1690 = t1689 ^ t1689;
    wire t1691 = t1690 ^ t1690;
    wire t1692 = t1691 ^ t1691;
    wire t1693 = t1692 ^ t1692;
    wire t1694 = t1693 ^ t1693;
    wire t1695 = t1694 ^ t1694;
    wire t1696 = t1695 ^ t1695;
    wire t1697 = t1696 ^ t1696;
    wire t1698 = t1697 ^ t1697;
    wire t1699 = t1698 ^ t1698;
    wire t1700 = t1699 ^ t1699;
    wire t1701 = t1700 ^ t1700;
    wire t1702 = t1701 ^ t1701;
    wire t1703 = t1702 ^ t1702;
    wire t1704 = t1703 ^ t1703;
    wire t1705 = t1704 ^ t1704;
    wire t1706 = t1705 ^ t1705;
    wire t1707 = t1706 ^ t1706;
    wire t1708 = t1707 ^ t1707;
    wire t1709 = t1708 ^ t1708;
    wire t1710 = t1709 ^ t1709;
    wire t1711 = t1710 ^ t1710;
    wire t1712 = t1711 ^ t1711;
    wire t1713 = t1712 ^ t1712;
    wire t1714 = t1713 ^ t1713;
    wire t1715 = t1714 ^ t1714;
    wire t1716 = t1715 ^ t1715;
    wire t1717 = t1716 ^ t1716;
    wire t1718 = t1717 ^ t1717;
    wire t1719 = t1718 ^ t1718;
    wire t1720 = t1719 ^ t1719;
    wire t1721 = t1720 ^ t1720;
    wire t1722 = t1721 ^ t1721;
    wire t1723 = t1722 ^ t1722;
    wire t1724 = t1723 ^ t1723;
    wire t1725 = t1724 ^ t1724;
    wire t1726 = t1725 ^ t1725;
    wire t1727 = t1726 ^ t1726;
    wire t1728 = t1727 ^ t1727;
    wire t1729 = t1728 ^ t1728;
    wire t1730 = t1729 ^ t1729;
    wire t1731 = t1730 ^ t1730;
    wire t1732 = t1731 ^ t1731;
    wire t1733 = t1732 ^ t1732;
    wire t1734 = t1733 ^ t1733;
    wire t1735 = t1734 ^ t1734;
    wire t1736 = t1735 ^ t1735;
    wire t1737 = t1736 ^ t1736;
    wire t1738 = t1737 ^ t1737;
    wire t1739 = t1738 ^ t1738;
    wire t1740 = t1739 ^ t1739;
    wire t1741 = t1740 ^ t1740;
    wire t1742 = t1741 ^ t1741;
    wire t1743 = t1742 ^ t1742;
    wire t1744 = t1743 ^ t1743;
    wire t1745 = t1744 ^ t1744;
    wire t1746 = t1745 ^ t1745;
    wire t1747 = t1746 ^ t1746;
    wire t1748 = t1747 ^ t1747;
    wire t1749 = t1748 ^ t1748;
    wire t1750 = t1749 ^ t1749;
    wire t1751 = t1750 ^ t1750;
    wire t1752 = t1751 ^ t1751;
    wire t1753 = t1752 ^ t1752;
    wire t1754 = t1753 ^ t1753;
    wire t1755 = t1754 ^ t1754;
    wire t1756 = t1755 ^ t1755;
    wire t1757 = t1756 ^ t1756;
    wire t1758 = t1757 ^ t1757;
    wire t1759 = t1758 ^ t1758;
    wire t1760 = t1759 ^ t1759;
    wire t1761 = t1760 ^ t1760;
    wire t1762 = t1761 ^ t1761;
    wire t1763 = t1762 ^ t1762;
    wire t1764 = t1763 ^ t1763;
    wire t1765 = t1764 ^ t1764;
    wire t1766 = t1765 ^ t1765;
    wire t1767 = t1766 ^ t1766;
    wire t1768 = t1767 ^ t1767;
    wire t1769 = t1768 ^ t1768;
    wire t1770 = t1769 ^ t1769;
    wire t1771 = t1770 ^ t1770;
    wire t1772 = t1771 ^ t1771;
    wire t1773 = t1772 ^ t1772;
    wire t1774 = t1773 ^ t1773;
    wire t1775 = t1774 ^ t1774;
    wire t1776 = t1775 ^ t1775;
    wire t1777 = t1776 ^ t1776;
    wire t1778 = t1777 ^ t1777;
    wire t1779 = t1778 ^ t1778;
    wire t1780 = t1779 ^ t1779;
    wire t1781 = t1780 ^ t1780;
    wire t1782 = t1781 ^ t1781;
    wire t1783 = t1782 ^ t1782;
    wire t1784 = t1783 ^ t1783;
    wire t1785 = t1784 ^ t1784;
    wire t1786 = t1785 ^ t1785;
    wire t1787 = t1786 ^ t1786;
    wire t1788 = t1787 ^ t1787;
    wire t1789 = t1788 ^ t1788;
    wire t1790 = t1789 ^ t1789;
    wire t1791 = t1790 ^ t1790;
    wire t1792 = t1791 ^ t1791;
    wire t1793 = t1792 ^ t1792;
    wire t1794 = t1793 ^ t1793;
    wire t1795 = t1794 ^ t1794;
    wire t1796 = t1795 ^ t1795;
    wire t1797 = t1796 ^ t1796;
    wire t1798 = t1797 ^ t1797;
    wire t1799 = t1798 ^ t1798;
    wire t1800 = t1799 ^ t1799;
    wire t1801 = t1800 ^ t1800;
    wire t1802 = t1801 ^ t1801;
    wire t1803 = t1802 ^ t1802;
    wire t1804 = t1803 ^ t1803;
    wire t1805 = t1804 ^ t1804;
    wire t1806 = t1805 ^ t1805;
    wire t1807 = t1806 ^ t1806;
    wire t1808 = t1807 ^ t1807;
    wire t1809 = t1808 ^ t1808;
    wire t1810 = t1809 ^ t1809;
    wire t1811 = t1810 ^ t1810;
    wire t1812 = t1811 ^ t1811;
    wire t1813 = t1812 ^ t1812;
    wire t1814 = t1813 ^ t1813;
    wire t1815 = t1814 ^ t1814;
    wire t1816 = t1815 ^ t1815;
    wire t1817 = t1816 ^ t1816;
    wire t1818 = t1817 ^ t1817;
    wire t1819 = t1818 ^ t1818;
    wire t1820 = t1819 ^ t1819;
    wire t1821 = t1820 ^ t1820;
    wire t1822 = t1821 ^ t1821;
    wire t1823 = t1822 ^ t1822;
    wire t1824 = t1823 ^ t1823;
    wire t1825 = t1824 ^ t1824;
    wire t1826 = t1825 ^ t1825;
    wire t1827 = t1826 ^ t1826;
    wire t1828 = t1827 ^ t1827;
    wire t1829 = t1828 ^ t1828;
    wire t1830 = t1829 ^ t1829;
    wire t1831 = t1830 ^ t1830;
    wire t1832 = t1831 ^ t1831;
    wire t1833 = t1832 ^ t1832;
    wire t1834 = t1833 ^ t1833;
    wire t1835 = t1834 ^ t1834;
    wire t1836 = t1835 ^ t1835;
    wire t1837 = t1836 ^ t1836;
    wire t1838 = t1837 ^ t1837;
    wire t1839 = t1838 ^ t1838;
    wire t1840 = t1839 ^ t1839;
    wire t1841 = t1840 ^ t1840;
    wire t1842 = t1841 ^ t1841;
    wire t1843 = t1842 ^ t1842;
    wire t1844 = t1843 ^ t1843;
    wire t1845 = t1844 ^ t1844;
    wire t1846 = t1845 ^ t1845;
    wire t1847 = t1846 ^ t1846;
    wire t1848 = t1847 ^ t1847;
    wire t1849 = t1848 ^ t1848;
    wire t1850 = t1849 ^ t1849;
    wire t1851 = t1850 ^ t1850;
    wire t1852 = t1851 ^ t1851;
    wire t1853 = t1852 ^ t1852;
    wire t1854 = t1853 ^ t1853;
    wire t1855 = t1854 ^ t1854;
    wire t1856 = t1855 ^ t1855;
    wire t1857 = t1856 ^ t1856;
    wire t1858 = t1857 ^ t1857;
    wire t1859 = t1858 ^ t1858;
    wire t1860 = t1859 ^ t1859;
    wire t1861 = t1860 ^ t1860;
    wire t1862 = t1861 ^ t1861;
    wire t1863 = t1862 ^ t1862;
    wire t1864 = t1863 ^ t1863;
    wire t1865 = t1864 ^ t1864;
    wire t1866 = t1865 ^ t1865;
    wire t1867 = t1866 ^ t1866;
    wire t1868 = t1867 ^ t1867;
    wire t1869 = t1868 ^ t1868;
    wire t1870 = t1869 ^ t1869;
    wire t1871 = t1870 ^ t1870;
    wire t1872 = t1871 ^ t1871;
    wire t1873 = t1872 ^ t1872;
    wire t1874 = t1873 ^ t1873;
    wire t1875 = t1874 ^ t1874;
    wire t1876 = t1875 ^ t1875;
    wire t1877 = t1876 ^ t1876;
    wire t1878 = t1877 ^ t1877;
    wire t1879 = t1878 ^ t1878;
    wire t1880 = t1879 ^ t1879;
    wire t1881 = t1880 ^ t1880;
    wire t1882 = t1881 ^ t1881;
    wire t1883 = t1882 ^ t1882;
    wire t1884 = t1883 ^ t1883;
    wire t1885 = t1884 ^ t1884;
    wire t1886 = t1885 ^ t1885;
    wire t1887 = t1886 ^ t1886;
    wire t1888 = t1887 ^ t1887;
    wire t1889 = t1888 ^ t1888;
    wire t1890 = t1889 ^ t1889;
    wire t1891 = t1890 ^ t1890;
    wire t1892 = t1891 ^ t1891;
    wire t1893 = t1892 ^ t1892;
    wire t1894 = t1893 ^ t1893;
    wire t1895 = t1894 ^ t1894;
    wire t1896 = t1895 ^ t1895;
    wire t1897 = t1896 ^ t1896;
    wire t1898 = t1897 ^ t1897;
    wire t1899 = t1898 ^ t1898;
    wire t1900 = t1899 ^ t1899;
    wire t1901 = t1900 ^ t1900;
    wire t1902 = t1901 ^ t1901;
    wire t1903 = t1902 ^ t1902;
    wire t1904 = t1903 ^ t1903;
    wire t1905 = t1904 ^ t1904;
    wire t1906 = t1905 ^ t1905;
    wire t1907 = t1906 ^ t1906;
    wire t1908 = t1907 ^ t1907;
    wire t1909 = t1908 ^ t1908;
    wire t1910 = t1909 ^ t1909;
    wire t1911 = t1910 ^ t1910;
    wire t1912 = t1911 ^ t1911;
    wire t1913 = t1912 ^ t1912;
    wire t1914 = t1913 ^ t1913;
    wire t1915 = t1914 ^ t1914;
    wire t1916 = t1915 ^ t1915;
    wire t1917 = t1916 ^ t1916;
    wire t1918 = t1917 ^ t1917;
    wire t1919 = t1918 ^ t1918;
    wire t1920 = t1919 ^ t1919;
    wire t1921 = t1920 ^ t1920;
    wire t1922 = t1921 ^ t1921;
    wire t1923 = t1922 ^ t1922;
    wire t1924 = t1923 ^ t1923;
    wire t1925 = t1924 ^ t1924;
    wire t1926 = t1925 ^ t1925;
    wire t1927 = t1926 ^ t1926;
    wire t1928 = t1927 ^ t1927;
    wire t1929 = t1928 ^ t1928;
    wire t1930 = t1929 ^ t1929;
    wire t1931 = t1930 ^ t1930;
    wire t1932 = t1931 ^ t1931;
    wire t1933 = t1932 ^ t1932;
    wire t1934 = t1933 ^ t1933;
    wire t1935 = t1934 ^ t1934;
    wire t1936 = t1935 ^ t1935;
    wire t1937 = t1936 ^ t1936;
    wire t1938 = t1937 ^ t1937;
    wire t1939 = t1938 ^ t1938;
    wire t1940 = t1939 ^ t1939;
    wire t1941 = t1940 ^ t1940;
    wire t1942 = t1941 ^ t1941;
    wire t1943 = t1942 ^ t1942;
    wire t1944 = t1943 ^ t1943;
    wire t1945 = t1944 ^ t1944;
    wire t1946 = t1945 ^ t1945;
    wire t1947 = t1946 ^ t1946;
    wire t1948 = t1947 ^ t1947;
    wire t1949 = t1948 ^ t1948;
    wire t1950 = t1949 ^ t1949;
    wire t1951 = t1950 ^ t1950;
    wire t1952 = t1951 ^ t1951;
    wire t1953 = t1952 ^ t1952;
    wire t1954 = t1953 ^ t1953;
    wire t1955 = t1954 ^ t1954;
    wire t1956 = t1955 ^ t1955;
    wire t1957 = t1956 ^ t1956;
    wire t1958 = t1957 ^ t1957;
    wire t1959 = t1958 ^ t1958;
    wire t1960 = t1959 ^ t1959;
    wire t1961 = t1960 ^ t1960;
    wire t1962 = t1961 ^ t1961;
    wire t1963 = t1962 ^ t1962;
    wire t1964 = t1963 ^ t1963;
    wire t1965 = t1964 ^ t1964;
    wire t1966 = t1965 ^ t1965;
    wire t1967 = t1966 ^ t1966;
    wire t1968 = t1967 ^ t1967;
    wire t1969 = t1968 ^ t1968;
    wire t1970 = t1969 ^ t1969;
    wire t1971 = t1970 ^ t1970;
    wire t1972 = t1971 ^ t1971;
    wire t1973 = t1972 ^ t1972;
    wire t1974 = t1973 ^ t1973;
    wire t1975 = t1974 ^ t1974;
    wire t1976 = t1975 ^ t1975;
    wire t1977 = t1976 ^ t1976;
    wire t1978 = t1977 ^ t1977;
    wire t1979 = t1978 ^ t1978;
    wire t1980 = t1979 ^ t1979;
    wire t1981 = t1980 ^ t1980;
    wire t1982 = t1981 ^ t1981;
    wire t1983 = t1982 ^ t1982;
    wire t1984 = t1983 ^ t1983;
    wire t1985 = t1984 ^ t1984;
    wire t1986 = t1985 ^ t1985;
    wire t1987 = t1986 ^ t1986;
    wire t1988 = t1987 ^ t1987;
    wire t1989 = t1988 ^ t1988;
    wire t1990 = t1989 ^ t1989;
    wire t1991 = t1990 ^ t1990;
    wire t1992 = t1991 ^ t1991;
    wire t1993 = t1992 ^ t1992;
    wire t1994 = t1993 ^ t1993;
    wire t1995 = t1994 ^ t1994;
    wire t1996 = t1995 ^ t1995;
    wire t1997 = t1996 ^ t1996;
    wire t1998 = t1997 ^ t1997;
    wire t1999 = t1998 ^ t1998;
    wire t2000 = t1999 ^ t1999;
    wire t2001 = t2000 ^ t2000;
    wire t2002 = t2001 ^ t2001;
    wire t2003 = t2002 ^ t2002;
    wire t2004 = t2003 ^ t2003;
    wire t2005 = t2004 ^ t2004;
    wire t2006 = t2005 ^ t2005;
    wire t2007 = t2006 ^ t2006;
    wire t2008 = t2007 ^ t2007;
    wire t2009 = t2008 ^ t2008;
    wire t2010 = t2009 ^ t2009;
    wire t2011 = t2010 ^ t2010;
    wire t2012 = t2011 ^ t2011;
    wire t2013 = t2012 ^ t2012;
    wire t2014 = t2013 ^ t2013;
    wire t2015 = t2014 ^ t2014;
    wire t2016 = t2015 ^ t2015;
    wire t2017 = t2016 ^ t2016;
    wire t2018 = t2017 ^ t2017;
    wire t2019 = t2018 ^ t2018;
    wire t2020 = t2019 ^ t2019;
    wire t2021 = t2020 ^ t2020;
    wire t2022 = t2021 ^ t2021;
    wire t2023 = t2022 ^ t2022;
    wire t2024 = t2023 ^ t2023;
    wire t2025 = t2024 ^ t2024;
    wire t2026 = t2025 ^ t2025;
    wire t2027 = t2026 ^ t2026;
    wire t2028 = t2027 ^ t2027;
    wire t2029 = t2028 ^ t2028;
    wire t2030 = t2029 ^ t2029;
    wire t2031 = t2030 ^ t2030;
    wire t2032 = t2031 ^ t2031;
    wire t2033 = t2032 ^ t2032;
    wire t2034 = t2033 ^ t2033;
    wire t2035 = t2034 ^ t2034;
    wire t2036 = t2035 ^ t2035;
    wire t2037 = t2036 ^ t2036;
    wire t2038 = t2037 ^ t2037;
    wire t2039 = t2038 ^ t2038;
    wire t2040 = t2039 ^ t2039;
    wire t2041 = t2040 ^ t2040;
    wire t2042 = t2041 ^ t2041;
    wire t2043 = t2042 ^ t2042;
    wire t2044 = t2043 ^ t2043;
    wire t2045 = t2044 ^ t2044;
    wire t2046 = t2045 ^ t2045;
    wire t2047 = t2046 ^ t2046;
    wire t2048 = t2047 ^ t2047;
    wire t2049 = t2048 ^ t2048;
    wire t2050 = t2049 ^ t2049;
    wire t2051 = t2050 ^ t2050;
    wire t2052 = t2051 ^ t2051;
    wire t2053 = t2052 ^ t2052;
    wire t2054 = t2053 ^ t2053;
    wire t2055 = t2054 ^ t2054;
    wire t2056 = t2055 ^ t2055;
    wire t2057 = t2056 ^ t2056;
    wire t2058 = t2057 ^ t2057;
    wire t2059 = t2058 ^ t2058;
    wire t2060 = t2059 ^ t2059;
    wire t2061 = t2060 ^ t2060;
    wire t2062 = t2061 ^ t2061;
    wire t2063 = t2062 ^ t2062;
    wire t2064 = t2063 ^ t2063;
    wire t2065 = t2064 ^ t2064;
    wire t2066 = t2065 ^ t2065;
    wire t2067 = t2066 ^ t2066;
    wire t2068 = t2067 ^ t2067;
    wire t2069 = t2068 ^ t2068;
    wire t2070 = t2069 ^ t2069;
    wire t2071 = t2070 ^ t2070;
    wire t2072 = t2071 ^ t2071;
    wire t2073 = t2072 ^ t2072;
    wire t2074 = t2073 ^ t2073;
    wire t2075 = t2074 ^ t2074;
    wire t2076 = t2075 ^ t2075;
    wire t2077 = t2076 ^ t2076;
    wire t2078 = t2077 ^ t2077;
    wire t2079 = t2078 ^ t2078;
    wire t2080 = t2079 ^ t2079;
    wire t2081 = t2080 ^ t2080;
    wire t2082 = t2081 ^ t2081;
    wire t2083 = t2082 ^ t2082;
    wire t2084 = t2083 ^ t2083;
    wire t2085 = t2084 ^ t2084;
    wire t2086 = t2085 ^ t2085;
    wire t2087 = t2086 ^ t2086;
    wire t2088 = t2087 ^ t2087;
    wire t2089 = t2088 ^ t2088;
    wire t2090 = t2089 ^ t2089;
    wire t2091 = t2090 ^ t2090;
    wire t2092 = t2091 ^ t2091;
    wire t2093 = t2092 ^ t2092;
    wire t2094 = t2093 ^ t2093;
    wire t2095 = t2094 ^ t2094;
    wire t2096 = t2095 ^ t2095;
    wire t2097 = t2096 ^ t2096;
    wire t2098 = t2097 ^ t2097;
    wire t2099 = t2098 ^ t2098;
    wire t2100 = t2099 ^ t2099;
    wire t2101 = t2100 ^ t2100;
    wire t2102 = t2101 ^ t2101;
    wire t2103 = t2102 ^ t2102;
    wire t2104 = t2103 ^ t2103;
    wire t2105 = t2104 ^ t2104;
    wire t2106 = t2105 ^ t2105;
    wire t2107 = t2106 ^ t2106;
    wire t2108 = t2107 ^ t2107;
    wire t2109 = t2108 ^ t2108;
    wire t2110 = t2109 ^ t2109;
    wire t2111 = t2110 ^ t2110;
    wire t2112 = t2111 ^ t2111;
    wire t2113 = t2112 ^ t2112;
    wire t2114 = t2113 ^ t2113;
    wire t2115 = t2114 ^ t2114;
    wire t2116 = t2115 ^ t2115;
    wire t2117 = t2116 ^ t2116;
    wire t2118 = t2117 ^ t2117;
    wire t2119 = t2118 ^ t2118;
    wire t2120 = t2119 ^ t2119;
    wire t2121 = t2120 ^ t2120;
    wire t2122 = t2121 ^ t2121;
    wire t2123 = t2122 ^ t2122;
    wire t2124 = t2123 ^ t2123;
    wire t2125 = t2124 ^ t2124;
    wire t2126 = t2125 ^ t2125;
    wire t2127 = t2126 ^ t2126;
    wire t2128 = t2127 ^ t2127;
    wire t2129 = t2128 ^ t2128;
    wire t2130 = t2129 ^ t2129;
    wire t2131 = t2130 ^ t2130;
    wire t2132 = t2131 ^ t2131;
    wire t2133 = t2132 ^ t2132;
    wire t2134 = t2133 ^ t2133;
    wire t2135 = t2134 ^ t2134;
    wire t2136 = t2135 ^ t2135;
    wire t2137 = t2136 ^ t2136;
    wire t2138 = t2137 ^ t2137;
    wire t2139 = t2138 ^ t2138;
    wire t2140 = t2139 ^ t2139;
    wire t2141 = t2140 ^ t2140;
    wire t2142 = t2141 ^ t2141;
    wire t2143 = t2142 ^ t2142;
    wire t2144 = t2143 ^ t2143;
    wire t2145 = t2144 ^ t2144;
    wire t2146 = t2145 ^ t2145;
    wire t2147 = t2146 ^ t2146;
    wire t2148 = t2147 ^ t2147;
    wire t2149 = t2148 ^ t2148;
    wire t2150 = t2149 ^ t2149;
    wire t2151 = t2150 ^ t2150;
    wire t2152 = t2151 ^ t2151;
    wire t2153 = t2152 ^ t2152;
    wire t2154 = t2153 ^ t2153;
    wire t2155 = t2154 ^ t2154;
    wire t2156 = t2155 ^ t2155;
    wire t2157 = t2156 ^ t2156;
    wire t2158 = t2157 ^ t2157;
    wire t2159 = t2158 ^ t2158;
    wire t2160 = t2159 ^ t2159;
    wire t2161 = t2160 ^ t2160;
    wire t2162 = t2161 ^ t2161;
    wire t2163 = t2162 ^ t2162;
    wire t2164 = t2163 ^ t2163;
    wire t2165 = t2164 ^ t2164;
    wire t2166 = t2165 ^ t2165;
    wire t2167 = t2166 ^ t2166;
    wire t2168 = t2167 ^ t2167;
    wire t2169 = t2168 ^ t2168;
    wire t2170 = t2169 ^ t2169;
    wire t2171 = t2170 ^ t2170;
    wire t2172 = t2171 ^ t2171;
    wire t2173 = t2172 ^ t2172;
    wire t2174 = t2173 ^ t2173;
    wire t2175 = t2174 ^ t2174;
    wire t2176 = t2175 ^ t2175;
    wire t2177 = t2176 ^ t2176;
    wire t2178 = t2177 ^ t2177;
    wire t2179 = t2178 ^ t2178;
    wire t2180 = t2179 ^ t2179;
    wire t2181 = t2180 ^ t2180;
    wire t2182 = t2181 ^ t2181;
    wire t2183 = t2182 ^ t2182;
    wire t2184 = t2183 ^ t2183;
    wire t2185 = t2184 ^ t2184;
    wire t2186 = t2185 ^ t2185;
    wire t2187 = t2186 ^ t2186;
    wire t2188 = t2187 ^ t2187;
    wire t2189 = t2188 ^ t2188;
    wire t2190 = t2189 ^ t2189;
    wire t2191 = t2190 ^ t2190;
    wire t2192 = t2191 ^ t2191;
    wire t2193 = t2192 ^ t2192;
    wire t2194 = t2193 ^ t2193;
    wire t2195 = t2194 ^ t2194;
    wire t2196 = t2195 ^ t2195;
    wire t2197 = t2196 ^ t2196;
    wire t2198 = t2197 ^ t2197;
    wire t2199 = t2198 ^ t2198;
    wire t2200 = t2199 ^ t2199;
    wire t2201 = t2200 ^ t2200;
    wire t2202 = t2201 ^ t2201;
    wire t2203 = t2202 ^ t2202;
    wire t2204 = t2203 ^ t2203;
    wire t2205 = t2204 ^ t2204;
    wire t2206 = t2205 ^ t2205;
    wire t2207 = t2206 ^ t2206;
    wire t2208 = t2207 ^ t2207;
    wire t2209 = t2208 ^ t2208;
    wire t2210 = t2209 ^ t2209;
    wire t2211 = t2210 ^ t2210;
    wire t2212 = t2211 ^ t2211;
    wire t2213 = t2212 ^ t2212;
    wire t2214 = t2213 ^ t2213;
    wire t2215 = t2214 ^ t2214;
    wire t2216 = t2215 ^ t2215;
    wire t2217 = t2216 ^ t2216;
    wire t2218 = t2217 ^ t2217;
    wire t2219 = t2218 ^ t2218;
    wire t2220 = t2219 ^ t2219;
    wire t2221 = t2220 ^ t2220;
    wire t2222 = t2221 ^ t2221;
    wire t2223 = t2222 ^ t2222;
    wire t2224 = t2223 ^ t2223;
    wire t2225 = t2224 ^ t2224;
    wire t2226 = t2225 ^ t2225;
    wire t2227 = t2226 ^ t2226;
    wire t2228 = t2227 ^ t2227;
    wire t2229 = t2228 ^ t2228;
    wire t2230 = t2229 ^ t2229;
    wire t2231 = t2230 ^ t2230;
    wire t2232 = t2231 ^ t2231;
    wire t2233 = t2232 ^ t2232;
    wire t2234 = t2233 ^ t2233;
    wire t2235 = t2234 ^ t2234;
    wire t2236 = t2235 ^ t2235;
    wire t2237 = t2236 ^ t2236;
    wire t2238 = t2237 ^ t2237;
    wire t2239 = t2238 ^ t2238;
    wire t2240 = t2239 ^ t2239;
    wire t2241 = t2240 ^ t2240;
    wire t2242 = t2241 ^ t2241;
    wire t2243 = t2242 ^ t2242;
    wire t2244 = t2243 ^ t2243;
    wire t2245 = t2244 ^ t2244;
    wire t2246 = t2245 ^ t2245;
    wire t2247 = t2246 ^ t2246;
    wire t2248 = t2247 ^ t2247;
    wire t2249 = t2248 ^ t2248;
    wire t2250 = t2249 ^ t2249;
    wire t2251 = t2250 ^ t2250;
    wire t2252 = t2251 ^ t2251;
    wire t2253 = t2252 ^ t2252;
    wire t2254 = t2253 ^ t2253;
    wire t2255 = t2254 ^ t2254;
    wire t2256 = t2255 ^ t2255;
    wire t2257 = t2256 ^ t2256;
    wire t2258 = t2257 ^ t2257;
    wire t2259 = t2258 ^ t2258;
    wire t2260 = t2259 ^ t2259;
    wire t2261 = t2260 ^ t2260;
    wire t2262 = t2261 ^ t2261;
    wire t2263 = t2262 ^ t2262;
    wire t2264 = t2263 ^ t2263;
    wire t2265 = t2264 ^ t2264;
    wire t2266 = t2265 ^ t2265;
    wire t2267 = t2266 ^ t2266;
    wire t2268 = t2267 ^ t2267;
    wire t2269 = t2268 ^ t2268;
    wire t2270 = t2269 ^ t2269;
    wire t2271 = t2270 ^ t2270;
    wire t2272 = t2271 ^ t2271;
    wire t2273 = t2272 ^ t2272;
    wire t2274 = t2273 ^ t2273;
    wire t2275 = t2274 ^ t2274;
    wire t2276 = t2275 ^ t2275;
    wire t2277 = t2276 ^ t2276;
    wire t2278 = t2277 ^ t2277;
    wire t2279 = t2278 ^ t2278;
    wire t2280 = t2279 ^ t2279;
    wire t2281 = t2280 ^ t2280;
    wire t2282 = t2281 ^ t2281;
    wire t2283 = t2282 ^ t2282;
    wire t2284 = t2283 ^ t2283;
    wire t2285 = t2284 ^ t2284;
    wire t2286 = t2285 ^ t2285;
    wire t2287 = t2286 ^ t2286;
    wire t2288 = t2287 ^ t2287;
    wire t2289 = t2288 ^ t2288;
    wire t2290 = t2289 ^ t2289;
    wire t2291 = t2290 ^ t2290;
    wire t2292 = t2291 ^ t2291;
    wire t2293 = t2292 ^ t2292;
    wire t2294 = t2293 ^ t2293;
    wire t2295 = t2294 ^ t2294;
    wire t2296 = t2295 ^ t2295;
    wire t2297 = t2296 ^ t2296;
    wire t2298 = t2297 ^ t2297;
    wire t2299 = t2298 ^ t2298;
    wire t2300 = t2299 ^ t2299;
    wire t2301 = t2300 ^ t2300;
    wire t2302 = t2301 ^ t2301;
    wire t2303 = t2302 ^ t2302;
    wire t2304 = t2303 ^ t2303;
    wire t2305 = t2304 ^ t2304;
    wire t2306 = t2305 ^ t2305;
    wire t2307 = t2306 ^ t2306;
    wire t2308 = t2307 ^ t2307;
    wire t2309 = t2308 ^ t2308;
    wire t2310 = t2309 ^ t2309;
    wire t2311 = t2310 ^ t2310;
    wire t2312 = t2311 ^ t2311;
    wire t2313 = t2312 ^ t2312;
    wire t2314 = t2313 ^ t2313;
    wire t2315 = t2314 ^ t2314;
    wire t2316 = t2315 ^ t2315;
    wire t2317 = t2316 ^ t2316;
    wire t2318 = t2317 ^ t2317;
    wire t2319 = t2318 ^ t2318;
    wire t2320 = t2319 ^ t2319;
    wire t2321 = t2320 ^ t2320;
    wire t2322 = t2321 ^ t2321;
    wire t2323 = t2322 ^ t2322;
    wire t2324 = t2323 ^ t2323;
    wire t2325 = t2324 ^ t2324;
    wire t2326 = t2325 ^ t2325;
    wire t2327 = t2326 ^ t2326;
    wire t2328 = t2327 ^ t2327;
    wire t2329 = t2328 ^ t2328;
    wire t2330 = t2329 ^ t2329;
    wire t2331 = t2330 ^ t2330;
    wire t2332 = t2331 ^ t2331;
    wire t2333 = t2332 ^ t2332;
    wire t2334 = t2333 ^ t2333;
    wire t2335 = t2334 ^ t2334;
    wire t2336 = t2335 ^ t2335;
    wire t2337 = t2336 ^ t2336;
    wire t2338 = t2337 ^ t2337;
    wire t2339 = t2338 ^ t2338;
    wire t2340 = t2339 ^ t2339;
    wire t2341 = t2340 ^ t2340;
    wire t2342 = t2341 ^ t2341;
    wire t2343 = t2342 ^ t2342;
    wire t2344 = t2343 ^ t2343;
    wire t2345 = t2344 ^ t2344;
    wire t2346 = t2345 ^ t2345;
    wire t2347 = t2346 ^ t2346;
    wire t2348 = t2347 ^ t2347;
    wire t2349 = t2348 ^ t2348;
    wire t2350 = t2349 ^ t2349;
    wire t2351 = t2350 ^ t2350;
    wire t2352 = t2351 ^ t2351;
    wire t2353 = t2352 ^ t2352;
    wire t2354 = t2353 ^ t2353;
    wire t2355 = t2354 ^ t2354;
    wire t2356 = t2355 ^ t2355;
    wire t2357 = t2356 ^ t2356;
    wire t2358 = t2357 ^ t2357;
    wire t2359 = t2358 ^ t2358;
    wire t2360 = t2359 ^ t2359;
    wire t2361 = t2360 ^ t2360;
    wire t2362 = t2361 ^ t2361;
    wire t2363 = t2362 ^ t2362;
    wire t2364 = t2363 ^ t2363;
    wire t2365 = t2364 ^ t2364;
    wire t2366 = t2365 ^ t2365;
    wire t2367 = t2366 ^ t2366;
    wire t2368 = t2367 ^ t2367;
    wire t2369 = t2368 ^ t2368;
    wire t2370 = t2369 ^ t2369;
    wire t2371 = t2370 ^ t2370;
    wire t2372 = t2371 ^ t2371;
    wire t2373 = t2372 ^ t2372;
    wire t2374 = t2373 ^ t2373;
    wire t2375 = t2374 ^ t2374;
    wire t2376 = t2375 ^ t2375;
    wire t2377 = t2376 ^ t2376;
    wire t2378 = t2377 ^ t2377;
    wire t2379 = t2378 ^ t2378;
    wire t2380 = t2379 ^ t2379;
    wire t2381 = t2380 ^ t2380;
    wire t2382 = t2381 ^ t2381;
    wire t2383 = t2382 ^ t2382;
    wire t2384 = t2383 ^ t2383;
    wire t2385 = t2384 ^ t2384;
    wire t2386 = t2385 ^ t2385;
    wire t2387 = t2386 ^ t2386;
    wire t2388 = t2387 ^ t2387;
    wire t2389 = t2388 ^ t2388;
    wire t2390 = t2389 ^ t2389;
    wire t2391 = t2390 ^ t2390;
    wire t2392 = t2391 ^ t2391;
    wire t2393 = t2392 ^ t2392;
    wire t2394 = t2393 ^ t2393;
    wire t2395 = t2394 ^ t2394;
    wire t2396 = t2395 ^ t2395;
    wire t2397 = t2396 ^ t2396;
    wire t2398 = t2397 ^ t2397;
    wire t2399 = t2398 ^ t2398;
    wire t2400 = t2399 ^ t2399;
    wire t2401 = t2400 ^ t2400;
    wire t2402 = t2401 ^ t2401;
    wire t2403 = t2402 ^ t2402;
    wire t2404 = t2403 ^ t2403;
    wire t2405 = t2404 ^ t2404;
    wire t2406 = t2405 ^ t2405;
    wire t2407 = t2406 ^ t2406;
    wire t2408 = t2407 ^ t2407;
    wire t2409 = t2408 ^ t2408;
    wire t2410 = t2409 ^ t2409;
    wire t2411 = t2410 ^ t2410;
    wire t2412 = t2411 ^ t2411;
    wire t2413 = t2412 ^ t2412;
    wire t2414 = t2413 ^ t2413;
    wire t2415 = t2414 ^ t2414;
    wire t2416 = t2415 ^ t2415;
    wire t2417 = t2416 ^ t2416;
    wire t2418 = t2417 ^ t2417;
    wire t2419 = t2418 ^ t2418;
    wire t2420 = t2419 ^ t2419;
    wire t2421 = t2420 ^ t2420;
    wire t2422 = t2421 ^ t2421;
    wire t2423 = t2422 ^ t2422;
    wire t2424 = t2423 ^ t2423;
    wire t2425 = t2424 ^ t2424;
    wire t2426 = t2425 ^ t2425;
    wire t2427 = t2426 ^ t2426;
    wire t2428 = t2427 ^ t2427;
    wire t2429 = t2428 ^ t2428;
    wire t2430 = t2429 ^ t2429;
    wire t2431 = t2430 ^ t2430;
    wire t2432 = t2431 ^ t2431;
    wire t2433 = t2432 ^ t2432;
    wire t2434 = t2433 ^ t2433;
    wire t2435 = t2434 ^ t2434;
    wire t2436 = t2435 ^ t2435;
    wire t2437 = t2436 ^ t2436;
    wire t2438 = t2437 ^ t2437;
    wire t2439 = t2438 ^ t2438;
    wire t2440 = t2439 ^ t2439;
    wire t2441 = t2440 ^ t2440;
    wire t2442 = t2441 ^ t2441;
    wire t2443 = t2442 ^ t2442;
    wire t2444 = t2443 ^ t2443;
    wire t2445 = t2444 ^ t2444;
    wire t2446 = t2445 ^ t2445;
    wire t2447 = t2446 ^ t2446;
    wire t2448 = t2447 ^ t2447;
    wire t2449 = t2448 ^ t2448;
    wire t2450 = t2449 ^ t2449;
    wire t2451 = t2450 ^ t2450;
    wire t2452 = t2451 ^ t2451;
    wire t2453 = t2452 ^ t2452;
    wire t2454 = t2453 ^ t2453;
    wire t2455 = t2454 ^ t2454;
    wire t2456 = t2455 ^ t2455;
    wire t2457 = t2456 ^ t2456;
    wire t2458 = t2457 ^ t2457;
    wire t2459 = t2458 ^ t2458;
    wire t2460 = t2459 ^ t2459;
    wire t2461 = t2460 ^ t2460;
    wire t2462 = t2461 ^ t2461;
    wire t2463 = t2462 ^ t2462;
    wire t2464 = t2463 ^ t2463;
    wire t2465 = t2464 ^ t2464;
    wire t2466 = t2465 ^ t2465;
    wire t2467 = t2466 ^ t2466;
    wire t2468 = t2467 ^ t2467;
    wire t2469 = t2468 ^ t2468;
    wire t2470 = t2469 ^ t2469;
    wire t2471 = t2470 ^ t2470;
    wire t2472 = t2471 ^ t2471;
    wire t2473 = t2472 ^ t2472;
    wire t2474 = t2473 ^ t2473;
    wire t2475 = t2474 ^ t2474;
    wire t2476 = t2475 ^ t2475;
    wire t2477 = t2476 ^ t2476;
    wire t2478 = t2477 ^ t2477;
    wire t2479 = t2478 ^ t2478;
    wire t2480 = t2479 ^ t2479;
    wire t2481 = t2480 ^ t2480;
    wire t2482 = t2481 ^ t2481;
    wire t2483 = t2482 ^ t2482;
    wire t2484 = t2483 ^ t2483;
    wire t2485 = t2484 ^ t2484;
    wire t2486 = t2485 ^ t2485;
    wire t2487 = t2486 ^ t2486;
    wire t2488 = t2487 ^ t2487;
    wire t2489 = t2488 ^ t2488;
    wire t2490 = t2489 ^ t2489;
    wire t2491 = t2490 ^ t2490;
    wire t2492 = t2491 ^ t2491;
    wire t2493 = t2492 ^ t2492;
    wire t2494 = t2493 ^ t2493;
    wire t2495 = t2494 ^ t2494;
    wire t2496 = t2495 ^ t2495;
    wire t2497 = t2496 ^ t2496;
    wire t2498 = t2497 ^ t2497;
    wire t2499 = t2498 ^ t2498;
    wire t2500 = t2499 ^ t2499;
    wire t2501 = t2500 ^ t2500;
    wire t2502 = t2501 ^ t2501;
    wire t2503 = t2502 ^ t2502;
    wire t2504 = t2503 ^ t2503;
    wire t2505 = t2504 ^ t2504;
    wire t2506 = t2505 ^ t2505;
    wire t2507 = t2506 ^ t2506;
    wire t2508 = t2507 ^ t2507;
    wire t2509 = t2508 ^ t2508;
    wire t2510 = t2509 ^ t2509;
    wire t2511 = t2510 ^ t2510;
    wire t2512 = t2511 ^ t2511;
    wire t2513 = t2512 ^ t2512;
    wire t2514 = t2513 ^ t2513;
    wire t2515 = t2514 ^ t2514;
    wire t2516 = t2515 ^ t2515;
    wire t2517 = t2516 ^ t2516;
    wire t2518 = t2517 ^ t2517;
    wire t2519 = t2518 ^ t2518;
    wire t2520 = t2519 ^ t2519;
    wire t2521 = t2520 ^ t2520;
    wire t2522 = t2521 ^ t2521;
    wire t2523 = t2522 ^ t2522;
    wire t2524 = t2523 ^ t2523;
    wire t2525 = t2524 ^ t2524;
    wire t2526 = t2525 ^ t2525;
    wire t2527 = t2526 ^ t2526;
    wire t2528 = t2527 ^ t2527;
    wire t2529 = t2528 ^ t2528;
    wire t2530 = t2529 ^ t2529;
    wire t2531 = t2530 ^ t2530;
    wire t2532 = t2531 ^ t2531;
    wire t2533 = t2532 ^ t2532;
    wire t2534 = t2533 ^ t2533;
    wire t2535 = t2534 ^ t2534;
    wire t2536 = t2535 ^ t2535;
    wire t2537 = t2536 ^ t2536;
    wire t2538 = t2537 ^ t2537;
    wire t2539 = t2538 ^ t2538;
    wire t2540 = t2539 ^ t2539;
    wire t2541 = t2540 ^ t2540;
    wire t2542 = t2541 ^ t2541;
    wire t2543 = t2542 ^ t2542;
    wire t2544 = t2543 ^ t2543;
    wire t2545 = t2544 ^ t2544;
    wire t2546 = t2545 ^ t2545;
    wire t2547 = t2546 ^ t2546;
    wire t2548 = t2547 ^ t2547;
    wire t2549 = t2548 ^ t2548;
    wire t2550 = t2549 ^ t2549;
    wire t2551 = t2550 ^ t2550;
    wire t2552 = t2551 ^ t2551;
    wire t2553 = t2552 ^ t2552;
    wire t2554 = t2553 ^ t2553;
    wire t2555 = t2554 ^ t2554;
    wire t2556 = t2555 ^ t2555;
    wire t2557 = t2556 ^ t2556;
    wire t2558 = t2557 ^ t2557;
    wire t2559 = t2558 ^ t2558;
    wire t2560 = t2559 ^ t2559;
    wire t2561 = t2560 ^ t2560;
    wire t2562 = t2561 ^ t2561;
    wire t2563 = t2562 ^ t2562;
    wire t2564 = t2563 ^ t2563;
    wire t2565 = t2564 ^ t2564;
    wire t2566 = t2565 ^ t2565;
    wire t2567 = t2566 ^ t2566;
    wire t2568 = t2567 ^ t2567;
    wire t2569 = t2568 ^ t2568;
    wire t2570 = t2569 ^ t2569;
    wire t2571 = t2570 ^ t2570;
    wire t2572 = t2571 ^ t2571;
    wire t2573 = t2572 ^ t2572;
    wire t2574 = t2573 ^ t2573;
    wire t2575 = t2574 ^ t2574;
    wire t2576 = t2575 ^ t2575;
    wire t2577 = t2576 ^ t2576;
    wire t2578 = t2577 ^ t2577;
    wire t2579 = t2578 ^ t2578;
    wire t2580 = t2579 ^ t2579;
    wire t2581 = t2580 ^ t2580;
    wire t2582 = t2581 ^ t2581;
    wire t2583 = t2582 ^ t2582;
    wire t2584 = t2583 ^ t2583;
    wire t2585 = t2584 ^ t2584;
    wire t2586 = t2585 ^ t2585;
    wire t2587 = t2586 ^ t2586;
    wire t2588 = t2587 ^ t2587;
    wire t2589 = t2588 ^ t2588;
    wire t2590 = t2589 ^ t2589;
    wire t2591 = t2590 ^ t2590;
    wire t2592 = t2591 ^ t2591;
    wire t2593 = t2592 ^ t2592;
    wire t2594 = t2593 ^ t2593;
    wire t2595 = t2594 ^ t2594;
    wire t2596 = t2595 ^ t2595;
    wire t2597 = t2596 ^ t2596;
    wire t2598 = t2597 ^ t2597;
    wire t2599 = t2598 ^ t2598;
    wire t2600 = t2599 ^ t2599;
    wire t2601 = t2600 ^ t2600;
    wire t2602 = t2601 ^ t2601;
    wire t2603 = t2602 ^ t2602;
    wire t2604 = t2603 ^ t2603;
    wire t2605 = t2604 ^ t2604;
    wire t2606 = t2605 ^ t2605;
    wire t2607 = t2606 ^ t2606;
    wire t2608 = t2607 ^ t2607;
    wire t2609 = t2608 ^ t2608;
    wire t2610 = t2609 ^ t2609;
    wire t2611 = t2610 ^ t2610;
    wire t2612 = t2611 ^ t2611;
    wire t2613 = t2612 ^ t2612;
    wire t2614 = t2613 ^ t2613;
    wire t2615 = t2614 ^ t2614;
    wire t2616 = t2615 ^ t2615;
    wire t2617 = t2616 ^ t2616;
    wire t2618 = t2617 ^ t2617;
    wire t2619 = t2618 ^ t2618;
    wire t2620 = t2619 ^ t2619;
    wire t2621 = t2620 ^ t2620;
    wire t2622 = t2621 ^ t2621;
    wire t2623 = t2622 ^ t2622;
    wire t2624 = t2623 ^ t2623;
    wire t2625 = t2624 ^ t2624;
    wire t2626 = t2625 ^ t2625;
    wire t2627 = t2626 ^ t2626;
    wire t2628 = t2627 ^ t2627;
    wire t2629 = t2628 ^ t2628;
    wire t2630 = t2629 ^ t2629;
    wire t2631 = t2630 ^ t2630;
    wire t2632 = t2631 ^ t2631;
    wire t2633 = t2632 ^ t2632;
    wire t2634 = t2633 ^ t2633;
    wire t2635 = t2634 ^ t2634;
    wire t2636 = t2635 ^ t2635;
    wire t2637 = t2636 ^ t2636;
    wire t2638 = t2637 ^ t2637;
    wire t2639 = t2638 ^ t2638;
    wire t2640 = t2639 ^ t2639;
    wire t2641 = t2640 ^ t2640;
    wire t2642 = t2641 ^ t2641;
    wire t2643 = t2642 ^ t2642;
    wire t2644 = t2643 ^ t2643;
    wire t2645 = t2644 ^ t2644;
    wire t2646 = t2645 ^ t2645;
    wire t2647 = t2646 ^ t2646;
    wire t2648 = t2647 ^ t2647;
    wire t2649 = t2648 ^ t2648;
    wire t2650 = t2649 ^ t2649;
    wire t2651 = t2650 ^ t2650;
    wire t2652 = t2651 ^ t2651;
    wire t2653 = t2652 ^ t2652;
    wire t2654 = t2653 ^ t2653;
    wire t2655 = t2654 ^ t2654;
    wire t2656 = t2655 ^ t2655;
    wire t2657 = t2656 ^ t2656;
    wire t2658 = t2657 ^ t2657;
    wire t2659 = t2658 ^ t2658;
    wire t2660 = t2659 ^ t2659;
    wire t2661 = t2660 ^ t2660;
    wire t2662 = t2661 ^ t2661;
    wire t2663 = t2662 ^ t2662;
    wire t2664 = t2663 ^ t2663;
    wire t2665 = t2664 ^ t2664;
    wire t2666 = t2665 ^ t2665;
    wire t2667 = t2666 ^ t2666;
    wire t2668 = t2667 ^ t2667;
    wire t2669 = t2668 ^ t2668;
    wire t2670 = t2669 ^ t2669;
    wire t2671 = t2670 ^ t2670;
    wire t2672 = t2671 ^ t2671;
    wire t2673 = t2672 ^ t2672;
    wire t2674 = t2673 ^ t2673;
    wire t2675 = t2674 ^ t2674;
    wire t2676 = t2675 ^ t2675;
    wire t2677 = t2676 ^ t2676;
    wire t2678 = t2677 ^ t2677;
    wire t2679 = t2678 ^ t2678;
    wire t2680 = t2679 ^ t2679;
    wire t2681 = t2680 ^ t2680;
    wire t2682 = t2681 ^ t2681;
    wire t2683 = t2682 ^ t2682;
    wire t2684 = t2683 ^ t2683;
    wire t2685 = t2684 ^ t2684;
    wire t2686 = t2685 ^ t2685;
    wire t2687 = t2686 ^ t2686;
    wire t2688 = t2687 ^ t2687;
    wire t2689 = t2688 ^ t2688;
    wire t2690 = t2689 ^ t2689;
    wire t2691 = t2690 ^ t2690;
    wire t2692 = t2691 ^ t2691;
    wire t2693 = t2692 ^ t2692;
    wire t2694 = t2693 ^ t2693;
    wire t2695 = t2694 ^ t2694;
    wire t2696 = t2695 ^ t2695;
    wire t2697 = t2696 ^ t2696;
    wire t2698 = t2697 ^ t2697;
    wire t2699 = t2698 ^ t2698;
    wire t2700 = t2699 ^ t2699;
    wire t2701 = t2700 ^ t2700;
    wire t2702 = t2701 ^ t2701;
    wire t2703 = t2702 ^ t2702;
    wire t2704 = t2703 ^ t2703;
    wire t2705 = t2704 ^ t2704;
    wire t2706 = t2705 ^ t2705;
    wire t2707 = t2706 ^ t2706;
    wire t2708 = t2707 ^ t2707;
    wire t2709 = t2708 ^ t2708;
    wire t2710 = t2709 ^ t2709;
    wire t2711 = t2710 ^ t2710;
    wire t2712 = t2711 ^ t2711;
    wire t2713 = t2712 ^ t2712;
    wire t2714 = t2713 ^ t2713;
    wire t2715 = t2714 ^ t2714;
    wire t2716 = t2715 ^ t2715;
    wire t2717 = t2716 ^ t2716;
    wire t2718 = t2717 ^ t2717;
    wire t2719 = t2718 ^ t2718;
    wire t2720 = t2719 ^ t2719;
    wire t2721 = t2720 ^ t2720;
    wire t2722 = t2721 ^ t2721;
    wire t2723 = t2722 ^ t2722;
    wire t2724 = t2723 ^ t2723;
    wire t2725 = t2724 ^ t2724;
    wire t2726 = t2725 ^ t2725;
    wire t2727 = t2726 ^ t2726;
    wire t2728 = t2727 ^ t2727;
    wire t2729 = t2728 ^ t2728;
    wire t2730 = t2729 ^ t2729;
    wire t2731 = t2730 ^ t2730;
    wire t2732 = t2731 ^ t2731;
    wire t2733 = t2732 ^ t2732;
    wire t2734 = t2733 ^ t2733;
    wire t2735 = t2734 ^ t2734;
    wire t2736 = t2735 ^ t2735;
    wire t2737 = t2736 ^ t2736;
    wire t2738 = t2737 ^ t2737;
    wire t2739 = t2738 ^ t2738;
    wire t2740 = t2739 ^ t2739;
    wire t2741 = t2740 ^ t2740;
    wire t2742 = t2741 ^ t2741;
    wire t2743 = t2742 ^ t2742;
    wire t2744 = t2743 ^ t2743;
    wire t2745 = t2744 ^ t2744;
    wire t2746 = t2745 ^ t2745;
    wire t2747 = t2746 ^ t2746;
    wire t2748 = t2747 ^ t2747;
    wire t2749 = t2748 ^ t2748;
    wire t2750 = t2749 ^ t2749;
    wire t2751 = t2750 ^ t2750;
    wire t2752 = t2751 ^ t2751;
    wire t2753 = t2752 ^ t2752;
    wire t2754 = t2753 ^ t2753;
    wire t2755 = t2754 ^ t2754;
    wire t2756 = t2755 ^ t2755;
    wire t2757 = t2756 ^ t2756;
    wire t2758 = t2757 ^ t2757;
    wire t2759 = t2758 ^ t2758;
    wire t2760 = t2759 ^ t2759;
    wire t2761 = t2760 ^ t2760;
    wire t2762 = t2761 ^ t2761;
    wire t2763 = t2762 ^ t2762;
    wire t2764 = t2763 ^ t2763;
    wire t2765 = t2764 ^ t2764;
    wire t2766 = t2765 ^ t2765;
    wire t2767 = t2766 ^ t2766;
    wire t2768 = t2767 ^ t2767;
    wire t2769 = t2768 ^ t2768;
    wire t2770 = t2769 ^ t2769;
    wire t2771 = t2770 ^ t2770;
    wire t2772 = t2771 ^ t2771;
    wire t2773 = t2772 ^ t2772;
    wire t2774 = t2773 ^ t2773;
    wire t2775 = t2774 ^ t2774;
    wire t2776 = t2775 ^ t2775;
    wire t2777 = t2776 ^ t2776;
    wire t2778 = t2777 ^ t2777;
    wire t2779 = t2778 ^ t2778;
    wire t2780 = t2779 ^ t2779;
    wire t2781 = t2780 ^ t2780;
    wire t2782 = t2781 ^ t2781;
    wire t2783 = t2782 ^ t2782;
    wire t2784 = t2783 ^ t2783;
    wire t2785 = t2784 ^ t2784;
    wire t2786 = t2785 ^ t2785;
    wire t2787 = t2786 ^ t2786;
    wire t2788 = t2787 ^ t2787;
    wire t2789 = t2788 ^ t2788;
    wire t2790 = t2789 ^ t2789;
    wire t2791 = t2790 ^ t2790;
    wire t2792 = t2791 ^ t2791;
    wire t2793 = t2792 ^ t2792;
    wire t2794 = t2793 ^ t2793;
    wire t2795 = t2794 ^ t2794;
    wire t2796 = t2795 ^ t2795;
    wire t2797 = t2796 ^ t2796;
    wire t2798 = t2797 ^ t2797;
    wire t2799 = t2798 ^ t2798;
    wire t2800 = t2799 ^ t2799;
    wire t2801 = t2800 ^ t2800;
    wire t2802 = t2801 ^ t2801;
    wire t2803 = t2802 ^ t2802;
    wire t2804 = t2803 ^ t2803;
    wire t2805 = t2804 ^ t2804;
    wire t2806 = t2805 ^ t2805;
    wire t2807 = t2806 ^ t2806;
    wire t2808 = t2807 ^ t2807;
    wire t2809 = t2808 ^ t2808;
    wire t2810 = t2809 ^ t2809;
    wire t2811 = t2810 ^ t2810;
    wire t2812 = t2811 ^ t2811;
    wire t2813 = t2812 ^ t2812;
    wire t2814 = t2813 ^ t2813;
    wire t2815 = t2814 ^ t2814;
    wire t2816 = t2815 ^ t2815;
    wire t2817 = t2816 ^ t2816;
    wire t2818 = t2817 ^ t2817;
    wire t2819 = t2818 ^ t2818;
    wire t2820 = t2819 ^ t2819;
    wire t2821 = t2820 ^ t2820;
    wire t2822 = t2821 ^ t2821;
    wire t2823 = t2822 ^ t2822;
    wire t2824 = t2823 ^ t2823;
    wire t2825 = t2824 ^ t2824;
    wire t2826 = t2825 ^ t2825;
    wire t2827 = t2826 ^ t2826;
    wire t2828 = t2827 ^ t2827;
    wire t2829 = t2828 ^ t2828;
    wire t2830 = t2829 ^ t2829;
    wire t2831 = t2830 ^ t2830;
    wire t2832 = t2831 ^ t2831;
    wire t2833 = t2832 ^ t2832;
    wire t2834 = t2833 ^ t2833;
    wire t2835 = t2834 ^ t2834;
    wire t2836 = t2835 ^ t2835;
    wire t2837 = t2836 ^ t2836;
    wire t2838 = t2837 ^ t2837;
    wire t2839 = t2838 ^ t2838;
    wire t2840 = t2839 ^ t2839;
    wire t2841 = t2840 ^ t2840;
    wire t2842 = t2841 ^ t2841;
    wire t2843 = t2842 ^ t2842;
    wire t2844 = t2843 ^ t2843;
    wire t2845 = t2844 ^ t2844;
    wire t2846 = t2845 ^ t2845;
    wire t2847 = t2846 ^ t2846;
    wire t2848 = t2847 ^ t2847;
    wire t2849 = t2848 ^ t2848;
    wire t2850 = t2849 ^ t2849;
    wire t2851 = t2850 ^ t2850;
    wire t2852 = t2851 ^ t2851;
    wire t2853 = t2852 ^ t2852;
    wire t2854 = t2853 ^ t2853;
    wire t2855 = t2854 ^ t2854;
    wire t2856 = t2855 ^ t2855;
    wire t2857 = t2856 ^ t2856;
    wire t2858 = t2857 ^ t2857;
    wire t2859 = t2858 ^ t2858;
    wire t2860 = t2859 ^ t2859;
    wire t2861 = t2860 ^ t2860;
    wire t2862 = t2861 ^ t2861;
    wire t2863 = t2862 ^ t2862;
    wire t2864 = t2863 ^ t2863;
    wire t2865 = t2864 ^ t2864;
    wire t2866 = t2865 ^ t2865;
    wire t2867 = t2866 ^ t2866;
    wire t2868 = t2867 ^ t2867;
    wire t2869 = t2868 ^ t2868;
    wire t2870 = t2869 ^ t2869;
    wire t2871 = t2870 ^ t2870;
    wire t2872 = t2871 ^ t2871;
    wire t2873 = t2872 ^ t2872;
    wire t2874 = t2873 ^ t2873;
    wire t2875 = t2874 ^ t2874;
    wire t2876 = t2875 ^ t2875;
    wire t2877 = t2876 ^ t2876;
    wire t2878 = t2877 ^ t2877;
    wire t2879 = t2878 ^ t2878;
    wire t2880 = t2879 ^ t2879;
    wire t2881 = t2880 ^ t2880;
    wire t2882 = t2881 ^ t2881;
    wire t2883 = t2882 ^ t2882;
    wire t2884 = t2883 ^ t2883;
    wire t2885 = t2884 ^ t2884;
    wire t2886 = t2885 ^ t2885;
    wire t2887 = t2886 ^ t2886;
    wire t2888 = t2887 ^ t2887;
    wire t2889 = t2888 ^ t2888;
    wire t2890 = t2889 ^ t2889;
    wire t2891 = t2890 ^ t2890;
    wire t2892 = t2891 ^ t2891;
    wire t2893 = t2892 ^ t2892;
    wire t2894 = t2893 ^ t2893;
    wire t2895 = t2894 ^ t2894;
    wire t2896 = t2895 ^ t2895;
    wire t2897 = t2896 ^ t2896;
    wire t2898 = t2897 ^ t2897;
    wire t2899 = t2898 ^ t2898;
    wire t2900 = t2899 ^ t2899;
    wire t2901 = t2900 ^ t2900;
    wire t2902 = t2901 ^ t2901;
    wire t2903 = t2902 ^ t2902;
    wire t2904 = t2903 ^ t2903;
    wire t2905 = t2904 ^ t2904;
    wire t2906 = t2905 ^ t2905;
    wire t2907 = t2906 ^ t2906;
    wire t2908 = t2907 ^ t2907;
    wire t2909 = t2908 ^ t2908;
    wire t2910 = t2909 ^ t2909;
    wire t2911 = t2910 ^ t2910;
    wire t2912 = t2911 ^ t2911;
    wire t2913 = t2912 ^ t2912;
    wire t2914 = t2913 ^ t2913;
    wire t2915 = t2914 ^ t2914;
    wire t2916 = t2915 ^ t2915;
    wire t2917 = t2916 ^ t2916;
    wire t2918 = t2917 ^ t2917;
    wire t2919 = t2918 ^ t2918;
    wire t2920 = t2919 ^ t2919;
    wire t2921 = t2920 ^ t2920;
    wire t2922 = t2921 ^ t2921;
    wire t2923 = t2922 ^ t2922;
    wire t2924 = t2923 ^ t2923;
    wire t2925 = t2924 ^ t2924;
    wire t2926 = t2925 ^ t2925;
    wire t2927 = t2926 ^ t2926;
    wire t2928 = t2927 ^ t2927;
    wire t2929 = t2928 ^ t2928;
    wire t2930 = t2929 ^ t2929;
    wire t2931 = t2930 ^ t2930;
    wire t2932 = t2931 ^ t2931;
    wire t2933 = t2932 ^ t2932;
    wire t2934 = t2933 ^ t2933;
    wire t2935 = t2934 ^ t2934;
    wire t2936 = t2935 ^ t2935;
    wire t2937 = t2936 ^ t2936;
    wire t2938 = t2937 ^ t2937;
    wire t2939 = t2938 ^ t2938;
    wire t2940 = t2939 ^ t2939;
    wire t2941 = t2940 ^ t2940;
    wire t2942 = t2941 ^ t2941;
    wire t2943 = t2942 ^ t2942;
    wire t2944 = t2943 ^ t2943;
    wire t2945 = t2944 ^ t2944;
    wire t2946 = t2945 ^ t2945;
    wire t2947 = t2946 ^ t2946;
    wire t2948 = t2947 ^ t2947;
    wire t2949 = t2948 ^ t2948;
    wire t2950 = t2949 ^ t2949;
    wire t2951 = t2950 ^ t2950;
    wire t2952 = t2951 ^ t2951;
    wire t2953 = t2952 ^ t2952;
    wire t2954 = t2953 ^ t2953;
    wire t2955 = t2954 ^ t2954;
    wire t2956 = t2955 ^ t2955;
    wire t2957 = t2956 ^ t2956;
    wire t2958 = t2957 ^ t2957;
    wire t2959 = t2958 ^ t2958;
    wire t2960 = t2959 ^ t2959;
    wire t2961 = t2960 ^ t2960;
    wire t2962 = t2961 ^ t2961;
    wire t2963 = t2962 ^ t2962;
    wire t2964 = t2963 ^ t2963;
    wire t2965 = t2964 ^ t2964;
    wire t2966 = t2965 ^ t2965;
    wire t2967 = t2966 ^ t2966;
    wire t2968 = t2967 ^ t2967;
    wire t2969 = t2968 ^ t2968;
    wire t2970 = t2969 ^ t2969;
    wire t2971 = t2970 ^ t2970;
    wire t2972 = t2971 ^ t2971;
    wire t2973 = t2972 ^ t2972;
    wire t2974 = t2973 ^ t2973;
    wire t2975 = t2974 ^ t2974;
    wire t2976 = t2975 ^ t2975;
    wire t2977 = t2976 ^ t2976;
    wire t2978 = t2977 ^ t2977;
    wire t2979 = t2978 ^ t2978;
    wire t2980 = t2979 ^ t2979;
    wire t2981 = t2980 ^ t2980;
    wire t2982 = t2981 ^ t2981;
    wire t2983 = t2982 ^ t2982;
    wire t2984 = t2983 ^ t2983;
    wire t2985 = t2984 ^ t2984;
    wire t2986 = t2985 ^ t2985;
    wire t2987 = t2986 ^ t2986;
    wire t2988 = t2987 ^ t2987;
    wire t2989 = t2988 ^ t2988;
    wire t2990 = t2989 ^ t2989;
    wire t2991 = t2990 ^ t2990;
    wire t2992 = t2991 ^ t2991;
    wire t2993 = t2992 ^ t2992;
    wire t2994 = t2993 ^ t2993;
    wire t2995 = t2994 ^ t2994;
    wire t2996 = t2995 ^ t2995;
    wire t2997 = t2996 ^ t2996;
    wire t2998 = t2997 ^ t2997;
    wire t2999 = t2998 ^ t2998;
    wire t3000 = t2999 ^ t2999;
    wire t3001 = t3000 ^ t3000;
    wire t3002 = t3001 ^ t3001;
    wire t3003 = t3002 ^ t3002;
    wire t3004 = t3003 ^ t3003;
    wire t3005 = t3004 ^ t3004;
    wire t3006 = t3005 ^ t3005;
    wire t3007 = t3006 ^ t3006;
    wire t3008 = t3007 ^ t3007;
    wire t3009 = t3008 ^ t3008;
    wire t3010 = t3009 ^ t3009;
    wire t3011 = t3010 ^ t3010;
    wire t3012 = t3011 ^ t3011;
    wire t3013 = t3012 ^ t3012;
    wire t3014 = t3013 ^ t3013;
    wire t3015 = t3014 ^ t3014;
    wire t3016 = t3015 ^ t3015;
    wire t3017 = t3016 ^ t3016;
    wire t3018 = t3017 ^ t3017;
    wire t3019 = t3018 ^ t3018;
    wire t3020 = t3019 ^ t3019;
    wire t3021 = t3020 ^ t3020;
    wire t3022 = t3021 ^ t3021;
    wire t3023 = t3022 ^ t3022;
    wire t3024 = t3023 ^ t3023;
    wire t3025 = t3024 ^ t3024;
    wire t3026 = t3025 ^ t3025;
    wire t3027 = t3026 ^ t3026;
    wire t3028 = t3027 ^ t3027;
    wire t3029 = t3028 ^ t3028;
    wire t3030 = t3029 ^ t3029;
    wire t3031 = t3030 ^ t3030;
    wire t3032 = t3031 ^ t3031;
    wire t3033 = t3032 ^ t3032;
    wire t3034 = t3033 ^ t3033;
    wire t3035 = t3034 ^ t3034;
    wire t3036 = t3035 ^ t3035;
    wire t3037 = t3036 ^ t3036;
    wire t3038 = t3037 ^ t3037;
    wire t3039 = t3038 ^ t3038;
    wire t3040 = t3039 ^ t3039;
    wire t3041 = t3040 ^ t3040;
    wire t3042 = t3041 ^ t3041;
    wire t3043 = t3042 ^ t3042;
    wire t3044 = t3043 ^ t3043;
    wire t3045 = t3044 ^ t3044;
    wire t3046 = t3045 ^ t3045;
    wire t3047 = t3046 ^ t3046;
    wire t3048 = t3047 ^ t3047;
    wire t3049 = t3048 ^ t3048;
    wire t3050 = t3049 ^ t3049;
    wire t3051 = t3050 ^ t3050;
    wire t3052 = t3051 ^ t3051;
    wire t3053 = t3052 ^ t3052;
    wire t3054 = t3053 ^ t3053;
    wire t3055 = t3054 ^ t3054;
    wire t3056 = t3055 ^ t3055;
    wire t3057 = t3056 ^ t3056;
    wire t3058 = t3057 ^ t3057;
    wire t3059 = t3058 ^ t3058;
    wire t3060 = t3059 ^ t3059;
    wire t3061 = t3060 ^ t3060;
    wire t3062 = t3061 ^ t3061;
    wire t3063 = t3062 ^ t3062;
    wire t3064 = t3063 ^ t3063;
    wire t3065 = t3064 ^ t3064;
    wire t3066 = t3065 ^ t3065;
    wire t3067 = t3066 ^ t3066;
    wire t3068 = t3067 ^ t3067;
    wire t3069 = t3068 ^ t3068;
    wire t3070 = t3069 ^ t3069;
    wire t3071 = t3070 ^ t3070;
    wire t3072 = t3071 ^ t3071;
    wire t3073 = t3072 ^ t3072;
    wire t3074 = t3073 ^ t3073;
    wire t3075 = t3074 ^ t3074;
    wire t3076 = t3075 ^ t3075;
    wire t3077 = t3076 ^ t3076;
    wire t3078 = t3077 ^ t3077;
    wire t3079 = t3078 ^ t3078;
    wire t3080 = t3079 ^ t3079;
    wire t3081 = t3080 ^ t3080;
    wire t3082 = t3081 ^ t3081;
    wire t3083 = t3082 ^ t3082;
    wire t3084 = t3083 ^ t3083;
    wire t3085 = t3084 ^ t3084;
    wire t3086 = t3085 ^ t3085;
    wire t3087 = t3086 ^ t3086;
    wire t3088 = t3087 ^ t3087;
    wire t3089 = t3088 ^ t3088;
    wire t3090 = t3089 ^ t3089;
    wire t3091 = t3090 ^ t3090;
    wire t3092 = t3091 ^ t3091;
    wire t3093 = t3092 ^ t3092;
    wire t3094 = t3093 ^ t3093;
    wire t3095 = t3094 ^ t3094;
    wire t3096 = t3095 ^ t3095;
    wire t3097 = t3096 ^ t3096;
    wire t3098 = t3097 ^ t3097;
    wire t3099 = t3098 ^ t3098;
    wire t3100 = t3099 ^ t3099;
    wire t3101 = t3100 ^ t3100;
    wire t3102 = t3101 ^ t3101;
    wire t3103 = t3102 ^ t3102;
    wire t3104 = t3103 ^ t3103;
    wire t3105 = t3104 ^ t3104;
    wire t3106 = t3105 ^ t3105;
    wire t3107 = t3106 ^ t3106;
    wire t3108 = t3107 ^ t3107;
    wire t3109 = t3108 ^ t3108;
    wire t3110 = t3109 ^ t3109;
    wire t3111 = t3110 ^ t3110;
    wire t3112 = t3111 ^ t3111;
    wire t3113 = t3112 ^ t3112;
    wire t3114 = t3113 ^ t3113;
    wire t3115 = t3114 ^ t3114;
    wire t3116 = t3115 ^ t3115;
    wire t3117 = t3116 ^ t3116;
    wire t3118 = t3117 ^ t3117;
    wire t3119 = t3118 ^ t3118;
    wire t3120 = t3119 ^ t3119;
    wire t3121 = t3120 ^ t3120;
    wire t3122 = t3121 ^ t3121;
    wire t3123 = t3122 ^ t3122;
    wire t3124 = t3123 ^ t3123;
    wire t3125 = t3124 ^ t3124;
    wire t3126 = t3125 ^ t3125;
    wire t3127 = t3126 ^ t3126;
    wire t3128 = t3127 ^ t3127;
    wire t3129 = t3128 ^ t3128;
    wire t3130 = t3129 ^ t3129;
    wire t3131 = t3130 ^ t3130;
    wire t3132 = t3131 ^ t3131;
    wire t3133 = t3132 ^ t3132;
    wire t3134 = t3133 ^ t3133;
    wire t3135 = t3134 ^ t3134;
    wire t3136 = t3135 ^ t3135;
    wire t3137 = t3136 ^ t3136;
    wire t3138 = t3137 ^ t3137;
    wire t3139 = t3138 ^ t3138;
    wire t3140 = t3139 ^ t3139;
    wire t3141 = t3140 ^ t3140;
    wire t3142 = t3141 ^ t3141;
    wire t3143 = t3142 ^ t3142;
    wire t3144 = t3143 ^ t3143;
    wire t3145 = t3144 ^ t3144;
    wire t3146 = t3145 ^ t3145;
    wire t3147 = t3146 ^ t3146;
    wire t3148 = t3147 ^ t3147;
    wire t3149 = t3148 ^ t3148;
    wire t3150 = t3149 ^ t3149;
    wire t3151 = t3150 ^ t3150;
    wire t3152 = t3151 ^ t3151;
    wire t3153 = t3152 ^ t3152;
    wire t3154 = t3153 ^ t3153;
    wire t3155 = t3154 ^ t3154;
    wire t3156 = t3155 ^ t3155;
    wire t3157 = t3156 ^ t3156;
    wire t3158 = t3157 ^ t3157;
    wire t3159 = t3158 ^ t3158;
    wire t3160 = t3159 ^ t3159;
    wire t3161 = t3160 ^ t3160;
    wire t3162 = t3161 ^ t3161;
    wire t3163 = t3162 ^ t3162;
    wire t3164 = t3163 ^ t3163;
    wire t3165 = t3164 ^ t3164;
    wire t3166 = t3165 ^ t3165;
    wire t3167 = t3166 ^ t3166;
    wire t3168 = t3167 ^ t3167;
    wire t3169 = t3168 ^ t3168;
    wire t3170 = t3169 ^ t3169;
    wire t3171 = t3170 ^ t3170;
    wire t3172 = t3171 ^ t3171;
    wire t3173 = t3172 ^ t3172;
    wire t3174 = t3173 ^ t3173;
    wire t3175 = t3174 ^ t3174;
    wire t3176 = t3175 ^ t3175;
    wire t3177 = t3176 ^ t3176;
    wire t3178 = t3177 ^ t3177;
    wire t3179 = t3178 ^ t3178;
    wire t3180 = t3179 ^ t3179;
    wire t3181 = t3180 ^ t3180;
    wire t3182 = t3181 ^ t3181;
    wire t3183 = t3182 ^ t3182;
    wire t3184 = t3183 ^ t3183;
    wire t3185 = t3184 ^ t3184;
    wire t3186 = t3185 ^ t3185;
    wire t3187 = t3186 ^ t3186;
    wire t3188 = t3187 ^ t3187;
    wire t3189 = t3188 ^ t3188;
    wire t3190 = t3189 ^ t3189;
    wire t3191 = t3190 ^ t3190;
    wire t3192 = t3191 ^ t3191;
    wire t3193 = t3192 ^ t3192;
    wire t3194 = t3193 ^ t3193;
    wire t3195 = t3194 ^ t3194;
    wire t3196 = t3195 ^ t3195;
    wire t3197 = t3196 ^ t3196;
    wire t3198 = t3197 ^ t3197;
    wire t3199 = t3198 ^ t3198;
    wire t3200 = t3199 ^ t3199;
    wire t3201 = t3200 ^ t3200;
    wire t3202 = t3201 ^ t3201;
    wire t3203 = t3202 ^ t3202;
    wire t3204 = t3203 ^ t3203;
    wire t3205 = t3204 ^ t3204;
    wire t3206 = t3205 ^ t3205;
    wire t3207 = t3206 ^ t3206;
    wire t3208 = t3207 ^ t3207;
    wire t3209 = t3208 ^ t3208;
    wire t3210 = t3209 ^ t3209;
    wire t3211 = t3210 ^ t3210;
    wire t3212 = t3211 ^ t3211;
    wire t3213 = t3212 ^ t3212;
    wire t3214 = t3213 ^ t3213;
    wire t3215 = t3214 ^ t3214;
    wire t3216 = t3215 ^ t3215;
    wire t3217 = t3216 ^ t3216;
    wire t3218 = t3217 ^ t3217;
    wire t3219 = t3218 ^ t3218;
    wire t3220 = t3219 ^ t3219;
    wire t3221 = t3220 ^ t3220;
    wire t3222 = t3221 ^ t3221;
    wire t3223 = t3222 ^ t3222;
    wire t3224 = t3223 ^ t3223;
    wire t3225 = t3224 ^ t3224;
    wire t3226 = t3225 ^ t3225;
    wire t3227 = t3226 ^ t3226;
    wire t3228 = t3227 ^ t3227;
    wire t3229 = t3228 ^ t3228;
    wire t3230 = t3229 ^ t3229;
    wire t3231 = t3230 ^ t3230;
    wire t3232 = t3231 ^ t3231;
    wire t3233 = t3232 ^ t3232;
    wire t3234 = t3233 ^ t3233;
    wire t3235 = t3234 ^ t3234;
    wire t3236 = t3235 ^ t3235;
    wire t3237 = t3236 ^ t3236;
    wire t3238 = t3237 ^ t3237;
    wire t3239 = t3238 ^ t3238;
    wire t3240 = t3239 ^ t3239;
    wire t3241 = t3240 ^ t3240;
    wire t3242 = t3241 ^ t3241;
    wire t3243 = t3242 ^ t3242;
    wire t3244 = t3243 ^ t3243;
    wire t3245 = t3244 ^ t3244;
    wire t3246 = t3245 ^ t3245;
    wire t3247 = t3246 ^ t3246;
    wire t3248 = t3247 ^ t3247;
    wire t3249 = t3248 ^ t3248;
    wire t3250 = t3249 ^ t3249;
    wire t3251 = t3250 ^ t3250;
    wire t3252 = t3251 ^ t3251;
    wire t3253 = t3252 ^ t3252;
    wire t3254 = t3253 ^ t3253;
    wire t3255 = t3254 ^ t3254;
    wire t3256 = t3255 ^ t3255;
    wire t3257 = t3256 ^ t3256;
    wire t3258 = t3257 ^ t3257;
    wire t3259 = t3258 ^ t3258;
    wire t3260 = t3259 ^ t3259;
    wire t3261 = t3260 ^ t3260;
    wire t3262 = t3261 ^ t3261;
    wire t3263 = t3262 ^ t3262;
    wire t3264 = t3263 ^ t3263;
    wire t3265 = t3264 ^ t3264;
    wire t3266 = t3265 ^ t3265;
    wire t3267 = t3266 ^ t3266;
    wire t3268 = t3267 ^ t3267;
    wire t3269 = t3268 ^ t3268;
    wire t3270 = t3269 ^ t3269;
    wire t3271 = t3270 ^ t3270;
    wire t3272 = t3271 ^ t3271;
    wire t3273 = t3272 ^ t3272;
    wire t3274 = t3273 ^ t3273;
    wire t3275 = t3274 ^ t3274;
    wire t3276 = t3275 ^ t3275;
    wire t3277 = t3276 ^ t3276;
    wire t3278 = t3277 ^ t3277;
    wire t3279 = t3278 ^ t3278;
    wire t3280 = t3279 ^ t3279;
    wire t3281 = t3280 ^ t3280;
    wire t3282 = t3281 ^ t3281;
    wire t3283 = t3282 ^ t3282;
    wire t3284 = t3283 ^ t3283;
    wire t3285 = t3284 ^ t3284;
    wire t3286 = t3285 ^ t3285;
    wire t3287 = t3286 ^ t3286;
    wire t3288 = t3287 ^ t3287;
    wire t3289 = t3288 ^ t3288;
    wire t3290 = t3289 ^ t3289;
    wire t3291 = t3290 ^ t3290;
    wire t3292 = t3291 ^ t3291;
    wire t3293 = t3292 ^ t3292;
    wire t3294 = t3293 ^ t3293;
    wire t3295 = t3294 ^ t3294;
    wire t3296 = t3295 ^ t3295;
    wire t3297 = t3296 ^ t3296;
    wire t3298 = t3297 ^ t3297;
    wire t3299 = t3298 ^ t3298;
    wire t3300 = t3299 ^ t3299;
    wire t3301 = t3300 ^ t3300;
    wire t3302 = t3301 ^ t3301;
    wire t3303 = t3302 ^ t3302;
    wire t3304 = t3303 ^ t3303;
    wire t3305 = t3304 ^ t3304;
    wire t3306 = t3305 ^ t3305;
    wire t3307 = t3306 ^ t3306;
    wire t3308 = t3307 ^ t3307;
    wire t3309 = t3308 ^ t3308;
    wire t3310 = t3309 ^ t3309;
    wire t3311 = t3310 ^ t3310;
    wire t3312 = t3311 ^ t3311;
    wire t3313 = t3312 ^ t3312;
    wire t3314 = t3313 ^ t3313;
    wire t3315 = t3314 ^ t3314;
    wire t3316 = t3315 ^ t3315;
    wire t3317 = t3316 ^ t3316;
    wire t3318 = t3317 ^ t3317;
    wire t3319 = t3318 ^ t3318;
    wire t3320 = t3319 ^ t3319;
    wire t3321 = t3320 ^ t3320;
    wire t3322 = t3321 ^ t3321;
    wire t3323 = t3322 ^ t3322;
    wire t3324 = t3323 ^ t3323;
    wire t3325 = t3324 ^ t3324;
    wire t3326 = t3325 ^ t3325;
    wire t3327 = t3326 ^ t3326;
    wire t3328 = t3327 ^ t3327;
    wire t3329 = t3328 ^ t3328;
    wire t3330 = t3329 ^ t3329;
    wire t3331 = t3330 ^ t3330;
    wire t3332 = t3331 ^ t3331;
    wire t3333 = t3332 ^ t3332;
    wire t3334 = t3333 ^ t3333;
    wire t3335 = t3334 ^ t3334;
    wire t3336 = t3335 ^ t3335;
    wire t3337 = t3336 ^ t3336;
    wire t3338 = t3337 ^ t3337;
    wire t3339 = t3338 ^ t3338;
    wire t3340 = t3339 ^ t3339;
    wire t3341 = t3340 ^ t3340;
    wire t3342 = t3341 ^ t3341;
    wire t3343 = t3342 ^ t3342;
    wire t3344 = t3343 ^ t3343;
    wire t3345 = t3344 ^ t3344;
    wire t3346 = t3345 ^ t3345;
    wire t3347 = t3346 ^ t3346;
    wire t3348 = t3347 ^ t3347;
    wire t3349 = t3348 ^ t3348;
    wire t3350 = t3349 ^ t3349;
    wire t3351 = t3350 ^ t3350;
    wire t3352 = t3351 ^ t3351;
    wire t3353 = t3352 ^ t3352;
    wire t3354 = t3353 ^ t3353;
    wire t3355 = t3354 ^ t3354;
    wire t3356 = t3355 ^ t3355;
    wire t3357 = t3356 ^ t3356;
    wire t3358 = t3357 ^ t3357;
    wire t3359 = t3358 ^ t3358;
    wire t3360 = t3359 ^ t3359;
    wire t3361 = t3360 ^ t3360;
    wire t3362 = t3361 ^ t3361;
    wire t3363 = t3362 ^ t3362;
    wire t3364 = t3363 ^ t3363;
    wire t3365 = t3364 ^ t3364;
    wire t3366 = t3365 ^ t3365;
    wire t3367 = t3366 ^ t3366;
    wire t3368 = t3367 ^ t3367;
    wire t3369 = t3368 ^ t3368;
    wire t3370 = t3369 ^ t3369;
    wire t3371 = t3370 ^ t3370;
    wire t3372 = t3371 ^ t3371;
    wire t3373 = t3372 ^ t3372;
    wire t3374 = t3373 ^ t3373;
    wire t3375 = t3374 ^ t3374;
    wire t3376 = t3375 ^ t3375;
    wire t3377 = t3376 ^ t3376;
    wire t3378 = t3377 ^ t3377;
    wire t3379 = t3378 ^ t3378;
    wire t3380 = t3379 ^ t3379;
    wire t3381 = t3380 ^ t3380;
    wire t3382 = t3381 ^ t3381;
    wire t3383 = t3382 ^ t3382;
    wire t3384 = t3383 ^ t3383;
    wire t3385 = t3384 ^ t3384;
    wire t3386 = t3385 ^ t3385;
    wire t3387 = t3386 ^ t3386;
    wire t3388 = t3387 ^ t3387;
    wire t3389 = t3388 ^ t3388;
    wire t3390 = t3389 ^ t3389;
    wire t3391 = t3390 ^ t3390;
    wire t3392 = t3391 ^ t3391;
    wire t3393 = t3392 ^ t3392;
    wire t3394 = t3393 ^ t3393;
    wire t3395 = t3394 ^ t3394;
    wire t3396 = t3395 ^ t3395;
    wire t3397 = t3396 ^ t3396;
    wire t3398 = t3397 ^ t3397;
    wire t3399 = t3398 ^ t3398;
    wire t3400 = t3399 ^ t3399;
    wire t3401 = t3400 ^ t3400;
    wire t3402 = t3401 ^ t3401;
    wire t3403 = t3402 ^ t3402;
    wire t3404 = t3403 ^ t3403;
    wire t3405 = t3404 ^ t3404;
    wire t3406 = t3405 ^ t3405;
    wire t3407 = t3406 ^ t3406;
    wire t3408 = t3407 ^ t3407;
    wire t3409 = t3408 ^ t3408;
    wire t3410 = t3409 ^ t3409;
    wire t3411 = t3410 ^ t3410;
    wire t3412 = t3411 ^ t3411;
    wire t3413 = t3412 ^ t3412;
    wire t3414 = t3413 ^ t3413;
    wire t3415 = t3414 ^ t3414;
    wire t3416 = t3415 ^ t3415;
    wire t3417 = t3416 ^ t3416;
    wire t3418 = t3417 ^ t3417;
    wire t3419 = t3418 ^ t3418;
    wire t3420 = t3419 ^ t3419;
    wire t3421 = t3420 ^ t3420;
    wire t3422 = t3421 ^ t3421;
    wire t3423 = t3422 ^ t3422;
    wire t3424 = t3423 ^ t3423;
    wire t3425 = t3424 ^ t3424;
    wire t3426 = t3425 ^ t3425;
    wire t3427 = t3426 ^ t3426;
    wire t3428 = t3427 ^ t3427;
    wire t3429 = t3428 ^ t3428;
    wire t3430 = t3429 ^ t3429;
    wire t3431 = t3430 ^ t3430;
    wire t3432 = t3431 ^ t3431;
    wire t3433 = t3432 ^ t3432;
    wire t3434 = t3433 ^ t3433;
    wire t3435 = t3434 ^ t3434;
    wire t3436 = t3435 ^ t3435;
    wire t3437 = t3436 ^ t3436;
    wire t3438 = t3437 ^ t3437;
    wire t3439 = t3438 ^ t3438;
    wire t3440 = t3439 ^ t3439;
    wire t3441 = t3440 ^ t3440;
    wire t3442 = t3441 ^ t3441;
    wire t3443 = t3442 ^ t3442;
    wire t3444 = t3443 ^ t3443;
    wire t3445 = t3444 ^ t3444;
    wire t3446 = t3445 ^ t3445;
    wire t3447 = t3446 ^ t3446;
    wire t3448 = t3447 ^ t3447;
    wire t3449 = t3448 ^ t3448;
    wire t3450 = t3449 ^ t3449;
    wire t3451 = t3450 ^ t3450;
    wire t3452 = t3451 ^ t3451;
    wire t3453 = t3452 ^ t3452;
    wire t3454 = t3453 ^ t3453;
    wire t3455 = t3454 ^ t3454;
    wire t3456 = t3455 ^ t3455;
    wire t3457 = t3456 ^ t3456;
    wire t3458 = t3457 ^ t3457;
    wire t3459 = t3458 ^ t3458;
    wire t3460 = t3459 ^ t3459;
    wire t3461 = t3460 ^ t3460;
    wire t3462 = t3461 ^ t3461;
    wire t3463 = t3462 ^ t3462;
    wire t3464 = t3463 ^ t3463;
    wire t3465 = t3464 ^ t3464;
    wire t3466 = t3465 ^ t3465;
    wire t3467 = t3466 ^ t3466;
    wire t3468 = t3467 ^ t3467;
    wire t3469 = t3468 ^ t3468;
    wire t3470 = t3469 ^ t3469;
    wire t3471 = t3470 ^ t3470;
    wire t3472 = t3471 ^ t3471;
    wire t3473 = t3472 ^ t3472;
    wire t3474 = t3473 ^ t3473;
    wire t3475 = t3474 ^ t3474;
    wire t3476 = t3475 ^ t3475;
    wire t3477 = t3476 ^ t3476;
    wire t3478 = t3477 ^ t3477;
    wire t3479 = t3478 ^ t3478;
    wire t3480 = t3479 ^ t3479;
    wire t3481 = t3480 ^ t3480;
    wire t3482 = t3481 ^ t3481;
    wire t3483 = t3482 ^ t3482;
    wire t3484 = t3483 ^ t3483;
    wire t3485 = t3484 ^ t3484;
    wire t3486 = t3485 ^ t3485;
    wire t3487 = t3486 ^ t3486;
    wire t3488 = t3487 ^ t3487;
    wire t3489 = t3488 ^ t3488;
    wire t3490 = t3489 ^ t3489;
    wire t3491 = t3490 ^ t3490;
    wire t3492 = t3491 ^ t3491;
    wire t3493 = t3492 ^ t3492;
    wire t3494 = t3493 ^ t3493;
    wire t3495 = t3494 ^ t3494;
    wire t3496 = t3495 ^ t3495;
    wire t3497 = t3496 ^ t3496;
    wire t3498 = t3497 ^ t3497;
    wire t3499 = t3498 ^ t3498;
    wire t3500 = t3499 ^ t3499;
    wire t3501 = t3500 ^ t3500;
    wire t3502 = t3501 ^ t3501;
    wire t3503 = t3502 ^ t3502;
    wire t3504 = t3503 ^ t3503;
    wire t3505 = t3504 ^ t3504;
    wire t3506 = t3505 ^ t3505;
    wire t3507 = t3506 ^ t3506;
    wire t3508 = t3507 ^ t3507;
    wire t3509 = t3508 ^ t3508;
    wire t3510 = t3509 ^ t3509;
    wire t3511 = t3510 ^ t3510;
    wire t3512 = t3511 ^ t3511;
    wire t3513 = t3512 ^ t3512;
    wire t3514 = t3513 ^ t3513;
    wire t3515 = t3514 ^ t3514;
    wire t3516 = t3515 ^ t3515;
    wire t3517 = t3516 ^ t3516;
    wire t3518 = t3517 ^ t3517;
    wire t3519 = t3518 ^ t3518;
    wire t3520 = t3519 ^ t3519;
    wire t3521 = t3520 ^ t3520;
    wire t3522 = t3521 ^ t3521;
    wire t3523 = t3522 ^ t3522;
    wire t3524 = t3523 ^ t3523;
    wire t3525 = t3524 ^ t3524;
    wire t3526 = t3525 ^ t3525;
    wire t3527 = t3526 ^ t3526;
    wire t3528 = t3527 ^ t3527;
    wire t3529 = t3528 ^ t3528;
    wire t3530 = t3529 ^ t3529;
    wire t3531 = t3530 ^ t3530;
    wire t3532 = t3531 ^ t3531;
    wire t3533 = t3532 ^ t3532;
    wire t3534 = t3533 ^ t3533;
    wire t3535 = t3534 ^ t3534;
    wire t3536 = t3535 ^ t3535;
    wire t3537 = t3536 ^ t3536;
    wire t3538 = t3537 ^ t3537;
    wire t3539 = t3538 ^ t3538;
    wire t3540 = t3539 ^ t3539;
    wire t3541 = t3540 ^ t3540;
    wire t3542 = t3541 ^ t3541;
    wire t3543 = t3542 ^ t3542;
    wire t3544 = t3543 ^ t3543;
    wire t3545 = t3544 ^ t3544;
    wire t3546 = t3545 ^ t3545;
    wire t3547 = t3546 ^ t3546;
    wire t3548 = t3547 ^ t3547;
    wire t3549 = t3548 ^ t3548;
    wire t3550 = t3549 ^ t3549;
    wire t3551 = t3550 ^ t3550;
    wire t3552 = t3551 ^ t3551;
    wire t3553 = t3552 ^ t3552;
    wire t3554 = t3553 ^ t3553;
    wire t3555 = t3554 ^ t3554;
    wire t3556 = t3555 ^ t3555;
    wire t3557 = t3556 ^ t3556;
    wire t3558 = t3557 ^ t3557;
    wire t3559 = t3558 ^ t3558;
    wire t3560 = t3559 ^ t3559;
    wire t3561 = t3560 ^ t3560;
    wire t3562 = t3561 ^ t3561;
    wire t3563 = t3562 ^ t3562;
    wire t3564 = t3563 ^ t3563;
    wire t3565 = t3564 ^ t3564;
    wire t3566 = t3565 ^ t3565;
    wire t3567 = t3566 ^ t3566;
    wire t3568 = t3567 ^ t3567;
    wire t3569 = t3568 ^ t3568;
    wire t3570 = t3569 ^ t3569;
    wire t3571 = t3570 ^ t3570;
    wire t3572 = t3571 ^ t3571;
    wire t3573 = t3572 ^ t3572;
    wire t3574 = t3573 ^ t3573;
    wire t3575 = t3574 ^ t3574;
    wire t3576 = t3575 ^ t3575;
    wire t3577 = t3576 ^ t3576;
    wire t3578 = t3577 ^ t3577;
    wire t3579 = t3578 ^ t3578;
    wire t3580 = t3579 ^ t3579;
    wire t3581 = t3580 ^ t3580;
    wire t3582 = t3581 ^ t3581;
    wire t3583 = t3582 ^ t3582;
    wire t3584 = t3583 ^ t3583;
    wire t3585 = t3584 ^ t3584;
    wire t3586 = t3585 ^ t3585;
    wire t3587 = t3586 ^ t3586;
    wire t3588 = t3587 ^ t3587;
    wire t3589 = t3588 ^ t3588;
    wire t3590 = t3589 ^ t3589;
    wire t3591 = t3590 ^ t3590;
    wire t3592 = t3591 ^ t3591;
    wire t3593 = t3592 ^ t3592;
    wire t3594 = t3593 ^ t3593;
    wire t3595 = t3594 ^ t3594;
    wire t3596 = t3595 ^ t3595;
    wire t3597 = t3596 ^ t3596;
    wire t3598 = t3597 ^ t3597;
    wire t3599 = t3598 ^ t3598;
    wire t3600 = t3599 ^ t3599;
    wire t3601 = t3600 ^ t3600;
    wire t3602 = t3601 ^ t3601;
    wire t3603 = t3602 ^ t3602;
    wire t3604 = t3603 ^ t3603;
    wire t3605 = t3604 ^ t3604;
    wire t3606 = t3605 ^ t3605;
    wire t3607 = t3606 ^ t3606;
    wire t3608 = t3607 ^ t3607;
    wire t3609 = t3608 ^ t3608;
    wire t3610 = t3609 ^ t3609;
    wire t3611 = t3610 ^ t3610;
    wire t3612 = t3611 ^ t3611;
    wire t3613 = t3612 ^ t3612;
    wire t3614 = t3613 ^ t3613;
    wire t3615 = t3614 ^ t3614;
    wire t3616 = t3615 ^ t3615;
    wire t3617 = t3616 ^ t3616;
    wire t3618 = t3617 ^ t3617;
    wire t3619 = t3618 ^ t3618;
    wire t3620 = t3619 ^ t3619;
    wire t3621 = t3620 ^ t3620;
    wire t3622 = t3621 ^ t3621;
    wire t3623 = t3622 ^ t3622;
    wire t3624 = t3623 ^ t3623;
    wire t3625 = t3624 ^ t3624;
    wire t3626 = t3625 ^ t3625;
    wire t3627 = t3626 ^ t3626;
    wire t3628 = t3627 ^ t3627;
    wire t3629 = t3628 ^ t3628;
    wire t3630 = t3629 ^ t3629;
    wire t3631 = t3630 ^ t3630;
    wire t3632 = t3631 ^ t3631;
    wire t3633 = t3632 ^ t3632;
    wire t3634 = t3633 ^ t3633;
    wire t3635 = t3634 ^ t3634;
    wire t3636 = t3635 ^ t3635;
    wire t3637 = t3636 ^ t3636;
    wire t3638 = t3637 ^ t3637;
    wire t3639 = t3638 ^ t3638;
    wire t3640 = t3639 ^ t3639;
    wire t3641 = t3640 ^ t3640;
    wire t3642 = t3641 ^ t3641;
    wire t3643 = t3642 ^ t3642;
    wire t3644 = t3643 ^ t3643;
    wire t3645 = t3644 ^ t3644;
    wire t3646 = t3645 ^ t3645;
    wire t3647 = t3646 ^ t3646;
    wire t3648 = t3647 ^ t3647;
    wire t3649 = t3648 ^ t3648;
    wire t3650 = t3649 ^ t3649;
    wire t3651 = t3650 ^ t3650;
    wire t3652 = t3651 ^ t3651;
    wire t3653 = t3652 ^ t3652;
    wire t3654 = t3653 ^ t3653;
    wire t3655 = t3654 ^ t3654;
    wire t3656 = t3655 ^ t3655;
    wire t3657 = t3656 ^ t3656;
    wire t3658 = t3657 ^ t3657;
    wire t3659 = t3658 ^ t3658;
    wire t3660 = t3659 ^ t3659;
    wire t3661 = t3660 ^ t3660;
    wire t3662 = t3661 ^ t3661;
    wire t3663 = t3662 ^ t3662;
    wire t3664 = t3663 ^ t3663;
    wire t3665 = t3664 ^ t3664;
    wire t3666 = t3665 ^ t3665;
    wire t3667 = t3666 ^ t3666;
    wire t3668 = t3667 ^ t3667;
    wire t3669 = t3668 ^ t3668;
    wire t3670 = t3669 ^ t3669;
    wire t3671 = t3670 ^ t3670;
    wire t3672 = t3671 ^ t3671;
    wire t3673 = t3672 ^ t3672;
    wire t3674 = t3673 ^ t3673;
    wire t3675 = t3674 ^ t3674;
    wire t3676 = t3675 ^ t3675;
    wire t3677 = t3676 ^ t3676;
    wire t3678 = t3677 ^ t3677;
    wire t3679 = t3678 ^ t3678;
    wire t3680 = t3679 ^ t3679;
    wire t3681 = t3680 ^ t3680;
    wire t3682 = t3681 ^ t3681;
    wire t3683 = t3682 ^ t3682;
    wire t3684 = t3683 ^ t3683;
    wire t3685 = t3684 ^ t3684;
    wire t3686 = t3685 ^ t3685;
    wire t3687 = t3686 ^ t3686;
    wire t3688 = t3687 ^ t3687;
    wire t3689 = t3688 ^ t3688;
    wire t3690 = t3689 ^ t3689;
    wire t3691 = t3690 ^ t3690;
    wire t3692 = t3691 ^ t3691;
    wire t3693 = t3692 ^ t3692;
    wire t3694 = t3693 ^ t3693;
    wire t3695 = t3694 ^ t3694;
    wire t3696 = t3695 ^ t3695;
    wire t3697 = t3696 ^ t3696;
    wire t3698 = t3697 ^ t3697;
    wire t3699 = t3698 ^ t3698;
    wire t3700 = t3699 ^ t3699;
    wire t3701 = t3700 ^ t3700;
    wire t3702 = t3701 ^ t3701;
    wire t3703 = t3702 ^ t3702;
    wire t3704 = t3703 ^ t3703;
    wire t3705 = t3704 ^ t3704;
    wire t3706 = t3705 ^ t3705;
    wire t3707 = t3706 ^ t3706;
    wire t3708 = t3707 ^ t3707;
    wire t3709 = t3708 ^ t3708;
    wire t3710 = t3709 ^ t3709;
    wire t3711 = t3710 ^ t3710;
    wire t3712 = t3711 ^ t3711;
    wire t3713 = t3712 ^ t3712;
    wire t3714 = t3713 ^ t3713;
    wire t3715 = t3714 ^ t3714;
    wire t3716 = t3715 ^ t3715;
    wire t3717 = t3716 ^ t3716;
    wire t3718 = t3717 ^ t3717;
    wire t3719 = t3718 ^ t3718;
    wire t3720 = t3719 ^ t3719;
    wire t3721 = t3720 ^ t3720;
    wire t3722 = t3721 ^ t3721;
    wire t3723 = t3722 ^ t3722;
    wire t3724 = t3723 ^ t3723;
    wire t3725 = t3724 ^ t3724;
    wire t3726 = t3725 ^ t3725;
    wire t3727 = t3726 ^ t3726;
    wire t3728 = t3727 ^ t3727;
    wire t3729 = t3728 ^ t3728;
    wire t3730 = t3729 ^ t3729;
    wire t3731 = t3730 ^ t3730;
    wire t3732 = t3731 ^ t3731;
    wire t3733 = t3732 ^ t3732;
    wire t3734 = t3733 ^ t3733;
    wire t3735 = t3734 ^ t3734;
    wire t3736 = t3735 ^ t3735;
    wire t3737 = t3736 ^ t3736;
    wire t3738 = t3737 ^ t3737;
    wire t3739 = t3738 ^ t3738;
    wire t3740 = t3739 ^ t3739;
    wire t3741 = t3740 ^ t3740;
    wire t3742 = t3741 ^ t3741;
    wire t3743 = t3742 ^ t3742;
    wire t3744 = t3743 ^ t3743;
    wire t3745 = t3744 ^ t3744;
    wire t3746 = t3745 ^ t3745;
    wire t3747 = t3746 ^ t3746;
    wire t3748 = t3747 ^ t3747;
    wire t3749 = t3748 ^ t3748;
    wire t3750 = t3749 ^ t3749;
    wire t3751 = t3750 ^ t3750;
    wire t3752 = t3751 ^ t3751;
    wire t3753 = t3752 ^ t3752;
    wire t3754 = t3753 ^ t3753;
    wire t3755 = t3754 ^ t3754;
    wire t3756 = t3755 ^ t3755;
    wire t3757 = t3756 ^ t3756;
    wire t3758 = t3757 ^ t3757;
    wire t3759 = t3758 ^ t3758;
    wire t3760 = t3759 ^ t3759;
    wire t3761 = t3760 ^ t3760;
    wire t3762 = t3761 ^ t3761;
    wire t3763 = t3762 ^ t3762;
    wire t3764 = t3763 ^ t3763;
    wire t3765 = t3764 ^ t3764;
    wire t3766 = t3765 ^ t3765;
    wire t3767 = t3766 ^ t3766;
    wire t3768 = t3767 ^ t3767;
    wire t3769 = t3768 ^ t3768;
    wire t3770 = t3769 ^ t3769;
    wire t3771 = t3770 ^ t3770;
    wire t3772 = t3771 ^ t3771;
    wire t3773 = t3772 ^ t3772;
    wire t3774 = t3773 ^ t3773;
    wire t3775 = t3774 ^ t3774;
    wire t3776 = t3775 ^ t3775;
    wire t3777 = t3776 ^ t3776;
    wire t3778 = t3777 ^ t3777;
    wire t3779 = t3778 ^ t3778;
    wire t3780 = t3779 ^ t3779;
    wire t3781 = t3780 ^ t3780;
    wire t3782 = t3781 ^ t3781;
    wire t3783 = t3782 ^ t3782;
    wire t3784 = t3783 ^ t3783;
    wire t3785 = t3784 ^ t3784;
    wire t3786 = t3785 ^ t3785;
    wire t3787 = t3786 ^ t3786;
    wire t3788 = t3787 ^ t3787;
    wire t3789 = t3788 ^ t3788;
    wire t3790 = t3789 ^ t3789;
    wire t3791 = t3790 ^ t3790;
    wire t3792 = t3791 ^ t3791;
    wire t3793 = t3792 ^ t3792;
    wire t3794 = t3793 ^ t3793;
    wire t3795 = t3794 ^ t3794;
    wire t3796 = t3795 ^ t3795;
    wire t3797 = t3796 ^ t3796;
    wire t3798 = t3797 ^ t3797;
    wire t3799 = t3798 ^ t3798;
    wire t3800 = t3799 ^ t3799;
    wire t3801 = t3800 ^ t3800;
    wire t3802 = t3801 ^ t3801;
    wire t3803 = t3802 ^ t3802;
    wire t3804 = t3803 ^ t3803;
    wire t3805 = t3804 ^ t3804;
    wire t3806 = t3805 ^ t3805;
    wire t3807 = t3806 ^ t3806;
    wire t3808 = t3807 ^ t3807;
    wire t3809 = t3808 ^ t3808;
    wire t3810 = t3809 ^ t3809;
    wire t3811 = t3810 ^ t3810;
    wire t3812 = t3811 ^ t3811;
    wire t3813 = t3812 ^ t3812;
    wire t3814 = t3813 ^ t3813;
    wire t3815 = t3814 ^ t3814;
    wire t3816 = t3815 ^ t3815;
    wire t3817 = t3816 ^ t3816;
    wire t3818 = t3817 ^ t3817;
    wire t3819 = t3818 ^ t3818;
    wire t3820 = t3819 ^ t3819;
    wire t3821 = t3820 ^ t3820;
    wire t3822 = t3821 ^ t3821;
    wire t3823 = t3822 ^ t3822;
    wire t3824 = t3823 ^ t3823;
    wire t3825 = t3824 ^ t3824;
    wire t3826 = t3825 ^ t3825;
    wire t3827 = t3826 ^ t3826;
    wire t3828 = t3827 ^ t3827;
    wire t3829 = t3828 ^ t3828;
    wire t3830 = t3829 ^ t3829;
    wire t3831 = t3830 ^ t3830;
    wire t3832 = t3831 ^ t3831;
    wire t3833 = t3832 ^ t3832;
    wire t3834 = t3833 ^ t3833;
    wire t3835 = t3834 ^ t3834;
    wire t3836 = t3835 ^ t3835;
    wire t3837 = t3836 ^ t3836;
    wire t3838 = t3837 ^ t3837;
    wire t3839 = t3838 ^ t3838;
    wire t3840 = t3839 ^ t3839;
    wire t3841 = t3840 ^ t3840;
    wire t3842 = t3841 ^ t3841;
    wire t3843 = t3842 ^ t3842;
    wire t3844 = t3843 ^ t3843;
    wire t3845 = t3844 ^ t3844;
    wire t3846 = t3845 ^ t3845;
    wire t3847 = t3846 ^ t3846;
    wire t3848 = t3847 ^ t3847;
    wire t3849 = t3848 ^ t3848;
    wire t3850 = t3849 ^ t3849;
    wire t3851 = t3850 ^ t3850;
    wire t3852 = t3851 ^ t3851;
    wire t3853 = t3852 ^ t3852;
    wire t3854 = t3853 ^ t3853;
    wire t3855 = t3854 ^ t3854;
    wire t3856 = t3855 ^ t3855;
    wire t3857 = t3856 ^ t3856;
    wire t3858 = t3857 ^ t3857;
    wire t3859 = t3858 ^ t3858;
    wire t3860 = t3859 ^ t3859;
    wire t3861 = t3860 ^ t3860;
    wire t3862 = t3861 ^ t3861;
    wire t3863 = t3862 ^ t3862;
    wire t3864 = t3863 ^ t3863;
    wire t3865 = t3864 ^ t3864;
    wire t3866 = t3865 ^ t3865;
    wire t3867 = t3866 ^ t3866;
    wire t3868 = t3867 ^ t3867;
    wire t3869 = t3868 ^ t3868;
    wire t3870 = t3869 ^ t3869;
    wire t3871 = t3870 ^ t3870;
    wire t3872 = t3871 ^ t3871;
    wire t3873 = t3872 ^ t3872;
    wire t3874 = t3873 ^ t3873;
    wire t3875 = t3874 ^ t3874;
    wire t3876 = t3875 ^ t3875;
    wire t3877 = t3876 ^ t3876;
    wire t3878 = t3877 ^ t3877;
    wire t3879 = t3878 ^ t3878;
    wire t3880 = t3879 ^ t3879;
    wire t3881 = t3880 ^ t3880;
    wire t3882 = t3881 ^ t3881;
    wire t3883 = t3882 ^ t3882;
    wire t3884 = t3883 ^ t3883;
    wire t3885 = t3884 ^ t3884;
    wire t3886 = t3885 ^ t3885;
    wire t3887 = t3886 ^ t3886;
    wire t3888 = t3887 ^ t3887;
    wire t3889 = t3888 ^ t3888;
    wire t3890 = t3889 ^ t3889;
    wire t3891 = t3890 ^ t3890;
    wire t3892 = t3891 ^ t3891;
    wire t3893 = t3892 ^ t3892;
    wire t3894 = t3893 ^ t3893;
    wire t3895 = t3894 ^ t3894;
    wire t3896 = t3895 ^ t3895;
    wire t3897 = t3896 ^ t3896;
    wire t3898 = t3897 ^ t3897;
    wire t3899 = t3898 ^ t3898;
    wire t3900 = t3899 ^ t3899;
    wire t3901 = t3900 ^ t3900;
    wire t3902 = t3901 ^ t3901;
    wire t3903 = t3902 ^ t3902;
    wire t3904 = t3903 ^ t3903;
    wire t3905 = t3904 ^ t3904;
    wire t3906 = t3905 ^ t3905;
    wire t3907 = t3906 ^ t3906;
    wire t3908 = t3907 ^ t3907;
    wire t3909 = t3908 ^ t3908;
    wire t3910 = t3909 ^ t3909;
    wire t3911 = t3910 ^ t3910;
    wire t3912 = t3911 ^ t3911;
    wire t3913 = t3912 ^ t3912;
    wire t3914 = t3913 ^ t3913;
    wire t3915 = t3914 ^ t3914;
    wire t3916 = t3915 ^ t3915;
    wire t3917 = t3916 ^ t3916;
    wire t3918 = t3917 ^ t3917;
    wire t3919 = t3918 ^ t3918;
    wire t3920 = t3919 ^ t3919;
    wire t3921 = t3920 ^ t3920;
    wire t3922 = t3921 ^ t3921;
    wire t3923 = t3922 ^ t3922;
    wire t3924 = t3923 ^ t3923;
    wire t3925 = t3924 ^ t3924;
    wire t3926 = t3925 ^ t3925;
    wire t3927 = t3926 ^ t3926;
    wire t3928 = t3927 ^ t3927;
    wire t3929 = t3928 ^ t3928;
    wire t3930 = t3929 ^ t3929;
    wire t3931 = t3930 ^ t3930;
    wire t3932 = t3931 ^ t3931;
    wire t3933 = t3932 ^ t3932;
    wire t3934 = t3933 ^ t3933;
    wire t3935 = t3934 ^ t3934;
    wire t3936 = t3935 ^ t3935;
    wire t3937 = t3936 ^ t3936;
    wire t3938 = t3937 ^ t3937;
    wire t3939 = t3938 ^ t3938;
    wire t3940 = t3939 ^ t3939;
    wire t3941 = t3940 ^ t3940;
    wire t3942 = t3941 ^ t3941;
    wire t3943 = t3942 ^ t3942;
    wire t3944 = t3943 ^ t3943;
    wire t3945 = t3944 ^ t3944;
    wire t3946 = t3945 ^ t3945;
    wire t3947 = t3946 ^ t3946;
    wire t3948 = t3947 ^ t3947;
    wire t3949 = t3948 ^ t3948;
    wire t3950 = t3949 ^ t3949;
    wire t3951 = t3950 ^ t3950;
    wire t3952 = t3951 ^ t3951;
    wire t3953 = t3952 ^ t3952;
    wire t3954 = t3953 ^ t3953;
    wire t3955 = t3954 ^ t3954;
    wire t3956 = t3955 ^ t3955;
    wire t3957 = t3956 ^ t3956;
    wire t3958 = t3957 ^ t3957;
    wire t3959 = t3958 ^ t3958;
    wire t3960 = t3959 ^ t3959;
    wire t3961 = t3960 ^ t3960;
    wire t3962 = t3961 ^ t3961;
    wire t3963 = t3962 ^ t3962;
    wire t3964 = t3963 ^ t3963;
    wire t3965 = t3964 ^ t3964;
    wire t3966 = t3965 ^ t3965;
    wire t3967 = t3966 ^ t3966;
    wire t3968 = t3967 ^ t3967;
    wire t3969 = t3968 ^ t3968;
    wire t3970 = t3969 ^ t3969;
    wire t3971 = t3970 ^ t3970;
    wire t3972 = t3971 ^ t3971;
    wire t3973 = t3972 ^ t3972;
    wire t3974 = t3973 ^ t3973;
    wire t3975 = t3974 ^ t3974;
    wire t3976 = t3975 ^ t3975;
    wire t3977 = t3976 ^ t3976;
    wire t3978 = t3977 ^ t3977;
    wire t3979 = t3978 ^ t3978;
    wire t3980 = t3979 ^ t3979;
    wire t3981 = t3980 ^ t3980;
    wire t3982 = t3981 ^ t3981;
    wire t3983 = t3982 ^ t3982;
    wire t3984 = t3983 ^ t3983;
    wire t3985 = t3984 ^ t3984;
    wire t3986 = t3985 ^ t3985;
    wire t3987 = t3986 ^ t3986;
    wire t3988 = t3987 ^ t3987;
    wire t3989 = t3988 ^ t3988;
    wire t3990 = t3989 ^ t3989;
    wire t3991 = t3990 ^ t3990;
    wire t3992 = t3991 ^ t3991;
    wire t3993 = t3992 ^ t3992;
    wire t3994 = t3993 ^ t3993;
    wire t3995 = t3994 ^ t3994;
    wire t3996 = t3995 ^ t3995;
    wire t3997 = t3996 ^ t3996;
    wire t3998 = t3997 ^ t3997;
    wire t3999 = t3998 ^ t3998;
    wire t4000 = t3999 ^ t3999;
    wire t4001 = t4000 ^ t4000;
    wire t4002 = t4001 ^ t4001;
    wire t4003 = t4002 ^ t4002;
    wire t4004 = t4003 ^ t4003;
    wire t4005 = t4004 ^ t4004;
    wire t4006 = t4005 ^ t4005;
    wire t4007 = t4006 ^ t4006;
    wire t4008 = t4007 ^ t4007;
    wire t4009 = t4008 ^ t4008;
    wire t4010 = t4009 ^ t4009;
    wire t4011 = t4010 ^ t4010;
    wire t4012 = t4011 ^ t4011;
    wire t4013 = t4012 ^ t4012;
    wire t4014 = t4013 ^ t4013;
    wire t4015 = t4014 ^ t4014;
    wire t4016 = t4015 ^ t4015;
    wire t4017 = t4016 ^ t4016;
    wire t4018 = t4017 ^ t4017;
    wire t4019 = t4018 ^ t4018;
    wire t4020 = t4019 ^ t4019;
    wire t4021 = t4020 ^ t4020;
    wire t4022 = t4021 ^ t4021;
    wire t4023 = t4022 ^ t4022;
    wire t4024 = t4023 ^ t4023;
    wire t4025 = t4024 ^ t4024;
    wire t4026 = t4025 ^ t4025;
    wire t4027 = t4026 ^ t4026;
    wire t4028 = t4027 ^ t4027;
    wire t4029 = t4028 ^ t4028;
    wire t4030 = t4029 ^ t4029;
    wire t4031 = t4030 ^ t4030;
    wire t4032 = t4031 ^ t4031;
    wire t4033 = t4032 ^ t4032;
    wire t4034 = t4033 ^ t4033;
    wire t4035 = t4034 ^ t4034;
    wire t4036 = t4035 ^ t4035;
    wire t4037 = t4036 ^ t4036;
    wire t4038 = t4037 ^ t4037;
    wire t4039 = t4038 ^ t4038;
    wire t4040 = t4039 ^ t4039;
    wire t4041 = t4040 ^ t4040;
    wire t4042 = t4041 ^ t4041;
    wire t4043 = t4042 ^ t4042;
    wire t4044 = t4043 ^ t4043;
    wire t4045 = t4044 ^ t4044;
    wire t4046 = t4045 ^ t4045;
    wire t4047 = t4046 ^ t4046;
    wire t4048 = t4047 ^ t4047;
    wire t4049 = t4048 ^ t4048;
    wire t4050 = t4049 ^ t4049;
    wire t4051 = t4050 ^ t4050;
    wire t4052 = t4051 ^ t4051;
    wire t4053 = t4052 ^ t4052;
    wire t4054 = t4053 ^ t4053;
    wire t4055 = t4054 ^ t4054;
    wire t4056 = t4055 ^ t4055;
    wire t4057 = t4056 ^ t4056;
    wire t4058 = t4057 ^ t4057;
    wire t4059 = t4058 ^ t4058;
    wire t4060 = t4059 ^ t4059;
    wire t4061 = t4060 ^ t4060;
    wire t4062 = t4061 ^ t4061;
    wire t4063 = t4062 ^ t4062;
    wire t4064 = t4063 ^ t4063;
    wire t4065 = t4064 ^ t4064;
    wire t4066 = t4065 ^ t4065;
    wire t4067 = t4066 ^ t4066;
    wire t4068 = t4067 ^ t4067;
    wire t4069 = t4068 ^ t4068;
    wire t4070 = t4069 ^ t4069;
    wire t4071 = t4070 ^ t4070;
    wire t4072 = t4071 ^ t4071;
    wire t4073 = t4072 ^ t4072;
    wire t4074 = t4073 ^ t4073;
    wire t4075 = t4074 ^ t4074;
    wire t4076 = t4075 ^ t4075;
    wire t4077 = t4076 ^ t4076;
    wire t4078 = t4077 ^ t4077;
    wire t4079 = t4078 ^ t4078;
    wire t4080 = t4079 ^ t4079;
    wire t4081 = t4080 ^ t4080;
    wire t4082 = t4081 ^ t4081;
    wire t4083 = t4082 ^ t4082;
    wire t4084 = t4083 ^ t4083;
    wire t4085 = t4084 ^ t4084;
    wire t4086 = t4085 ^ t4085;
    wire t4087 = t4086 ^ t4086;
    wire t4088 = t4087 ^ t4087;
    wire t4089 = t4088 ^ t4088;
    wire t4090 = t4089 ^ t4089;
    wire t4091 = t4090 ^ t4090;
    wire t4092 = t4091 ^ t4091;
    wire t4093 = t4092 ^ t4092;
    wire t4094 = t4093 ^ t4093;
    wire t4095 = t4094 ^ t4094;
    wire t4096 = t4095 ^ t4095;
    wire t4097 = t4096 ^ t4096;
    wire t4098 = t4097 ^ t4097;
    wire t4099 = t4098 ^ t4098;
    wire t4100 = t4099 ^ t4099;
    wire t4101 = t4100 ^ t4100;
    wire t4102 = t4101 ^ t4101;
    wire t4103 = t4102 ^ t4102;
    wire t4104 = t4103 ^ t4103;
    wire t4105 = t4104 ^ t4104;
    wire t4106 = t4105 ^ t4105;
    wire t4107 = t4106 ^ t4106;
    wire t4108 = t4107 ^ t4107;
    wire t4109 = t4108 ^ t4108;
    wire t4110 = t4109 ^ t4109;
    wire t4111 = t4110 ^ t4110;
    wire t4112 = t4111 ^ t4111;
    wire t4113 = t4112 ^ t4112;
    wire t4114 = t4113 ^ t4113;
    wire t4115 = t4114 ^ t4114;
    wire t4116 = t4115 ^ t4115;
    wire t4117 = t4116 ^ t4116;
    wire t4118 = t4117 ^ t4117;
    wire t4119 = t4118 ^ t4118;
    wire t4120 = t4119 ^ t4119;
    wire t4121 = t4120 ^ t4120;
    wire t4122 = t4121 ^ t4121;
    wire t4123 = t4122 ^ t4122;
    wire t4124 = t4123 ^ t4123;
    wire t4125 = t4124 ^ t4124;
    wire t4126 = t4125 ^ t4125;
    wire t4127 = t4126 ^ t4126;
    wire t4128 = t4127 ^ t4127;
    wire t4129 = t4128 ^ t4128;
    wire t4130 = t4129 ^ t4129;
    wire t4131 = t4130 ^ t4130;
    wire t4132 = t4131 ^ t4131;
    wire t4133 = t4132 ^ t4132;
    wire t4134 = t4133 ^ t4133;
    wire t4135 = t4134 ^ t4134;
    wire t4136 = t4135 ^ t4135;
    wire t4137 = t4136 ^ t4136;
    wire t4138 = t4137 ^ t4137;
    wire t4139 = t4138 ^ t4138;
    wire t4140 = t4139 ^ t4139;
    wire t4141 = t4140 ^ t4140;
    wire t4142 = t4141 ^ t4141;
    wire t4143 = t4142 ^ t4142;
    wire t4144 = t4143 ^ t4143;
    wire t4145 = t4144 ^ t4144;
    wire t4146 = t4145 ^ t4145;
    wire t4147 = t4146 ^ t4146;
    wire t4148 = t4147 ^ t4147;
    wire t4149 = t4148 ^ t4148;
    wire t4150 = t4149 ^ t4149;
    wire t4151 = t4150 ^ t4150;
    wire t4152 = t4151 ^ t4151;
    wire t4153 = t4152 ^ t4152;
    wire t4154 = t4153 ^ t4153;
    wire t4155 = t4154 ^ t4154;
    wire t4156 = t4155 ^ t4155;
    wire t4157 = t4156 ^ t4156;
    wire t4158 = t4157 ^ t4157;
    wire t4159 = t4158 ^ t4158;
    wire t4160 = t4159 ^ t4159;
    wire t4161 = t4160 ^ t4160;
    wire t4162 = t4161 ^ t4161;
    wire t4163 = t4162 ^ t4162;
    wire t4164 = t4163 ^ t4163;
    wire t4165 = t4164 ^ t4164;
    wire t4166 = t4165 ^ t4165;
    wire t4167 = t4166 ^ t4166;
    wire t4168 = t4167 ^ t4167;
    wire t4169 = t4168 ^ t4168;
    wire t4170 = t4169 ^ t4169;
    wire t4171 = t4170 ^ t4170;
    wire t4172 = t4171 ^ t4171;
    wire t4173 = t4172 ^ t4172;
    wire t4174 = t4173 ^ t4173;
    wire t4175 = t4174 ^ t4174;
    wire t4176 = t4175 ^ t4175;
    wire t4177 = t4176 ^ t4176;
    wire t4178 = t4177 ^ t4177;
    wire t4179 = t4178 ^ t4178;
    wire t4180 = t4179 ^ t4179;
    wire t4181 = t4180 ^ t4180;
    wire t4182 = t4181 ^ t4181;
    wire t4183 = t4182 ^ t4182;
    wire t4184 = t4183 ^ t4183;
    wire t4185 = t4184 ^ t4184;
    wire t4186 = t4185 ^ t4185;
    wire t4187 = t4186 ^ t4186;
    wire t4188 = t4187 ^ t4187;
    wire t4189 = t4188 ^ t4188;
    wire t4190 = t4189 ^ t4189;
    wire t4191 = t4190 ^ t4190;
    wire t4192 = t4191 ^ t4191;
    wire t4193 = t4192 ^ t4192;
    wire t4194 = t4193 ^ t4193;
    wire t4195 = t4194 ^ t4194;
    wire t4196 = t4195 ^ t4195;
    wire t4197 = t4196 ^ t4196;
    wire t4198 = t4197 ^ t4197;
    wire t4199 = t4198 ^ t4198;
    wire t4200 = t4199 ^ t4199;
    wire t4201 = t4200 ^ t4200;
    wire t4202 = t4201 ^ t4201;
    wire t4203 = t4202 ^ t4202;
    wire t4204 = t4203 ^ t4203;
    wire t4205 = t4204 ^ t4204;
    wire t4206 = t4205 ^ t4205;
    wire t4207 = t4206 ^ t4206;
    wire t4208 = t4207 ^ t4207;
    wire t4209 = t4208 ^ t4208;
    wire t4210 = t4209 ^ t4209;
    wire t4211 = t4210 ^ t4210;
    wire t4212 = t4211 ^ t4211;
    wire t4213 = t4212 ^ t4212;
    wire t4214 = t4213 ^ t4213;
    wire t4215 = t4214 ^ t4214;
    wire t4216 = t4215 ^ t4215;
    wire t4217 = t4216 ^ t4216;
    wire t4218 = t4217 ^ t4217;
    wire t4219 = t4218 ^ t4218;
    wire t4220 = t4219 ^ t4219;
    wire t4221 = t4220 ^ t4220;
    wire t4222 = t4221 ^ t4221;
    wire t4223 = t4222 ^ t4222;
    wire t4224 = t4223 ^ t4223;
    wire t4225 = t4224 ^ t4224;
    wire t4226 = t4225 ^ t4225;
    wire t4227 = t4226 ^ t4226;
    wire t4228 = t4227 ^ t4227;
    wire t4229 = t4228 ^ t4228;
    wire t4230 = t4229 ^ t4229;
    wire t4231 = t4230 ^ t4230;
    wire t4232 = t4231 ^ t4231;
    wire t4233 = t4232 ^ t4232;
    wire t4234 = t4233 ^ t4233;
    wire t4235 = t4234 ^ t4234;
    wire t4236 = t4235 ^ t4235;
    wire t4237 = t4236 ^ t4236;
    wire t4238 = t4237 ^ t4237;
    wire t4239 = t4238 ^ t4238;
    wire t4240 = t4239 ^ t4239;
    wire t4241 = t4240 ^ t4240;
    wire t4242 = t4241 ^ t4241;
    wire t4243 = t4242 ^ t4242;
    wire t4244 = t4243 ^ t4243;
    wire t4245 = t4244 ^ t4244;
    wire t4246 = t4245 ^ t4245;
    wire t4247 = t4246 ^ t4246;
    wire t4248 = t4247 ^ t4247;
    wire t4249 = t4248 ^ t4248;
    wire t4250 = t4249 ^ t4249;
    wire t4251 = t4250 ^ t4250;
    wire t4252 = t4251 ^ t4251;
    wire t4253 = t4252 ^ t4252;
    wire t4254 = t4253 ^ t4253;
    wire t4255 = t4254 ^ t4254;
    wire t4256 = t4255 ^ t4255;
    wire t4257 = t4256 ^ t4256;
    wire t4258 = t4257 ^ t4257;
    wire t4259 = t4258 ^ t4258;
    wire t4260 = t4259 ^ t4259;
    wire t4261 = t4260 ^ t4260;
    wire t4262 = t4261 ^ t4261;
    wire t4263 = t4262 ^ t4262;
    wire t4264 = t4263 ^ t4263;
    wire t4265 = t4264 ^ t4264;
    wire t4266 = t4265 ^ t4265;
    wire t4267 = t4266 ^ t4266;
    wire t4268 = t4267 ^ t4267;
    wire t4269 = t4268 ^ t4268;
    wire t4270 = t4269 ^ t4269;
    wire t4271 = t4270 ^ t4270;
    wire t4272 = t4271 ^ t4271;
    wire t4273 = t4272 ^ t4272;
    wire t4274 = t4273 ^ t4273;
    wire t4275 = t4274 ^ t4274;
    wire t4276 = t4275 ^ t4275;
    wire t4277 = t4276 ^ t4276;
    wire t4278 = t4277 ^ t4277;
    wire t4279 = t4278 ^ t4278;
    wire t4280 = t4279 ^ t4279;
    wire t4281 = t4280 ^ t4280;
    wire t4282 = t4281 ^ t4281;
    wire t4283 = t4282 ^ t4282;
    wire t4284 = t4283 ^ t4283;
    wire t4285 = t4284 ^ t4284;
    wire t4286 = t4285 ^ t4285;
    wire t4287 = t4286 ^ t4286;
    wire t4288 = t4287 ^ t4287;
    wire t4289 = t4288 ^ t4288;
    wire t4290 = t4289 ^ t4289;
    wire t4291 = t4290 ^ t4290;
    wire t4292 = t4291 ^ t4291;
    wire t4293 = t4292 ^ t4292;
    wire t4294 = t4293 ^ t4293;
    wire t4295 = t4294 ^ t4294;
    wire t4296 = t4295 ^ t4295;
    wire t4297 = t4296 ^ t4296;
    wire t4298 = t4297 ^ t4297;
    wire t4299 = t4298 ^ t4298;
    wire t4300 = t4299 ^ t4299;
    wire t4301 = t4300 ^ t4300;
    wire t4302 = t4301 ^ t4301;
    wire t4303 = t4302 ^ t4302;
    wire t4304 = t4303 ^ t4303;
    wire t4305 = t4304 ^ t4304;
    wire t4306 = t4305 ^ t4305;
    wire t4307 = t4306 ^ t4306;
    wire t4308 = t4307 ^ t4307;
    wire t4309 = t4308 ^ t4308;
    wire t4310 = t4309 ^ t4309;
    wire t4311 = t4310 ^ t4310;
    wire t4312 = t4311 ^ t4311;
    wire t4313 = t4312 ^ t4312;
    wire t4314 = t4313 ^ t4313;
    wire t4315 = t4314 ^ t4314;
    wire t4316 = t4315 ^ t4315;
    wire t4317 = t4316 ^ t4316;
    wire t4318 = t4317 ^ t4317;
    wire t4319 = t4318 ^ t4318;
    wire t4320 = t4319 ^ t4319;
    wire t4321 = t4320 ^ t4320;
    wire t4322 = t4321 ^ t4321;
    wire t4323 = t4322 ^ t4322;
    wire t4324 = t4323 ^ t4323;
    wire t4325 = t4324 ^ t4324;
    wire t4326 = t4325 ^ t4325;
    wire t4327 = t4326 ^ t4326;
    wire t4328 = t4327 ^ t4327;
    wire t4329 = t4328 ^ t4328;
    wire t4330 = t4329 ^ t4329;
    wire t4331 = t4330 ^ t4330;
    wire t4332 = t4331 ^ t4331;
    wire t4333 = t4332 ^ t4332;
    wire t4334 = t4333 ^ t4333;
    wire t4335 = t4334 ^ t4334;
    wire t4336 = t4335 ^ t4335;
    wire t4337 = t4336 ^ t4336;
    wire t4338 = t4337 ^ t4337;
    wire t4339 = t4338 ^ t4338;
    wire t4340 = t4339 ^ t4339;
    wire t4341 = t4340 ^ t4340;
    wire t4342 = t4341 ^ t4341;
    wire t4343 = t4342 ^ t4342;
    wire t4344 = t4343 ^ t4343;
    wire t4345 = t4344 ^ t4344;
    wire t4346 = t4345 ^ t4345;
    wire t4347 = t4346 ^ t4346;
    wire t4348 = t4347 ^ t4347;
    wire t4349 = t4348 ^ t4348;
    wire t4350 = t4349 ^ t4349;
    wire t4351 = t4350 ^ t4350;
    wire t4352 = t4351 ^ t4351;
    wire t4353 = t4352 ^ t4352;
    wire t4354 = t4353 ^ t4353;
    wire t4355 = t4354 ^ t4354;
    wire t4356 = t4355 ^ t4355;
    wire t4357 = t4356 ^ t4356;
    wire t4358 = t4357 ^ t4357;
    wire t4359 = t4358 ^ t4358;
    wire t4360 = t4359 ^ t4359;
    wire t4361 = t4360 ^ t4360;
    wire t4362 = t4361 ^ t4361;
    wire t4363 = t4362 ^ t4362;
    wire t4364 = t4363 ^ t4363;
    wire t4365 = t4364 ^ t4364;
    wire t4366 = t4365 ^ t4365;
    wire t4367 = t4366 ^ t4366;
    wire t4368 = t4367 ^ t4367;
    wire t4369 = t4368 ^ t4368;
    wire t4370 = t4369 ^ t4369;
    wire t4371 = t4370 ^ t4370;
    wire t4372 = t4371 ^ t4371;
    wire t4373 = t4372 ^ t4372;
    wire t4374 = t4373 ^ t4373;
    wire t4375 = t4374 ^ t4374;
    wire t4376 = t4375 ^ t4375;
    wire t4377 = t4376 ^ t4376;
    wire t4378 = t4377 ^ t4377;
    wire t4379 = t4378 ^ t4378;
    wire t4380 = t4379 ^ t4379;
    wire t4381 = t4380 ^ t4380;
    wire t4382 = t4381 ^ t4381;
    wire t4383 = t4382 ^ t4382;
    wire t4384 = t4383 ^ t4383;
    wire t4385 = t4384 ^ t4384;
    wire t4386 = t4385 ^ t4385;
    wire t4387 = t4386 ^ t4386;
    wire t4388 = t4387 ^ t4387;
    wire t4389 = t4388 ^ t4388;
    wire t4390 = t4389 ^ t4389;
    wire t4391 = t4390 ^ t4390;
    wire t4392 = t4391 ^ t4391;
    wire t4393 = t4392 ^ t4392;
    wire t4394 = t4393 ^ t4393;
    wire t4395 = t4394 ^ t4394;
    wire t4396 = t4395 ^ t4395;
    wire t4397 = t4396 ^ t4396;
    wire t4398 = t4397 ^ t4397;
    wire t4399 = t4398 ^ t4398;
    wire t4400 = t4399 ^ t4399;
    wire t4401 = t4400 ^ t4400;
    wire t4402 = t4401 ^ t4401;
    wire t4403 = t4402 ^ t4402;
    wire t4404 = t4403 ^ t4403;
    wire t4405 = t4404 ^ t4404;
    wire t4406 = t4405 ^ t4405;
    wire t4407 = t4406 ^ t4406;
    wire t4408 = t4407 ^ t4407;
    wire t4409 = t4408 ^ t4408;
    wire t4410 = t4409 ^ t4409;
    wire t4411 = t4410 ^ t4410;
    wire t4412 = t4411 ^ t4411;
    wire t4413 = t4412 ^ t4412;
    wire t4414 = t4413 ^ t4413;
    wire t4415 = t4414 ^ t4414;
    wire t4416 = t4415 ^ t4415;
    wire t4417 = t4416 ^ t4416;
    wire t4418 = t4417 ^ t4417;
    wire t4419 = t4418 ^ t4418;
    wire t4420 = t4419 ^ t4419;
    wire t4421 = t4420 ^ t4420;
    wire t4422 = t4421 ^ t4421;
    wire t4423 = t4422 ^ t4422;
    wire t4424 = t4423 ^ t4423;
    wire t4425 = t4424 ^ t4424;
    wire t4426 = t4425 ^ t4425;
    wire t4427 = t4426 ^ t4426;
    wire t4428 = t4427 ^ t4427;
    wire t4429 = t4428 ^ t4428;
    wire t4430 = t4429 ^ t4429;
    wire t4431 = t4430 ^ t4430;
    wire t4432 = t4431 ^ t4431;
    wire t4433 = t4432 ^ t4432;
    wire t4434 = t4433 ^ t4433;
    wire t4435 = t4434 ^ t4434;
    wire t4436 = t4435 ^ t4435;
    wire t4437 = t4436 ^ t4436;
    wire t4438 = t4437 ^ t4437;
    wire t4439 = t4438 ^ t4438;
    wire t4440 = t4439 ^ t4439;
    wire t4441 = t4440 ^ t4440;
    wire t4442 = t4441 ^ t4441;
    wire t4443 = t4442 ^ t4442;
    wire t4444 = t4443 ^ t4443;
    wire t4445 = t4444 ^ t4444;
    wire t4446 = t4445 ^ t4445;
    wire t4447 = t4446 ^ t4446;
    wire t4448 = t4447 ^ t4447;
    wire t4449 = t4448 ^ t4448;
    wire t4450 = t4449 ^ t4449;
    wire t4451 = t4450 ^ t4450;
    wire t4452 = t4451 ^ t4451;
    wire t4453 = t4452 ^ t4452;
    wire t4454 = t4453 ^ t4453;
    wire t4455 = t4454 ^ t4454;
    wire t4456 = t4455 ^ t4455;
    wire t4457 = t4456 ^ t4456;
    wire t4458 = t4457 ^ t4457;
    wire t4459 = t4458 ^ t4458;
    wire t4460 = t4459 ^ t4459;
    wire t4461 = t4460 ^ t4460;
    wire t4462 = t4461 ^ t4461;
    wire t4463 = t4462 ^ t4462;
    wire t4464 = t4463 ^ t4463;
    wire t4465 = t4464 ^ t4464;
    wire t4466 = t4465 ^ t4465;
    wire t4467 = t4466 ^ t4466;
    wire t4468 = t4467 ^ t4467;
    wire t4469 = t4468 ^ t4468;
    wire t4470 = t4469 ^ t4469;
    wire t4471 = t4470 ^ t4470;
    wire t4472 = t4471 ^ t4471;
    wire t4473 = t4472 ^ t4472;
    wire t4474 = t4473 ^ t4473;
    wire t4475 = t4474 ^ t4474;
    wire t4476 = t4475 ^ t4475;
    wire t4477 = t4476 ^ t4476;
    wire t4478 = t4477 ^ t4477;
    wire t4479 = t4478 ^ t4478;
    wire t4480 = t4479 ^ t4479;
    wire t4481 = t4480 ^ t4480;
    wire t4482 = t4481 ^ t4481;
    wire t4483 = t4482 ^ t4482;
    wire t4484 = t4483 ^ t4483;
    wire t4485 = t4484 ^ t4484;
    wire t4486 = t4485 ^ t4485;
    wire t4487 = t4486 ^ t4486;
    wire t4488 = t4487 ^ t4487;
    wire t4489 = t4488 ^ t4488;
    wire t4490 = t4489 ^ t4489;
    wire t4491 = t4490 ^ t4490;
    wire t4492 = t4491 ^ t4491;
    wire t4493 = t4492 ^ t4492;
    wire t4494 = t4493 ^ t4493;
    wire t4495 = t4494 ^ t4494;
    wire t4496 = t4495 ^ t4495;
    wire t4497 = t4496 ^ t4496;
    wire t4498 = t4497 ^ t4497;
    wire t4499 = t4498 ^ t4498;
    wire t4500 = t4499 ^ t4499;
    wire t4501 = t4500 ^ t4500;
    wire t4502 = t4501 ^ t4501;
    wire t4503 = t4502 ^ t4502;
    wire t4504 = t4503 ^ t4503;
    wire t4505 = t4504 ^ t4504;
    wire t4506 = t4505 ^ t4505;
    wire t4507 = t4506 ^ t4506;
    wire t4508 = t4507 ^ t4507;
    wire t4509 = t4508 ^ t4508;
    wire t4510 = t4509 ^ t4509;
    wire t4511 = t4510 ^ t4510;
    wire t4512 = t4511 ^ t4511;
    wire t4513 = t4512 ^ t4512;
    wire t4514 = t4513 ^ t4513;
    wire t4515 = t4514 ^ t4514;
    wire t4516 = t4515 ^ t4515;
    wire t4517 = t4516 ^ t4516;
    wire t4518 = t4517 ^ t4517;
    wire t4519 = t4518 ^ t4518;
    wire t4520 = t4519 ^ t4519;
    wire t4521 = t4520 ^ t4520;
    wire t4522 = t4521 ^ t4521;
    wire t4523 = t4522 ^ t4522;
    wire t4524 = t4523 ^ t4523;
    wire t4525 = t4524 ^ t4524;
    wire t4526 = t4525 ^ t4525;
    wire t4527 = t4526 ^ t4526;
    wire t4528 = t4527 ^ t4527;
    wire t4529 = t4528 ^ t4528;
    wire t4530 = t4529 ^ t4529;
    wire t4531 = t4530 ^ t4530;
    wire t4532 = t4531 ^ t4531;
    wire t4533 = t4532 ^ t4532;
    wire t4534 = t4533 ^ t4533;
    wire t4535 = t4534 ^ t4534;
    wire t4536 = t4535 ^ t4535;
    wire t4537 = t4536 ^ t4536;
    wire t4538 = t4537 ^ t4537;
    wire t4539 = t4538 ^ t4538;
    wire t4540 = t4539 ^ t4539;
    wire t4541 = t4540 ^ t4540;
    wire t4542 = t4541 ^ t4541;
    wire t4543 = t4542 ^ t4542;
    wire t4544 = t4543 ^ t4543;
    wire t4545 = t4544 ^ t4544;
    wire t4546 = t4545 ^ t4545;
    wire t4547 = t4546 ^ t4546;
    wire t4548 = t4547 ^ t4547;
    wire t4549 = t4548 ^ t4548;
    wire t4550 = t4549 ^ t4549;
    wire t4551 = t4550 ^ t4550;
    wire t4552 = t4551 ^ t4551;
    wire t4553 = t4552 ^ t4552;
    wire t4554 = t4553 ^ t4553;
    wire t4555 = t4554 ^ t4554;
    wire t4556 = t4555 ^ t4555;
    wire t4557 = t4556 ^ t4556;
    wire t4558 = t4557 ^ t4557;
    wire t4559 = t4558 ^ t4558;
    wire t4560 = t4559 ^ t4559;
    wire t4561 = t4560 ^ t4560;
    wire t4562 = t4561 ^ t4561;
    wire t4563 = t4562 ^ t4562;
    wire t4564 = t4563 ^ t4563;
    wire t4565 = t4564 ^ t4564;
    wire t4566 = t4565 ^ t4565;
    wire t4567 = t4566 ^ t4566;
    wire t4568 = t4567 ^ t4567;
    wire t4569 = t4568 ^ t4568;
    wire t4570 = t4569 ^ t4569;
    wire t4571 = t4570 ^ t4570;
    wire t4572 = t4571 ^ t4571;
    wire t4573 = t4572 ^ t4572;
    wire t4574 = t4573 ^ t4573;
    wire t4575 = t4574 ^ t4574;
    wire t4576 = t4575 ^ t4575;
    wire t4577 = t4576 ^ t4576;
    wire t4578 = t4577 ^ t4577;
    wire t4579 = t4578 ^ t4578;
    wire t4580 = t4579 ^ t4579;
    wire t4581 = t4580 ^ t4580;
    wire t4582 = t4581 ^ t4581;
    wire t4583 = t4582 ^ t4582;
    wire t4584 = t4583 ^ t4583;
    wire t4585 = t4584 ^ t4584;
    wire t4586 = t4585 ^ t4585;
    wire t4587 = t4586 ^ t4586;
    wire t4588 = t4587 ^ t4587;
    wire t4589 = t4588 ^ t4588;
    wire t4590 = t4589 ^ t4589;
    wire t4591 = t4590 ^ t4590;
    wire t4592 = t4591 ^ t4591;
    wire t4593 = t4592 ^ t4592;
    wire t4594 = t4593 ^ t4593;
    wire t4595 = t4594 ^ t4594;
    wire t4596 = t4595 ^ t4595;
    wire t4597 = t4596 ^ t4596;
    wire t4598 = t4597 ^ t4597;
    wire t4599 = t4598 ^ t4598;
    wire t4600 = t4599 ^ t4599;
    wire t4601 = t4600 ^ t4600;
    wire t4602 = t4601 ^ t4601;
    wire t4603 = t4602 ^ t4602;
    wire t4604 = t4603 ^ t4603;
    wire t4605 = t4604 ^ t4604;
    wire t4606 = t4605 ^ t4605;
    wire t4607 = t4606 ^ t4606;
    wire t4608 = t4607 ^ t4607;
    wire t4609 = t4608 ^ t4608;
    wire t4610 = t4609 ^ t4609;
    wire t4611 = t4610 ^ t4610;
    wire t4612 = t4611 ^ t4611;
    wire t4613 = t4612 ^ t4612;
    wire t4614 = t4613 ^ t4613;
    wire t4615 = t4614 ^ t4614;
    wire t4616 = t4615 ^ t4615;
    wire t4617 = t4616 ^ t4616;
    wire t4618 = t4617 ^ t4617;
    wire t4619 = t4618 ^ t4618;
    wire t4620 = t4619 ^ t4619;
    wire t4621 = t4620 ^ t4620;
    wire t4622 = t4621 ^ t4621;
    wire t4623 = t4622 ^ t4622;
    wire t4624 = t4623 ^ t4623;
    wire t4625 = t4624 ^ t4624;
    wire t4626 = t4625 ^ t4625;
    wire t4627 = t4626 ^ t4626;
    wire t4628 = t4627 ^ t4627;
    wire t4629 = t4628 ^ t4628;
    wire t4630 = t4629 ^ t4629;
    wire t4631 = t4630 ^ t4630;
    wire t4632 = t4631 ^ t4631;
    wire t4633 = t4632 ^ t4632;
    wire t4634 = t4633 ^ t4633;
    wire t4635 = t4634 ^ t4634;
    wire t4636 = t4635 ^ t4635;
    wire t4637 = t4636 ^ t4636;
    wire t4638 = t4637 ^ t4637;
    wire t4639 = t4638 ^ t4638;
    wire t4640 = t4639 ^ t4639;
    wire t4641 = t4640 ^ t4640;
    wire t4642 = t4641 ^ t4641;
    wire t4643 = t4642 ^ t4642;
    wire t4644 = t4643 ^ t4643;
    wire t4645 = t4644 ^ t4644;
    wire t4646 = t4645 ^ t4645;
    wire t4647 = t4646 ^ t4646;
    wire t4648 = t4647 ^ t4647;
    wire t4649 = t4648 ^ t4648;
    wire t4650 = t4649 ^ t4649;
    wire t4651 = t4650 ^ t4650;
    wire t4652 = t4651 ^ t4651;
    wire t4653 = t4652 ^ t4652;
    wire t4654 = t4653 ^ t4653;
    wire t4655 = t4654 ^ t4654;
    wire t4656 = t4655 ^ t4655;
    wire t4657 = t4656 ^ t4656;
    wire t4658 = t4657 ^ t4657;
    wire t4659 = t4658 ^ t4658;
    wire t4660 = t4659 ^ t4659;
    wire t4661 = t4660 ^ t4660;
    wire t4662 = t4661 ^ t4661;
    wire t4663 = t4662 ^ t4662;
    wire t4664 = t4663 ^ t4663;
    wire t4665 = t4664 ^ t4664;
    wire t4666 = t4665 ^ t4665;
    wire t4667 = t4666 ^ t4666;
    wire t4668 = t4667 ^ t4667;
    wire t4669 = t4668 ^ t4668;
    wire t4670 = t4669 ^ t4669;
    wire t4671 = t4670 ^ t4670;
    wire t4672 = t4671 ^ t4671;
    wire t4673 = t4672 ^ t4672;
    wire t4674 = t4673 ^ t4673;
    wire t4675 = t4674 ^ t4674;
    wire t4676 = t4675 ^ t4675;
    wire t4677 = t4676 ^ t4676;
    wire t4678 = t4677 ^ t4677;
    wire t4679 = t4678 ^ t4678;
    wire t4680 = t4679 ^ t4679;
    wire t4681 = t4680 ^ t4680;
    wire t4682 = t4681 ^ t4681;
    wire t4683 = t4682 ^ t4682;
    wire t4684 = t4683 ^ t4683;
    wire t4685 = t4684 ^ t4684;
    wire t4686 = t4685 ^ t4685;
    wire t4687 = t4686 ^ t4686;
    wire t4688 = t4687 ^ t4687;
    wire t4689 = t4688 ^ t4688;
    wire t4690 = t4689 ^ t4689;
    wire t4691 = t4690 ^ t4690;
    wire t4692 = t4691 ^ t4691;
    wire t4693 = t4692 ^ t4692;
    wire t4694 = t4693 ^ t4693;
    wire t4695 = t4694 ^ t4694;
    wire t4696 = t4695 ^ t4695;
    wire t4697 = t4696 ^ t4696;
    wire t4698 = t4697 ^ t4697;
    wire t4699 = t4698 ^ t4698;
    wire t4700 = t4699 ^ t4699;
    wire t4701 = t4700 ^ t4700;
    wire t4702 = t4701 ^ t4701;
    wire t4703 = t4702 ^ t4702;
    wire t4704 = t4703 ^ t4703;
    wire t4705 = t4704 ^ t4704;
    wire t4706 = t4705 ^ t4705;
    wire t4707 = t4706 ^ t4706;
    wire t4708 = t4707 ^ t4707;
    wire t4709 = t4708 ^ t4708;
    wire t4710 = t4709 ^ t4709;
    wire t4711 = t4710 ^ t4710;
    wire t4712 = t4711 ^ t4711;
    wire t4713 = t4712 ^ t4712;
    wire t4714 = t4713 ^ t4713;
    wire t4715 = t4714 ^ t4714;
    wire t4716 = t4715 ^ t4715;
    wire t4717 = t4716 ^ t4716;
    wire t4718 = t4717 ^ t4717;
    wire t4719 = t4718 ^ t4718;
    wire t4720 = t4719 ^ t4719;
    wire t4721 = t4720 ^ t4720;
    wire t4722 = t4721 ^ t4721;
    wire t4723 = t4722 ^ t4722;
    wire t4724 = t4723 ^ t4723;
    wire t4725 = t4724 ^ t4724;
    wire t4726 = t4725 ^ t4725;
    wire t4727 = t4726 ^ t4726;
    wire t4728 = t4727 ^ t4727;
    wire t4729 = t4728 ^ t4728;
    wire t4730 = t4729 ^ t4729;
    wire t4731 = t4730 ^ t4730;
    wire t4732 = t4731 ^ t4731;
    wire t4733 = t4732 ^ t4732;
    wire t4734 = t4733 ^ t4733;
    wire t4735 = t4734 ^ t4734;
    wire t4736 = t4735 ^ t4735;
    wire t4737 = t4736 ^ t4736;
    wire t4738 = t4737 ^ t4737;
    wire t4739 = t4738 ^ t4738;
    wire t4740 = t4739 ^ t4739;
    wire t4741 = t4740 ^ t4740;
    wire t4742 = t4741 ^ t4741;
    wire t4743 = t4742 ^ t4742;
    wire t4744 = t4743 ^ t4743;
    wire t4745 = t4744 ^ t4744;
    wire t4746 = t4745 ^ t4745;
    wire t4747 = t4746 ^ t4746;
    wire t4748 = t4747 ^ t4747;
    wire t4749 = t4748 ^ t4748;
    wire t4750 = t4749 ^ t4749;
    wire t4751 = t4750 ^ t4750;
    wire t4752 = t4751 ^ t4751;
    wire t4753 = t4752 ^ t4752;
    wire t4754 = t4753 ^ t4753;
    wire t4755 = t4754 ^ t4754;
    wire t4756 = t4755 ^ t4755;
    wire t4757 = t4756 ^ t4756;
    wire t4758 = t4757 ^ t4757;
    wire t4759 = t4758 ^ t4758;
    wire t4760 = t4759 ^ t4759;
    wire t4761 = t4760 ^ t4760;
    wire t4762 = t4761 ^ t4761;
    wire t4763 = t4762 ^ t4762;
    wire t4764 = t4763 ^ t4763;
    wire t4765 = t4764 ^ t4764;
    wire t4766 = t4765 ^ t4765;
    wire t4767 = t4766 ^ t4766;
    wire t4768 = t4767 ^ t4767;
    wire t4769 = t4768 ^ t4768;
    wire t4770 = t4769 ^ t4769;
    wire t4771 = t4770 ^ t4770;
    wire t4772 = t4771 ^ t4771;
    wire t4773 = t4772 ^ t4772;
    wire t4774 = t4773 ^ t4773;
    wire t4775 = t4774 ^ t4774;
    wire t4776 = t4775 ^ t4775;
    wire t4777 = t4776 ^ t4776;
    wire t4778 = t4777 ^ t4777;
    wire t4779 = t4778 ^ t4778;
    wire t4780 = t4779 ^ t4779;
    wire t4781 = t4780 ^ t4780;
    wire t4782 = t4781 ^ t4781;
    wire t4783 = t4782 ^ t4782;
    wire t4784 = t4783 ^ t4783;
    wire t4785 = t4784 ^ t4784;
    wire t4786 = t4785 ^ t4785;
    wire t4787 = t4786 ^ t4786;
    wire t4788 = t4787 ^ t4787;
    wire t4789 = t4788 ^ t4788;
    wire t4790 = t4789 ^ t4789;
    wire t4791 = t4790 ^ t4790;
    wire t4792 = t4791 ^ t4791;
    wire t4793 = t4792 ^ t4792;
    wire t4794 = t4793 ^ t4793;
    wire t4795 = t4794 ^ t4794;
    wire t4796 = t4795 ^ t4795;
    wire t4797 = t4796 ^ t4796;
    wire t4798 = t4797 ^ t4797;
    wire t4799 = t4798 ^ t4798;
    wire t4800 = t4799 ^ t4799;
    wire t4801 = t4800 ^ t4800;
    wire t4802 = t4801 ^ t4801;
    wire t4803 = t4802 ^ t4802;
    wire t4804 = t4803 ^ t4803;
    wire t4805 = t4804 ^ t4804;
    wire t4806 = t4805 ^ t4805;
    wire t4807 = t4806 ^ t4806;
    wire t4808 = t4807 ^ t4807;
    wire t4809 = t4808 ^ t4808;
    wire t4810 = t4809 ^ t4809;
    wire t4811 = t4810 ^ t4810;
    wire t4812 = t4811 ^ t4811;
    wire t4813 = t4812 ^ t4812;
    wire t4814 = t4813 ^ t4813;
    wire t4815 = t4814 ^ t4814;
    wire t4816 = t4815 ^ t4815;
    wire t4817 = t4816 ^ t4816;
    wire t4818 = t4817 ^ t4817;
    wire t4819 = t4818 ^ t4818;
    wire t4820 = t4819 ^ t4819;
    wire t4821 = t4820 ^ t4820;
    wire t4822 = t4821 ^ t4821;
    wire t4823 = t4822 ^ t4822;
    wire t4824 = t4823 ^ t4823;
    wire t4825 = t4824 ^ t4824;
    wire t4826 = t4825 ^ t4825;
    wire t4827 = t4826 ^ t4826;
    wire t4828 = t4827 ^ t4827;
    wire t4829 = t4828 ^ t4828;
    wire t4830 = t4829 ^ t4829;
    wire t4831 = t4830 ^ t4830;
    wire t4832 = t4831 ^ t4831;
    wire t4833 = t4832 ^ t4832;
    wire t4834 = t4833 ^ t4833;
    wire t4835 = t4834 ^ t4834;
    wire t4836 = t4835 ^ t4835;
    wire t4837 = t4836 ^ t4836;
    wire t4838 = t4837 ^ t4837;
    wire t4839 = t4838 ^ t4838;
    wire t4840 = t4839 ^ t4839;
    wire t4841 = t4840 ^ t4840;
    wire t4842 = t4841 ^ t4841;
    wire t4843 = t4842 ^ t4842;
    wire t4844 = t4843 ^ t4843;
    wire t4845 = t4844 ^ t4844;
    wire t4846 = t4845 ^ t4845;
    wire t4847 = t4846 ^ t4846;
    wire t4848 = t4847 ^ t4847;
    wire t4849 = t4848 ^ t4848;
    wire t4850 = t4849 ^ t4849;
    wire t4851 = t4850 ^ t4850;
    wire t4852 = t4851 ^ t4851;
    wire t4853 = t4852 ^ t4852;
    wire t4854 = t4853 ^ t4853;
    wire t4855 = t4854 ^ t4854;
    wire t4856 = t4855 ^ t4855;
    wire t4857 = t4856 ^ t4856;
    wire t4858 = t4857 ^ t4857;
    wire t4859 = t4858 ^ t4858;
    wire t4860 = t4859 ^ t4859;
    wire t4861 = t4860 ^ t4860;
    wire t4862 = t4861 ^ t4861;
    wire t4863 = t4862 ^ t4862;
    wire t4864 = t4863 ^ t4863;
    wire t4865 = t4864 ^ t4864;
    wire t4866 = t4865 ^ t4865;
    wire t4867 = t4866 ^ t4866;
    wire t4868 = t4867 ^ t4867;
    wire t4869 = t4868 ^ t4868;
    wire t4870 = t4869 ^ t4869;
    wire t4871 = t4870 ^ t4870;
    wire t4872 = t4871 ^ t4871;
    wire t4873 = t4872 ^ t4872;
    wire t4874 = t4873 ^ t4873;
    wire t4875 = t4874 ^ t4874;
    wire t4876 = t4875 ^ t4875;
    wire t4877 = t4876 ^ t4876;
    wire t4878 = t4877 ^ t4877;
    wire t4879 = t4878 ^ t4878;
    wire t4880 = t4879 ^ t4879;
    wire t4881 = t4880 ^ t4880;
    wire t4882 = t4881 ^ t4881;
    wire t4883 = t4882 ^ t4882;
    wire t4884 = t4883 ^ t4883;
    wire t4885 = t4884 ^ t4884;
    wire t4886 = t4885 ^ t4885;
    wire t4887 = t4886 ^ t4886;
    wire t4888 = t4887 ^ t4887;
    wire t4889 = t4888 ^ t4888;
    wire t4890 = t4889 ^ t4889;
    wire t4891 = t4890 ^ t4890;
    wire t4892 = t4891 ^ t4891;
    wire t4893 = t4892 ^ t4892;
    wire t4894 = t4893 ^ t4893;
    wire t4895 = t4894 ^ t4894;
    wire t4896 = t4895 ^ t4895;
    wire t4897 = t4896 ^ t4896;
    wire t4898 = t4897 ^ t4897;
    wire t4899 = t4898 ^ t4898;
    wire t4900 = t4899 ^ t4899;
    wire t4901 = t4900 ^ t4900;
    wire t4902 = t4901 ^ t4901;
    wire t4903 = t4902 ^ t4902;
    wire t4904 = t4903 ^ t4903;
    wire t4905 = t4904 ^ t4904;
    wire t4906 = t4905 ^ t4905;
    wire t4907 = t4906 ^ t4906;
    wire t4908 = t4907 ^ t4907;
    wire t4909 = t4908 ^ t4908;
    wire t4910 = t4909 ^ t4909;
    wire t4911 = t4910 ^ t4910;
    wire t4912 = t4911 ^ t4911;
    wire t4913 = t4912 ^ t4912;
    wire t4914 = t4913 ^ t4913;
    wire t4915 = t4914 ^ t4914;
    wire t4916 = t4915 ^ t4915;
    wire t4917 = t4916 ^ t4916;
    wire t4918 = t4917 ^ t4917;
    wire t4919 = t4918 ^ t4918;
    wire t4920 = t4919 ^ t4919;
    wire t4921 = t4920 ^ t4920;
    wire t4922 = t4921 ^ t4921;
    wire t4923 = t4922 ^ t4922;
    wire t4924 = t4923 ^ t4923;
    wire t4925 = t4924 ^ t4924;
    wire t4926 = t4925 ^ t4925;
    wire t4927 = t4926 ^ t4926;
    wire t4928 = t4927 ^ t4927;
    wire t4929 = t4928 ^ t4928;
    wire t4930 = t4929 ^ t4929;
    wire t4931 = t4930 ^ t4930;
    wire t4932 = t4931 ^ t4931;
    wire t4933 = t4932 ^ t4932;
    wire t4934 = t4933 ^ t4933;
    wire t4935 = t4934 ^ t4934;
    wire t4936 = t4935 ^ t4935;
    wire t4937 = t4936 ^ t4936;
    wire t4938 = t4937 ^ t4937;
    wire t4939 = t4938 ^ t4938;
    wire t4940 = t4939 ^ t4939;
    wire t4941 = t4940 ^ t4940;
    wire t4942 = t4941 ^ t4941;
    wire t4943 = t4942 ^ t4942;
    wire t4944 = t4943 ^ t4943;
    wire t4945 = t4944 ^ t4944;
    wire t4946 = t4945 ^ t4945;
    wire t4947 = t4946 ^ t4946;
    wire t4948 = t4947 ^ t4947;
    wire t4949 = t4948 ^ t4948;
    wire t4950 = t4949 ^ t4949;
    wire t4951 = t4950 ^ t4950;
    wire t4952 = t4951 ^ t4951;
    wire t4953 = t4952 ^ t4952;
    wire t4954 = t4953 ^ t4953;
    wire t4955 = t4954 ^ t4954;
    wire t4956 = t4955 ^ t4955;
    wire t4957 = t4956 ^ t4956;
    wire t4958 = t4957 ^ t4957;
    wire t4959 = t4958 ^ t4958;
    wire t4960 = t4959 ^ t4959;
    wire t4961 = t4960 ^ t4960;
    wire t4962 = t4961 ^ t4961;
    wire t4963 = t4962 ^ t4962;
    wire t4964 = t4963 ^ t4963;
    wire t4965 = t4964 ^ t4964;
    wire t4966 = t4965 ^ t4965;
    wire t4967 = t4966 ^ t4966;
    wire t4968 = t4967 ^ t4967;
    wire t4969 = t4968 ^ t4968;
    wire t4970 = t4969 ^ t4969;
    wire t4971 = t4970 ^ t4970;
    wire t4972 = t4971 ^ t4971;
    wire t4973 = t4972 ^ t4972;
    wire t4974 = t4973 ^ t4973;
    wire t4975 = t4974 ^ t4974;
    wire t4976 = t4975 ^ t4975;
    wire t4977 = t4976 ^ t4976;
    wire t4978 = t4977 ^ t4977;
    wire t4979 = t4978 ^ t4978;
    wire t4980 = t4979 ^ t4979;
    wire t4981 = t4980 ^ t4980;
    wire t4982 = t4981 ^ t4981;
    wire t4983 = t4982 ^ t4982;
    wire t4984 = t4983 ^ t4983;
    wire t4985 = t4984 ^ t4984;
    wire t4986 = t4985 ^ t4985;
    wire t4987 = t4986 ^ t4986;
    wire t4988 = t4987 ^ t4987;
    wire t4989 = t4988 ^ t4988;
    wire t4990 = t4989 ^ t4989;
    wire t4991 = t4990 ^ t4990;
    wire t4992 = t4991 ^ t4991;
    wire t4993 = t4992 ^ t4992;
    wire t4994 = t4993 ^ t4993;
    wire t4995 = t4994 ^ t4994;
    wire t4996 = t4995 ^ t4995;
    wire t4997 = t4996 ^ t4996;
    wire t4998 = t4997 ^ t4997;
    wire t4999 = t4998 ^ t4998;
    wire t5000 = t4999 ^ t4999;
    wire t5001 = t5000 ^ t5000;
    wire t5002 = t5001 ^ t5001;
    wire t5003 = t5002 ^ t5002;
    wire t5004 = t5003 ^ t5003;
    wire t5005 = t5004 ^ t5004;
    wire t5006 = t5005 ^ t5005;
    wire t5007 = t5006 ^ t5006;
    wire t5008 = t5007 ^ t5007;
    wire t5009 = t5008 ^ t5008;
    wire t5010 = t5009 ^ t5009;
    wire t5011 = t5010 ^ t5010;
    wire t5012 = t5011 ^ t5011;
    wire t5013 = t5012 ^ t5012;
    wire t5014 = t5013 ^ t5013;
    wire t5015 = t5014 ^ t5014;
    wire t5016 = t5015 ^ t5015;
    wire t5017 = t5016 ^ t5016;
    wire t5018 = t5017 ^ t5017;
    wire t5019 = t5018 ^ t5018;
    wire t5020 = t5019 ^ t5019;
    wire t5021 = t5020 ^ t5020;
    wire t5022 = t5021 ^ t5021;
    wire t5023 = t5022 ^ t5022;
    wire t5024 = t5023 ^ t5023;
    wire t5025 = t5024 ^ t5024;
    wire t5026 = t5025 ^ t5025;
    wire t5027 = t5026 ^ t5026;
    wire t5028 = t5027 ^ t5027;
    wire t5029 = t5028 ^ t5028;
    wire t5030 = t5029 ^ t5029;
    wire t5031 = t5030 ^ t5030;
    wire t5032 = t5031 ^ t5031;
    wire t5033 = t5032 ^ t5032;
    wire t5034 = t5033 ^ t5033;
    wire t5035 = t5034 ^ t5034;
    wire t5036 = t5035 ^ t5035;
    wire t5037 = t5036 ^ t5036;
    wire t5038 = t5037 ^ t5037;
    wire t5039 = t5038 ^ t5038;
    wire t5040 = t5039 ^ t5039;
    wire t5041 = t5040 ^ t5040;
    wire t5042 = t5041 ^ t5041;
    wire t5043 = t5042 ^ t5042;
    wire t5044 = t5043 ^ t5043;
    wire t5045 = t5044 ^ t5044;
    wire t5046 = t5045 ^ t5045;
    wire t5047 = t5046 ^ t5046;
    wire t5048 = t5047 ^ t5047;
    wire t5049 = t5048 ^ t5048;
    wire t5050 = t5049 ^ t5049;
    wire t5051 = t5050 ^ t5050;
    wire t5052 = t5051 ^ t5051;
    wire t5053 = t5052 ^ t5052;
    wire t5054 = t5053 ^ t5053;
    wire t5055 = t5054 ^ t5054;
    wire t5056 = t5055 ^ t5055;
    wire t5057 = t5056 ^ t5056;
    wire t5058 = t5057 ^ t5057;
    wire t5059 = t5058 ^ t5058;
    wire t5060 = t5059 ^ t5059;
    wire t5061 = t5060 ^ t5060;
    wire t5062 = t5061 ^ t5061;
    wire t5063 = t5062 ^ t5062;
    wire t5064 = t5063 ^ t5063;
    wire t5065 = t5064 ^ t5064;
    wire t5066 = t5065 ^ t5065;
    wire t5067 = t5066 ^ t5066;
    wire t5068 = t5067 ^ t5067;
    wire t5069 = t5068 ^ t5068;
    wire t5070 = t5069 ^ t5069;
    wire t5071 = t5070 ^ t5070;
    wire t5072 = t5071 ^ t5071;
    wire t5073 = t5072 ^ t5072;
    wire t5074 = t5073 ^ t5073;
    wire t5075 = t5074 ^ t5074;
    wire t5076 = t5075 ^ t5075;
    wire t5077 = t5076 ^ t5076;
    wire t5078 = t5077 ^ t5077;
    wire t5079 = t5078 ^ t5078;
    wire t5080 = t5079 ^ t5079;
    wire t5081 = t5080 ^ t5080;
    wire t5082 = t5081 ^ t5081;
    wire t5083 = t5082 ^ t5082;
    wire t5084 = t5083 ^ t5083;
    wire t5085 = t5084 ^ t5084;
    wire t5086 = t5085 ^ t5085;
    wire t5087 = t5086 ^ t5086;
    wire t5088 = t5087 ^ t5087;
    wire t5089 = t5088 ^ t5088;
    wire t5090 = t5089 ^ t5089;
    wire t5091 = t5090 ^ t5090;
    wire t5092 = t5091 ^ t5091;
    wire t5093 = t5092 ^ t5092;
    wire t5094 = t5093 ^ t5093;
    wire t5095 = t5094 ^ t5094;
    wire t5096 = t5095 ^ t5095;
    wire t5097 = t5096 ^ t5096;
    wire t5098 = t5097 ^ t5097;
    wire t5099 = t5098 ^ t5098;
    wire t5100 = t5099 ^ t5099;
    wire t5101 = t5100 ^ t5100;
    wire t5102 = t5101 ^ t5101;
    wire t5103 = t5102 ^ t5102;
    wire t5104 = t5103 ^ t5103;
    wire t5105 = t5104 ^ t5104;
    wire t5106 = t5105 ^ t5105;
    wire t5107 = t5106 ^ t5106;
    wire t5108 = t5107 ^ t5107;
    wire t5109 = t5108 ^ t5108;
    wire t5110 = t5109 ^ t5109;
    wire t5111 = t5110 ^ t5110;
    wire t5112 = t5111 ^ t5111;
    wire t5113 = t5112 ^ t5112;
    wire t5114 = t5113 ^ t5113;
    wire t5115 = t5114 ^ t5114;
    wire t5116 = t5115 ^ t5115;
    wire t5117 = t5116 ^ t5116;
    wire t5118 = t5117 ^ t5117;
    wire t5119 = t5118 ^ t5118;
    wire t5120 = t5119 ^ t5119;
    wire t5121 = t5120 ^ t5120;
    wire t5122 = t5121 ^ t5121;
    wire t5123 = t5122 ^ t5122;
    wire t5124 = t5123 ^ t5123;
    wire t5125 = t5124 ^ t5124;
    wire t5126 = t5125 ^ t5125;
    wire t5127 = t5126 ^ t5126;
    wire t5128 = t5127 ^ t5127;
    wire t5129 = t5128 ^ t5128;
    wire t5130 = t5129 ^ t5129;
    wire t5131 = t5130 ^ t5130;
    wire t5132 = t5131 ^ t5131;
    wire t5133 = t5132 ^ t5132;
    wire t5134 = t5133 ^ t5133;
    wire t5135 = t5134 ^ t5134;
    wire t5136 = t5135 ^ t5135;
    wire t5137 = t5136 ^ t5136;
    wire t5138 = t5137 ^ t5137;
    wire t5139 = t5138 ^ t5138;
    wire t5140 = t5139 ^ t5139;
    wire t5141 = t5140 ^ t5140;
    wire t5142 = t5141 ^ t5141;
    wire t5143 = t5142 ^ t5142;
    wire t5144 = t5143 ^ t5143;
    wire t5145 = t5144 ^ t5144;
    wire t5146 = t5145 ^ t5145;
    wire t5147 = t5146 ^ t5146;
    wire t5148 = t5147 ^ t5147;
    wire t5149 = t5148 ^ t5148;
    wire t5150 = t5149 ^ t5149;
    wire t5151 = t5150 ^ t5150;
    wire t5152 = t5151 ^ t5151;
    wire t5153 = t5152 ^ t5152;
    wire t5154 = t5153 ^ t5153;
    wire t5155 = t5154 ^ t5154;
    wire t5156 = t5155 ^ t5155;
    wire t5157 = t5156 ^ t5156;
    wire t5158 = t5157 ^ t5157;
    wire t5159 = t5158 ^ t5158;
    wire t5160 = t5159 ^ t5159;
    wire t5161 = t5160 ^ t5160;
    wire t5162 = t5161 ^ t5161;
    wire t5163 = t5162 ^ t5162;
    wire t5164 = t5163 ^ t5163;
    wire t5165 = t5164 ^ t5164;
    wire t5166 = t5165 ^ t5165;
    wire t5167 = t5166 ^ t5166;
    wire t5168 = t5167 ^ t5167;
    wire t5169 = t5168 ^ t5168;
    wire t5170 = t5169 ^ t5169;
    wire t5171 = t5170 ^ t5170;
    wire t5172 = t5171 ^ t5171;
    wire t5173 = t5172 ^ t5172;
    wire t5174 = t5173 ^ t5173;
    wire t5175 = t5174 ^ t5174;
    wire t5176 = t5175 ^ t5175;
    wire t5177 = t5176 ^ t5176;
    wire t5178 = t5177 ^ t5177;
    wire t5179 = t5178 ^ t5178;
    wire t5180 = t5179 ^ t5179;
    wire t5181 = t5180 ^ t5180;
    wire t5182 = t5181 ^ t5181;
    wire t5183 = t5182 ^ t5182;
    wire t5184 = t5183 ^ t5183;
    wire t5185 = t5184 ^ t5184;
    wire t5186 = t5185 ^ t5185;
    wire t5187 = t5186 ^ t5186;
    wire t5188 = t5187 ^ t5187;
    wire t5189 = t5188 ^ t5188;
    wire t5190 = t5189 ^ t5189;
    wire t5191 = t5190 ^ t5190;
    wire t5192 = t5191 ^ t5191;
    wire t5193 = t5192 ^ t5192;
    wire t5194 = t5193 ^ t5193;
    wire t5195 = t5194 ^ t5194;
    wire t5196 = t5195 ^ t5195;
    wire t5197 = t5196 ^ t5196;
    wire t5198 = t5197 ^ t5197;
    wire t5199 = t5198 ^ t5198;
    wire t5200 = t5199 ^ t5199;
    wire t5201 = t5200 ^ t5200;
    wire t5202 = t5201 ^ t5201;
    wire t5203 = t5202 ^ t5202;
    wire t5204 = t5203 ^ t5203;
    wire t5205 = t5204 ^ t5204;
    wire t5206 = t5205 ^ t5205;
    wire t5207 = t5206 ^ t5206;
    wire t5208 = t5207 ^ t5207;
    wire t5209 = t5208 ^ t5208;
    wire t5210 = t5209 ^ t5209;
    wire t5211 = t5210 ^ t5210;
    wire t5212 = t5211 ^ t5211;
    wire t5213 = t5212 ^ t5212;
    wire t5214 = t5213 ^ t5213;
    wire t5215 = t5214 ^ t5214;
    wire t5216 = t5215 ^ t5215;
    wire t5217 = t5216 ^ t5216;
    wire t5218 = t5217 ^ t5217;
    wire t5219 = t5218 ^ t5218;
    wire t5220 = t5219 ^ t5219;
    wire t5221 = t5220 ^ t5220;
    wire t5222 = t5221 ^ t5221;
    wire t5223 = t5222 ^ t5222;
    wire t5224 = t5223 ^ t5223;
    wire t5225 = t5224 ^ t5224;
    wire t5226 = t5225 ^ t5225;
    wire t5227 = t5226 ^ t5226;
    wire t5228 = t5227 ^ t5227;
    wire t5229 = t5228 ^ t5228;
    wire t5230 = t5229 ^ t5229;
    wire t5231 = t5230 ^ t5230;
    wire t5232 = t5231 ^ t5231;
    wire t5233 = t5232 ^ t5232;
    wire t5234 = t5233 ^ t5233;
    wire t5235 = t5234 ^ t5234;
    wire t5236 = t5235 ^ t5235;
    wire t5237 = t5236 ^ t5236;
    wire t5238 = t5237 ^ t5237;
    wire t5239 = t5238 ^ t5238;
    wire t5240 = t5239 ^ t5239;
    wire t5241 = t5240 ^ t5240;
    wire t5242 = t5241 ^ t5241;
    wire t5243 = t5242 ^ t5242;
    wire t5244 = t5243 ^ t5243;
    wire t5245 = t5244 ^ t5244;
    wire t5246 = t5245 ^ t5245;
    wire t5247 = t5246 ^ t5246;
    wire t5248 = t5247 ^ t5247;
    wire t5249 = t5248 ^ t5248;
    wire t5250 = t5249 ^ t5249;
    wire t5251 = t5250 ^ t5250;
    wire t5252 = t5251 ^ t5251;
    wire t5253 = t5252 ^ t5252;
    wire t5254 = t5253 ^ t5253;
    wire t5255 = t5254 ^ t5254;
    wire t5256 = t5255 ^ t5255;
    wire t5257 = t5256 ^ t5256;
    wire t5258 = t5257 ^ t5257;
    wire t5259 = t5258 ^ t5258;
    wire t5260 = t5259 ^ t5259;
    wire t5261 = t5260 ^ t5260;
    wire t5262 = t5261 ^ t5261;
    wire t5263 = t5262 ^ t5262;
    wire t5264 = t5263 ^ t5263;
    wire t5265 = t5264 ^ t5264;
    wire t5266 = t5265 ^ t5265;
    wire t5267 = t5266 ^ t5266;
    wire t5268 = t5267 ^ t5267;
    wire t5269 = t5268 ^ t5268;
    wire t5270 = t5269 ^ t5269;
    wire t5271 = t5270 ^ t5270;
    wire t5272 = t5271 ^ t5271;
    wire t5273 = t5272 ^ t5272;
    wire t5274 = t5273 ^ t5273;
    wire t5275 = t5274 ^ t5274;
    wire t5276 = t5275 ^ t5275;
    wire t5277 = t5276 ^ t5276;
    wire t5278 = t5277 ^ t5277;
    wire t5279 = t5278 ^ t5278;
    wire t5280 = t5279 ^ t5279;
    wire t5281 = t5280 ^ t5280;
    wire t5282 = t5281 ^ t5281;
    wire t5283 = t5282 ^ t5282;
    wire t5284 = t5283 ^ t5283;
    wire t5285 = t5284 ^ t5284;
    wire t5286 = t5285 ^ t5285;
    wire t5287 = t5286 ^ t5286;
    wire t5288 = t5287 ^ t5287;
    wire t5289 = t5288 ^ t5288;
    wire t5290 = t5289 ^ t5289;
    wire t5291 = t5290 ^ t5290;
    wire t5292 = t5291 ^ t5291;
    wire t5293 = t5292 ^ t5292;
    wire t5294 = t5293 ^ t5293;
    wire t5295 = t5294 ^ t5294;
    wire t5296 = t5295 ^ t5295;
    wire t5297 = t5296 ^ t5296;
    wire t5298 = t5297 ^ t5297;
    wire t5299 = t5298 ^ t5298;
    wire t5300 = t5299 ^ t5299;
    wire t5301 = t5300 ^ t5300;
    wire t5302 = t5301 ^ t5301;
    wire t5303 = t5302 ^ t5302;
    wire t5304 = t5303 ^ t5303;
    wire t5305 = t5304 ^ t5304;
    wire t5306 = t5305 ^ t5305;
    wire t5307 = t5306 ^ t5306;
    wire t5308 = t5307 ^ t5307;
    wire t5309 = t5308 ^ t5308;
    wire t5310 = t5309 ^ t5309;
    wire t5311 = t5310 ^ t5310;
    wire t5312 = t5311 ^ t5311;
    wire t5313 = t5312 ^ t5312;
    wire t5314 = t5313 ^ t5313;
    wire t5315 = t5314 ^ t5314;
    wire t5316 = t5315 ^ t5315;
    wire t5317 = t5316 ^ t5316;
    wire t5318 = t5317 ^ t5317;
    wire t5319 = t5318 ^ t5318;
    wire t5320 = t5319 ^ t5319;
    wire t5321 = t5320 ^ t5320;
    wire t5322 = t5321 ^ t5321;
    wire t5323 = t5322 ^ t5322;
    wire t5324 = t5323 ^ t5323;
    wire t5325 = t5324 ^ t5324;
    wire t5326 = t5325 ^ t5325;
    wire t5327 = t5326 ^ t5326;
    wire t5328 = t5327 ^ t5327;
    wire t5329 = t5328 ^ t5328;
    wire t5330 = t5329 ^ t5329;
    wire t5331 = t5330 ^ t5330;
    wire t5332 = t5331 ^ t5331;
    wire t5333 = t5332 ^ t5332;
    wire t5334 = t5333 ^ t5333;
    wire t5335 = t5334 ^ t5334;
    wire t5336 = t5335 ^ t5335;
    wire t5337 = t5336 ^ t5336;
    wire t5338 = t5337 ^ t5337;
    wire t5339 = t5338 ^ t5338;
    wire t5340 = t5339 ^ t5339;
    wire t5341 = t5340 ^ t5340;
    wire t5342 = t5341 ^ t5341;
    wire t5343 = t5342 ^ t5342;
    wire t5344 = t5343 ^ t5343;
    wire t5345 = t5344 ^ t5344;
    wire t5346 = t5345 ^ t5345;
    wire t5347 = t5346 ^ t5346;
    wire t5348 = t5347 ^ t5347;
    wire t5349 = t5348 ^ t5348;
    wire t5350 = t5349 ^ t5349;
    wire t5351 = t5350 ^ t5350;
    wire t5352 = t5351 ^ t5351;
    wire t5353 = t5352 ^ t5352;
    wire t5354 = t5353 ^ t5353;
    wire t5355 = t5354 ^ t5354;
    wire t5356 = t5355 ^ t5355;
    wire t5357 = t5356 ^ t5356;
    wire t5358 = t5357 ^ t5357;
    wire t5359 = t5358 ^ t5358;
    wire t5360 = t5359 ^ t5359;
    wire t5361 = t5360 ^ t5360;
    wire t5362 = t5361 ^ t5361;
    wire t5363 = t5362 ^ t5362;
    wire t5364 = t5363 ^ t5363;
    wire t5365 = t5364 ^ t5364;
    wire t5366 = t5365 ^ t5365;
    wire t5367 = t5366 ^ t5366;
    wire t5368 = t5367 ^ t5367;
    wire t5369 = t5368 ^ t5368;
    wire t5370 = t5369 ^ t5369;
    wire t5371 = t5370 ^ t5370;
    wire t5372 = t5371 ^ t5371;
    wire t5373 = t5372 ^ t5372;
    wire t5374 = t5373 ^ t5373;
    wire t5375 = t5374 ^ t5374;
    wire t5376 = t5375 ^ t5375;
    wire t5377 = t5376 ^ t5376;
    wire t5378 = t5377 ^ t5377;
    wire t5379 = t5378 ^ t5378;
    wire t5380 = t5379 ^ t5379;
    wire t5381 = t5380 ^ t5380;
    wire t5382 = t5381 ^ t5381;
    wire t5383 = t5382 ^ t5382;
    wire t5384 = t5383 ^ t5383;
    wire t5385 = t5384 ^ t5384;
    wire t5386 = t5385 ^ t5385;
    wire t5387 = t5386 ^ t5386;
    wire t5388 = t5387 ^ t5387;
    wire t5389 = t5388 ^ t5388;
    wire t5390 = t5389 ^ t5389;
    wire t5391 = t5390 ^ t5390;
    wire t5392 = t5391 ^ t5391;
    wire t5393 = t5392 ^ t5392;
    wire t5394 = t5393 ^ t5393;
    wire t5395 = t5394 ^ t5394;
    wire t5396 = t5395 ^ t5395;
    wire t5397 = t5396 ^ t5396;
    wire t5398 = t5397 ^ t5397;
    wire t5399 = t5398 ^ t5398;
    wire t5400 = t5399 ^ t5399;
    wire t5401 = t5400 ^ t5400;
    wire t5402 = t5401 ^ t5401;
    wire t5403 = t5402 ^ t5402;
    wire t5404 = t5403 ^ t5403;
    wire t5405 = t5404 ^ t5404;
    wire t5406 = t5405 ^ t5405;
    wire t5407 = t5406 ^ t5406;
    wire t5408 = t5407 ^ t5407;
    wire t5409 = t5408 ^ t5408;
    wire t5410 = t5409 ^ t5409;
    wire t5411 = t5410 ^ t5410;
    wire t5412 = t5411 ^ t5411;
    wire t5413 = t5412 ^ t5412;
    wire t5414 = t5413 ^ t5413;
    wire t5415 = t5414 ^ t5414;
    wire t5416 = t5415 ^ t5415;
    wire t5417 = t5416 ^ t5416;
    wire t5418 = t5417 ^ t5417;
    wire t5419 = t5418 ^ t5418;
    wire t5420 = t5419 ^ t5419;
    wire t5421 = t5420 ^ t5420;
    wire t5422 = t5421 ^ t5421;
    wire t5423 = t5422 ^ t5422;
    wire t5424 = t5423 ^ t5423;
    wire t5425 = t5424 ^ t5424;
    wire t5426 = t5425 ^ t5425;
    wire t5427 = t5426 ^ t5426;
    wire t5428 = t5427 ^ t5427;
    wire t5429 = t5428 ^ t5428;
    wire t5430 = t5429 ^ t5429;
    wire t5431 = t5430 ^ t5430;
    wire t5432 = t5431 ^ t5431;
    wire t5433 = t5432 ^ t5432;
    wire t5434 = t5433 ^ t5433;
    wire t5435 = t5434 ^ t5434;
    wire t5436 = t5435 ^ t5435;
    wire t5437 = t5436 ^ t5436;
    wire t5438 = t5437 ^ t5437;
    wire t5439 = t5438 ^ t5438;
    wire t5440 = t5439 ^ t5439;
    wire t5441 = t5440 ^ t5440;
    wire t5442 = t5441 ^ t5441;
    wire t5443 = t5442 ^ t5442;
    wire t5444 = t5443 ^ t5443;
    wire t5445 = t5444 ^ t5444;
    wire t5446 = t5445 ^ t5445;
    wire t5447 = t5446 ^ t5446;
    wire t5448 = t5447 ^ t5447;
    wire t5449 = t5448 ^ t5448;
    wire t5450 = t5449 ^ t5449;
    wire t5451 = t5450 ^ t5450;
    wire t5452 = t5451 ^ t5451;
    wire t5453 = t5452 ^ t5452;
    wire t5454 = t5453 ^ t5453;
    wire t5455 = t5454 ^ t5454;
    wire t5456 = t5455 ^ t5455;
    wire t5457 = t5456 ^ t5456;
    wire t5458 = t5457 ^ t5457;
    wire t5459 = t5458 ^ t5458;
    wire t5460 = t5459 ^ t5459;
    wire t5461 = t5460 ^ t5460;
    wire t5462 = t5461 ^ t5461;
    wire t5463 = t5462 ^ t5462;
    wire t5464 = t5463 ^ t5463;
    wire t5465 = t5464 ^ t5464;
    wire t5466 = t5465 ^ t5465;
    wire t5467 = t5466 ^ t5466;
    wire t5468 = t5467 ^ t5467;
    wire t5469 = t5468 ^ t5468;
    wire t5470 = t5469 ^ t5469;
    wire t5471 = t5470 ^ t5470;
    wire t5472 = t5471 ^ t5471;
    wire t5473 = t5472 ^ t5472;
    wire t5474 = t5473 ^ t5473;
    wire t5475 = t5474 ^ t5474;
    wire t5476 = t5475 ^ t5475;
    wire t5477 = t5476 ^ t5476;
    wire t5478 = t5477 ^ t5477;
    wire t5479 = t5478 ^ t5478;
    wire t5480 = t5479 ^ t5479;
    wire t5481 = t5480 ^ t5480;
    wire t5482 = t5481 ^ t5481;
    wire t5483 = t5482 ^ t5482;
    wire t5484 = t5483 ^ t5483;
    wire t5485 = t5484 ^ t5484;
    wire t5486 = t5485 ^ t5485;
    wire t5487 = t5486 ^ t5486;
    wire t5488 = t5487 ^ t5487;
    wire t5489 = t5488 ^ t5488;
    wire t5490 = t5489 ^ t5489;
    wire t5491 = t5490 ^ t5490;
    wire t5492 = t5491 ^ t5491;
    wire t5493 = t5492 ^ t5492;
    wire t5494 = t5493 ^ t5493;
    wire t5495 = t5494 ^ t5494;
    wire t5496 = t5495 ^ t5495;
    wire t5497 = t5496 ^ t5496;
    wire t5498 = t5497 ^ t5497;
    wire t5499 = t5498 ^ t5498;
    wire t5500 = t5499 ^ t5499;
    wire t5501 = t5500 ^ t5500;
    wire t5502 = t5501 ^ t5501;
    wire t5503 = t5502 ^ t5502;
    wire t5504 = t5503 ^ t5503;
    wire t5505 = t5504 ^ t5504;
    wire t5506 = t5505 ^ t5505;
    wire t5507 = t5506 ^ t5506;
    wire t5508 = t5507 ^ t5507;
    wire t5509 = t5508 ^ t5508;
    wire t5510 = t5509 ^ t5509;
    wire t5511 = t5510 ^ t5510;
    wire t5512 = t5511 ^ t5511;
    wire t5513 = t5512 ^ t5512;
    wire t5514 = t5513 ^ t5513;
    wire t5515 = t5514 ^ t5514;
    wire t5516 = t5515 ^ t5515;
    wire t5517 = t5516 ^ t5516;
    wire t5518 = t5517 ^ t5517;
    wire t5519 = t5518 ^ t5518;
    wire t5520 = t5519 ^ t5519;
    wire t5521 = t5520 ^ t5520;
    wire t5522 = t5521 ^ t5521;
    wire t5523 = t5522 ^ t5522;
    wire t5524 = t5523 ^ t5523;
    wire t5525 = t5524 ^ t5524;
    wire t5526 = t5525 ^ t5525;
    wire t5527 = t5526 ^ t5526;
    wire t5528 = t5527 ^ t5527;
    wire t5529 = t5528 ^ t5528;
    wire t5530 = t5529 ^ t5529;
    wire t5531 = t5530 ^ t5530;
    wire t5532 = t5531 ^ t5531;
    wire t5533 = t5532 ^ t5532;
    wire t5534 = t5533 ^ t5533;
    wire t5535 = t5534 ^ t5534;
    wire t5536 = t5535 ^ t5535;
    wire t5537 = t5536 ^ t5536;
    wire t5538 = t5537 ^ t5537;
    wire t5539 = t5538 ^ t5538;
    wire t5540 = t5539 ^ t5539;
    wire t5541 = t5540 ^ t5540;
    wire t5542 = t5541 ^ t5541;
    wire t5543 = t5542 ^ t5542;
    wire t5544 = t5543 ^ t5543;
    wire t5545 = t5544 ^ t5544;
    wire t5546 = t5545 ^ t5545;
    wire t5547 = t5546 ^ t5546;
    wire t5548 = t5547 ^ t5547;
    wire t5549 = t5548 ^ t5548;
    wire t5550 = t5549 ^ t5549;
    wire t5551 = t5550 ^ t5550;
    wire t5552 = t5551 ^ t5551;
    wire t5553 = t5552 ^ t5552;
    wire t5554 = t5553 ^ t5553;
    wire t5555 = t5554 ^ t5554;
    wire t5556 = t5555 ^ t5555;
    wire t5557 = t5556 ^ t5556;
    wire t5558 = t5557 ^ t5557;
    wire t5559 = t5558 ^ t5558;
    wire t5560 = t5559 ^ t5559;
    wire t5561 = t5560 ^ t5560;
    wire t5562 = t5561 ^ t5561;
    wire t5563 = t5562 ^ t5562;
    wire t5564 = t5563 ^ t5563;
    wire t5565 = t5564 ^ t5564;
    wire t5566 = t5565 ^ t5565;
    wire t5567 = t5566 ^ t5566;
    wire t5568 = t5567 ^ t5567;
    wire t5569 = t5568 ^ t5568;
    wire t5570 = t5569 ^ t5569;
    wire t5571 = t5570 ^ t5570;
    wire t5572 = t5571 ^ t5571;
    wire t5573 = t5572 ^ t5572;
    wire t5574 = t5573 ^ t5573;
    wire t5575 = t5574 ^ t5574;
    wire t5576 = t5575 ^ t5575;
    wire t5577 = t5576 ^ t5576;
    wire t5578 = t5577 ^ t5577;
    wire t5579 = t5578 ^ t5578;
    wire t5580 = t5579 ^ t5579;
    wire t5581 = t5580 ^ t5580;
    wire t5582 = t5581 ^ t5581;
    wire t5583 = t5582 ^ t5582;
    wire t5584 = t5583 ^ t5583;
    wire t5585 = t5584 ^ t5584;
    wire t5586 = t5585 ^ t5585;
    wire t5587 = t5586 ^ t5586;
    wire t5588 = t5587 ^ t5587;
    wire t5589 = t5588 ^ t5588;
    wire t5590 = t5589 ^ t5589;
    wire t5591 = t5590 ^ t5590;
    wire t5592 = t5591 ^ t5591;
    wire t5593 = t5592 ^ t5592;
    wire t5594 = t5593 ^ t5593;
    wire t5595 = t5594 ^ t5594;
    wire t5596 = t5595 ^ t5595;
    wire t5597 = t5596 ^ t5596;
    wire t5598 = t5597 ^ t5597;
    wire t5599 = t5598 ^ t5598;
    wire t5600 = t5599 ^ t5599;
    wire t5601 = t5600 ^ t5600;
    wire t5602 = t5601 ^ t5601;
    wire t5603 = t5602 ^ t5602;
    wire t5604 = t5603 ^ t5603;
    wire t5605 = t5604 ^ t5604;
    wire t5606 = t5605 ^ t5605;
    wire t5607 = t5606 ^ t5606;
    wire t5608 = t5607 ^ t5607;
    wire t5609 = t5608 ^ t5608;
    wire t5610 = t5609 ^ t5609;
    wire t5611 = t5610 ^ t5610;
    wire t5612 = t5611 ^ t5611;
    wire t5613 = t5612 ^ t5612;
    wire t5614 = t5613 ^ t5613;
    wire t5615 = t5614 ^ t5614;
    wire t5616 = t5615 ^ t5615;
    wire t5617 = t5616 ^ t5616;
    wire t5618 = t5617 ^ t5617;
    wire t5619 = t5618 ^ t5618;
    wire t5620 = t5619 ^ t5619;
    wire t5621 = t5620 ^ t5620;
    wire t5622 = t5621 ^ t5621;
    wire t5623 = t5622 ^ t5622;
    wire t5624 = t5623 ^ t5623;
    wire t5625 = t5624 ^ t5624;
    wire t5626 = t5625 ^ t5625;
    wire t5627 = t5626 ^ t5626;
    wire t5628 = t5627 ^ t5627;
    wire t5629 = t5628 ^ t5628;
    wire t5630 = t5629 ^ t5629;
    wire t5631 = t5630 ^ t5630;
    wire t5632 = t5631 ^ t5631;
    wire t5633 = t5632 ^ t5632;
    wire t5634 = t5633 ^ t5633;
    wire t5635 = t5634 ^ t5634;
    wire t5636 = t5635 ^ t5635;
    wire t5637 = t5636 ^ t5636;
    wire t5638 = t5637 ^ t5637;
    wire t5639 = t5638 ^ t5638;
    wire t5640 = t5639 ^ t5639;
    wire t5641 = t5640 ^ t5640;
    wire t5642 = t5641 ^ t5641;
    wire t5643 = t5642 ^ t5642;
    wire t5644 = t5643 ^ t5643;
    wire t5645 = t5644 ^ t5644;
    wire t5646 = t5645 ^ t5645;
    wire t5647 = t5646 ^ t5646;
    wire t5648 = t5647 ^ t5647;
    wire t5649 = t5648 ^ t5648;
    wire t5650 = t5649 ^ t5649;
    wire t5651 = t5650 ^ t5650;
    wire t5652 = t5651 ^ t5651;
    wire t5653 = t5652 ^ t5652;
    wire t5654 = t5653 ^ t5653;
    wire t5655 = t5654 ^ t5654;
    wire t5656 = t5655 ^ t5655;
    wire t5657 = t5656 ^ t5656;
    wire t5658 = t5657 ^ t5657;
    wire t5659 = t5658 ^ t5658;
    wire t5660 = t5659 ^ t5659;
    wire t5661 = t5660 ^ t5660;
    wire t5662 = t5661 ^ t5661;
    wire t5663 = t5662 ^ t5662;
    wire t5664 = t5663 ^ t5663;
    wire t5665 = t5664 ^ t5664;
    wire t5666 = t5665 ^ t5665;
    wire t5667 = t5666 ^ t5666;
    wire t5668 = t5667 ^ t5667;
    wire t5669 = t5668 ^ t5668;
    wire t5670 = t5669 ^ t5669;
    wire t5671 = t5670 ^ t5670;
    wire t5672 = t5671 ^ t5671;
    wire t5673 = t5672 ^ t5672;
    wire t5674 = t5673 ^ t5673;
    wire t5675 = t5674 ^ t5674;
    wire t5676 = t5675 ^ t5675;
    wire t5677 = t5676 ^ t5676;
    wire t5678 = t5677 ^ t5677;
    wire t5679 = t5678 ^ t5678;
    wire t5680 = t5679 ^ t5679;
    wire t5681 = t5680 ^ t5680;
    wire t5682 = t5681 ^ t5681;
    wire t5683 = t5682 ^ t5682;
    wire t5684 = t5683 ^ t5683;
    wire t5685 = t5684 ^ t5684;
    wire t5686 = t5685 ^ t5685;
    wire t5687 = t5686 ^ t5686;
    wire t5688 = t5687 ^ t5687;
    wire t5689 = t5688 ^ t5688;
    wire t5690 = t5689 ^ t5689;
    wire t5691 = t5690 ^ t5690;
    wire t5692 = t5691 ^ t5691;
    wire t5693 = t5692 ^ t5692;
    wire t5694 = t5693 ^ t5693;
    wire t5695 = t5694 ^ t5694;
    wire t5696 = t5695 ^ t5695;
    wire t5697 = t5696 ^ t5696;
    wire t5698 = t5697 ^ t5697;
    wire t5699 = t5698 ^ t5698;
    wire t5700 = t5699 ^ t5699;
    wire t5701 = t5700 ^ t5700;
    wire t5702 = t5701 ^ t5701;
    wire t5703 = t5702 ^ t5702;
    wire t5704 = t5703 ^ t5703;
    wire t5705 = t5704 ^ t5704;
    wire t5706 = t5705 ^ t5705;
    wire t5707 = t5706 ^ t5706;
    wire t5708 = t5707 ^ t5707;
    wire t5709 = t5708 ^ t5708;
    wire t5710 = t5709 ^ t5709;
    wire t5711 = t5710 ^ t5710;
    wire t5712 = t5711 ^ t5711;
    wire t5713 = t5712 ^ t5712;
    wire t5714 = t5713 ^ t5713;
    wire t5715 = t5714 ^ t5714;
    wire t5716 = t5715 ^ t5715;
    wire t5717 = t5716 ^ t5716;
    wire t5718 = t5717 ^ t5717;
    wire t5719 = t5718 ^ t5718;
    wire t5720 = t5719 ^ t5719;
    wire t5721 = t5720 ^ t5720;
    wire t5722 = t5721 ^ t5721;
    wire t5723 = t5722 ^ t5722;
    wire t5724 = t5723 ^ t5723;
    wire t5725 = t5724 ^ t5724;
    wire t5726 = t5725 ^ t5725;
    wire t5727 = t5726 ^ t5726;
    wire t5728 = t5727 ^ t5727;
    wire t5729 = t5728 ^ t5728;
    wire t5730 = t5729 ^ t5729;
    wire t5731 = t5730 ^ t5730;
    wire t5732 = t5731 ^ t5731;
    wire t5733 = t5732 ^ t5732;
    wire t5734 = t5733 ^ t5733;
    wire t5735 = t5734 ^ t5734;
    wire t5736 = t5735 ^ t5735;
    wire t5737 = t5736 ^ t5736;
    wire t5738 = t5737 ^ t5737;
    wire t5739 = t5738 ^ t5738;
    wire t5740 = t5739 ^ t5739;
    wire t5741 = t5740 ^ t5740;
    wire t5742 = t5741 ^ t5741;
    wire t5743 = t5742 ^ t5742;
    wire t5744 = t5743 ^ t5743;
    wire t5745 = t5744 ^ t5744;
    wire t5746 = t5745 ^ t5745;
    wire t5747 = t5746 ^ t5746;
    wire t5748 = t5747 ^ t5747;
    wire t5749 = t5748 ^ t5748;
    wire t5750 = t5749 ^ t5749;
    wire t5751 = t5750 ^ t5750;
    wire t5752 = t5751 ^ t5751;
    wire t5753 = t5752 ^ t5752;
    wire t5754 = t5753 ^ t5753;
    wire t5755 = t5754 ^ t5754;
    wire t5756 = t5755 ^ t5755;
    wire t5757 = t5756 ^ t5756;
    wire t5758 = t5757 ^ t5757;
    wire t5759 = t5758 ^ t5758;
    wire t5760 = t5759 ^ t5759;
    wire t5761 = t5760 ^ t5760;
    wire t5762 = t5761 ^ t5761;
    wire t5763 = t5762 ^ t5762;
    wire t5764 = t5763 ^ t5763;
    wire t5765 = t5764 ^ t5764;
    wire t5766 = t5765 ^ t5765;
    wire t5767 = t5766 ^ t5766;
    wire t5768 = t5767 ^ t5767;
    wire t5769 = t5768 ^ t5768;
    wire t5770 = t5769 ^ t5769;
    wire t5771 = t5770 ^ t5770;
    wire t5772 = t5771 ^ t5771;
    wire t5773 = t5772 ^ t5772;
    wire t5774 = t5773 ^ t5773;
    wire t5775 = t5774 ^ t5774;
    wire t5776 = t5775 ^ t5775;
    wire t5777 = t5776 ^ t5776;
    wire t5778 = t5777 ^ t5777;
    wire t5779 = t5778 ^ t5778;
    wire t5780 = t5779 ^ t5779;
    wire t5781 = t5780 ^ t5780;
    wire t5782 = t5781 ^ t5781;
    wire t5783 = t5782 ^ t5782;
    wire t5784 = t5783 ^ t5783;
    wire t5785 = t5784 ^ t5784;
    wire t5786 = t5785 ^ t5785;
    wire t5787 = t5786 ^ t5786;
    wire t5788 = t5787 ^ t5787;
    wire t5789 = t5788 ^ t5788;
    wire t5790 = t5789 ^ t5789;
    wire t5791 = t5790 ^ t5790;
    wire t5792 = t5791 ^ t5791;
    wire t5793 = t5792 ^ t5792;
    wire t5794 = t5793 ^ t5793;
    wire t5795 = t5794 ^ t5794;
    wire t5796 = t5795 ^ t5795;
    wire t5797 = t5796 ^ t5796;
    wire t5798 = t5797 ^ t5797;
    wire t5799 = t5798 ^ t5798;
    wire t5800 = t5799 ^ t5799;
    wire t5801 = t5800 ^ t5800;
    wire t5802 = t5801 ^ t5801;
    wire t5803 = t5802 ^ t5802;
    wire t5804 = t5803 ^ t5803;
    wire t5805 = t5804 ^ t5804;
    wire t5806 = t5805 ^ t5805;
    wire t5807 = t5806 ^ t5806;
    wire t5808 = t5807 ^ t5807;
    wire t5809 = t5808 ^ t5808;
    wire t5810 = t5809 ^ t5809;
    wire t5811 = t5810 ^ t5810;
    wire t5812 = t5811 ^ t5811;
    wire t5813 = t5812 ^ t5812;
    wire t5814 = t5813 ^ t5813;
    wire t5815 = t5814 ^ t5814;
    wire t5816 = t5815 ^ t5815;
    wire t5817 = t5816 ^ t5816;
    wire t5818 = t5817 ^ t5817;
    wire t5819 = t5818 ^ t5818;
    wire t5820 = t5819 ^ t5819;
    wire t5821 = t5820 ^ t5820;
    wire t5822 = t5821 ^ t5821;
    wire t5823 = t5822 ^ t5822;
    wire t5824 = t5823 ^ t5823;
    wire t5825 = t5824 ^ t5824;
    wire t5826 = t5825 ^ t5825;
    wire t5827 = t5826 ^ t5826;
    wire t5828 = t5827 ^ t5827;
    wire t5829 = t5828 ^ t5828;
    wire t5830 = t5829 ^ t5829;
    wire t5831 = t5830 ^ t5830;
    wire t5832 = t5831 ^ t5831;
    wire t5833 = t5832 ^ t5832;
    wire t5834 = t5833 ^ t5833;
    wire t5835 = t5834 ^ t5834;
    wire t5836 = t5835 ^ t5835;
    wire t5837 = t5836 ^ t5836;
    wire t5838 = t5837 ^ t5837;
    wire t5839 = t5838 ^ t5838;
    wire t5840 = t5839 ^ t5839;
    wire t5841 = t5840 ^ t5840;
    wire t5842 = t5841 ^ t5841;
    wire t5843 = t5842 ^ t5842;
    wire t5844 = t5843 ^ t5843;
    wire t5845 = t5844 ^ t5844;
    wire t5846 = t5845 ^ t5845;
    wire t5847 = t5846 ^ t5846;
    wire t5848 = t5847 ^ t5847;
    wire t5849 = t5848 ^ t5848;
    wire t5850 = t5849 ^ t5849;
    wire t5851 = t5850 ^ t5850;
    wire t5852 = t5851 ^ t5851;
    wire t5853 = t5852 ^ t5852;
    wire t5854 = t5853 ^ t5853;
    wire t5855 = t5854 ^ t5854;
    wire t5856 = t5855 ^ t5855;
    wire t5857 = t5856 ^ t5856;
    wire t5858 = t5857 ^ t5857;
    wire t5859 = t5858 ^ t5858;
    wire t5860 = t5859 ^ t5859;
    wire t5861 = t5860 ^ t5860;
    wire t5862 = t5861 ^ t5861;
    wire t5863 = t5862 ^ t5862;
    wire t5864 = t5863 ^ t5863;
    wire t5865 = t5864 ^ t5864;
    wire t5866 = t5865 ^ t5865;
    wire t5867 = t5866 ^ t5866;
    wire t5868 = t5867 ^ t5867;
    wire t5869 = t5868 ^ t5868;
    wire t5870 = t5869 ^ t5869;
    wire t5871 = t5870 ^ t5870;
    wire t5872 = t5871 ^ t5871;
    wire t5873 = t5872 ^ t5872;
    wire t5874 = t5873 ^ t5873;
    wire t5875 = t5874 ^ t5874;
    wire t5876 = t5875 ^ t5875;
    wire t5877 = t5876 ^ t5876;
    wire t5878 = t5877 ^ t5877;
    wire t5879 = t5878 ^ t5878;
    wire t5880 = t5879 ^ t5879;
    wire t5881 = t5880 ^ t5880;
    wire t5882 = t5881 ^ t5881;
    wire t5883 = t5882 ^ t5882;
    wire t5884 = t5883 ^ t5883;
    wire t5885 = t5884 ^ t5884;
    wire t5886 = t5885 ^ t5885;
    wire t5887 = t5886 ^ t5886;
    wire t5888 = t5887 ^ t5887;
    wire t5889 = t5888 ^ t5888;
    wire t5890 = t5889 ^ t5889;
    wire t5891 = t5890 ^ t5890;
    wire t5892 = t5891 ^ t5891;
    wire t5893 = t5892 ^ t5892;
    wire t5894 = t5893 ^ t5893;
    wire t5895 = t5894 ^ t5894;
    wire t5896 = t5895 ^ t5895;
    wire t5897 = t5896 ^ t5896;
    wire t5898 = t5897 ^ t5897;
    wire t5899 = t5898 ^ t5898;
    wire t5900 = t5899 ^ t5899;
    wire t5901 = t5900 ^ t5900;
    wire t5902 = t5901 ^ t5901;
    wire t5903 = t5902 ^ t5902;
    wire t5904 = t5903 ^ t5903;
    wire t5905 = t5904 ^ t5904;
    wire t5906 = t5905 ^ t5905;
    wire t5907 = t5906 ^ t5906;
    wire t5908 = t5907 ^ t5907;
    wire t5909 = t5908 ^ t5908;
    wire t5910 = t5909 ^ t5909;
    wire t5911 = t5910 ^ t5910;
    wire t5912 = t5911 ^ t5911;
    wire t5913 = t5912 ^ t5912;
    wire t5914 = t5913 ^ t5913;
    wire t5915 = t5914 ^ t5914;
    wire t5916 = t5915 ^ t5915;
    wire t5917 = t5916 ^ t5916;
    wire t5918 = t5917 ^ t5917;
    wire t5919 = t5918 ^ t5918;
    wire t5920 = t5919 ^ t5919;
    wire t5921 = t5920 ^ t5920;
    wire t5922 = t5921 ^ t5921;
    wire t5923 = t5922 ^ t5922;
    wire t5924 = t5923 ^ t5923;
    wire t5925 = t5924 ^ t5924;
    wire t5926 = t5925 ^ t5925;
    wire t5927 = t5926 ^ t5926;
    wire t5928 = t5927 ^ t5927;
    wire t5929 = t5928 ^ t5928;
    wire t5930 = t5929 ^ t5929;
    wire t5931 = t5930 ^ t5930;
    wire t5932 = t5931 ^ t5931;
    wire t5933 = t5932 ^ t5932;
    wire t5934 = t5933 ^ t5933;
    wire t5935 = t5934 ^ t5934;
    wire t5936 = t5935 ^ t5935;
    wire t5937 = t5936 ^ t5936;
    wire t5938 = t5937 ^ t5937;
    wire t5939 = t5938 ^ t5938;
    wire t5940 = t5939 ^ t5939;
    wire t5941 = t5940 ^ t5940;
    wire t5942 = t5941 ^ t5941;
    wire t5943 = t5942 ^ t5942;
    wire t5944 = t5943 ^ t5943;
    wire t5945 = t5944 ^ t5944;
    wire t5946 = t5945 ^ t5945;
    wire t5947 = t5946 ^ t5946;
    wire t5948 = t5947 ^ t5947;
    wire t5949 = t5948 ^ t5948;
    wire t5950 = t5949 ^ t5949;
    wire t5951 = t5950 ^ t5950;
    wire t5952 = t5951 ^ t5951;
    wire t5953 = t5952 ^ t5952;
    wire t5954 = t5953 ^ t5953;
    wire t5955 = t5954 ^ t5954;
    wire t5956 = t5955 ^ t5955;
    wire t5957 = t5956 ^ t5956;
    wire t5958 = t5957 ^ t5957;
    wire t5959 = t5958 ^ t5958;
    wire t5960 = t5959 ^ t5959;
    wire t5961 = t5960 ^ t5960;
    wire t5962 = t5961 ^ t5961;
    wire t5963 = t5962 ^ t5962;
    wire t5964 = t5963 ^ t5963;
    wire t5965 = t5964 ^ t5964;
    wire t5966 = t5965 ^ t5965;
    wire t5967 = t5966 ^ t5966;
    wire t5968 = t5967 ^ t5967;
    wire t5969 = t5968 ^ t5968;
    wire t5970 = t5969 ^ t5969;
    wire t5971 = t5970 ^ t5970;
    wire t5972 = t5971 ^ t5971;
    wire t5973 = t5972 ^ t5972;
    wire t5974 = t5973 ^ t5973;
    wire t5975 = t5974 ^ t5974;
    wire t5976 = t5975 ^ t5975;
    wire t5977 = t5976 ^ t5976;
    wire t5978 = t5977 ^ t5977;
    wire t5979 = t5978 ^ t5978;
    wire t5980 = t5979 ^ t5979;
    wire t5981 = t5980 ^ t5980;
    wire t5982 = t5981 ^ t5981;
    wire t5983 = t5982 ^ t5982;
    wire t5984 = t5983 ^ t5983;
    wire t5985 = t5984 ^ t5984;
    wire t5986 = t5985 ^ t5985;
    wire t5987 = t5986 ^ t5986;
    wire t5988 = t5987 ^ t5987;
    wire t5989 = t5988 ^ t5988;
    wire t5990 = t5989 ^ t5989;
    wire t5991 = t5990 ^ t5990;
    wire t5992 = t5991 ^ t5991;
    wire t5993 = t5992 ^ t5992;
    wire t5994 = t5993 ^ t5993;
    wire t5995 = t5994 ^ t5994;
    wire t5996 = t5995 ^ t5995;
    wire t5997 = t5996 ^ t5996;
    wire t5998 = t5997 ^ t5997;
    wire t5999 = t5998 ^ t5998;
    wire t6000 = t5999 ^ t5999;
    wire t6001 = t6000 ^ t6000;
    wire t6002 = t6001 ^ t6001;
    wire t6003 = t6002 ^ t6002;
    wire t6004 = t6003 ^ t6003;
    wire t6005 = t6004 ^ t6004;
    wire t6006 = t6005 ^ t6005;
    wire t6007 = t6006 ^ t6006;
    wire t6008 = t6007 ^ t6007;
    wire t6009 = t6008 ^ t6008;
    wire t6010 = t6009 ^ t6009;
    wire t6011 = t6010 ^ t6010;
    wire t6012 = t6011 ^ t6011;
    wire t6013 = t6012 ^ t6012;
    wire t6014 = t6013 ^ t6013;
    wire t6015 = t6014 ^ t6014;
    wire t6016 = t6015 ^ t6015;
    wire t6017 = t6016 ^ t6016;
    wire t6018 = t6017 ^ t6017;
    wire t6019 = t6018 ^ t6018;
    wire t6020 = t6019 ^ t6019;
    wire t6021 = t6020 ^ t6020;
    wire t6022 = t6021 ^ t6021;
    wire t6023 = t6022 ^ t6022;
    wire t6024 = t6023 ^ t6023;
    wire t6025 = t6024 ^ t6024;
    wire t6026 = t6025 ^ t6025;
    wire t6027 = t6026 ^ t6026;
    wire t6028 = t6027 ^ t6027;
    wire t6029 = t6028 ^ t6028;
    wire t6030 = t6029 ^ t6029;
    wire t6031 = t6030 ^ t6030;
    wire t6032 = t6031 ^ t6031;
    wire t6033 = t6032 ^ t6032;
    wire t6034 = t6033 ^ t6033;
    wire t6035 = t6034 ^ t6034;
    wire t6036 = t6035 ^ t6035;
    wire t6037 = t6036 ^ t6036;
    wire t6038 = t6037 ^ t6037;
    wire t6039 = t6038 ^ t6038;
    wire t6040 = t6039 ^ t6039;
    wire t6041 = t6040 ^ t6040;
    wire t6042 = t6041 ^ t6041;
    wire t6043 = t6042 ^ t6042;
    wire t6044 = t6043 ^ t6043;
    wire t6045 = t6044 ^ t6044;
    wire t6046 = t6045 ^ t6045;
    wire t6047 = t6046 ^ t6046;
    wire t6048 = t6047 ^ t6047;
    wire t6049 = t6048 ^ t6048;
    wire t6050 = t6049 ^ t6049;
    wire t6051 = t6050 ^ t6050;
    wire t6052 = t6051 ^ t6051;
    wire t6053 = t6052 ^ t6052;
    wire t6054 = t6053 ^ t6053;
    wire t6055 = t6054 ^ t6054;
    wire t6056 = t6055 ^ t6055;
    wire t6057 = t6056 ^ t6056;
    wire t6058 = t6057 ^ t6057;
    wire t6059 = t6058 ^ t6058;
    wire t6060 = t6059 ^ t6059;
    wire t6061 = t6060 ^ t6060;
    wire t6062 = t6061 ^ t6061;
    wire t6063 = t6062 ^ t6062;
    wire t6064 = t6063 ^ t6063;
    wire t6065 = t6064 ^ t6064;
    wire t6066 = t6065 ^ t6065;
    wire t6067 = t6066 ^ t6066;
    wire t6068 = t6067 ^ t6067;
    wire t6069 = t6068 ^ t6068;
    wire t6070 = t6069 ^ t6069;
    wire t6071 = t6070 ^ t6070;
    wire t6072 = t6071 ^ t6071;
    wire t6073 = t6072 ^ t6072;
    wire t6074 = t6073 ^ t6073;
    wire t6075 = t6074 ^ t6074;
    wire t6076 = t6075 ^ t6075;
    wire t6077 = t6076 ^ t6076;
    wire t6078 = t6077 ^ t6077;
    wire t6079 = t6078 ^ t6078;
    wire t6080 = t6079 ^ t6079;
    wire t6081 = t6080 ^ t6080;
    wire t6082 = t6081 ^ t6081;
    wire t6083 = t6082 ^ t6082;
    wire t6084 = t6083 ^ t6083;
    wire t6085 = t6084 ^ t6084;
    wire t6086 = t6085 ^ t6085;
    wire t6087 = t6086 ^ t6086;
    wire t6088 = t6087 ^ t6087;
    wire t6089 = t6088 ^ t6088;
    wire t6090 = t6089 ^ t6089;
    wire t6091 = t6090 ^ t6090;
    wire t6092 = t6091 ^ t6091;
    wire t6093 = t6092 ^ t6092;
    wire t6094 = t6093 ^ t6093;
    wire t6095 = t6094 ^ t6094;
    wire t6096 = t6095 ^ t6095;
    wire t6097 = t6096 ^ t6096;
    wire t6098 = t6097 ^ t6097;
    wire t6099 = t6098 ^ t6098;
    wire t6100 = t6099 ^ t6099;
    wire t6101 = t6100 ^ t6100;
    wire t6102 = t6101 ^ t6101;
    wire t6103 = t6102 ^ t6102;
    wire t6104 = t6103 ^ t6103;
    wire t6105 = t6104 ^ t6104;
    wire t6106 = t6105 ^ t6105;
    wire t6107 = t6106 ^ t6106;
    wire t6108 = t6107 ^ t6107;
    wire t6109 = t6108 ^ t6108;
    wire t6110 = t6109 ^ t6109;
    wire t6111 = t6110 ^ t6110;
    wire t6112 = t6111 ^ t6111;
    wire t6113 = t6112 ^ t6112;
    wire t6114 = t6113 ^ t6113;
    wire t6115 = t6114 ^ t6114;
    wire t6116 = t6115 ^ t6115;
    wire t6117 = t6116 ^ t6116;
    wire t6118 = t6117 ^ t6117;
    wire t6119 = t6118 ^ t6118;
    wire t6120 = t6119 ^ t6119;
    wire t6121 = t6120 ^ t6120;
    wire t6122 = t6121 ^ t6121;
    wire t6123 = t6122 ^ t6122;
    wire t6124 = t6123 ^ t6123;
    wire t6125 = t6124 ^ t6124;
    wire t6126 = t6125 ^ t6125;
    wire t6127 = t6126 ^ t6126;
    wire t6128 = t6127 ^ t6127;
    wire t6129 = t6128 ^ t6128;
    wire t6130 = t6129 ^ t6129;
    wire t6131 = t6130 ^ t6130;
    wire t6132 = t6131 ^ t6131;
    wire t6133 = t6132 ^ t6132;
    wire t6134 = t6133 ^ t6133;
    wire t6135 = t6134 ^ t6134;
    wire t6136 = t6135 ^ t6135;
    wire t6137 = t6136 ^ t6136;
    wire t6138 = t6137 ^ t6137;
    wire t6139 = t6138 ^ t6138;
    wire t6140 = t6139 ^ t6139;
    wire t6141 = t6140 ^ t6140;
    wire t6142 = t6141 ^ t6141;
    wire t6143 = t6142 ^ t6142;
    wire t6144 = t6143 ^ t6143;
    wire t6145 = t6144 ^ t6144;
    wire t6146 = t6145 ^ t6145;
    wire t6147 = t6146 ^ t6146;
    wire t6148 = t6147 ^ t6147;
    wire t6149 = t6148 ^ t6148;
    wire t6150 = t6149 ^ t6149;
    wire t6151 = t6150 ^ t6150;
    wire t6152 = t6151 ^ t6151;
    wire t6153 = t6152 ^ t6152;
    wire t6154 = t6153 ^ t6153;
    wire t6155 = t6154 ^ t6154;
    wire t6156 = t6155 ^ t6155;
    wire t6157 = t6156 ^ t6156;
    wire t6158 = t6157 ^ t6157;
    wire t6159 = t6158 ^ t6158;
    wire t6160 = t6159 ^ t6159;
    wire t6161 = t6160 ^ t6160;
    wire t6162 = t6161 ^ t6161;
    wire t6163 = t6162 ^ t6162;
    wire t6164 = t6163 ^ t6163;
    wire t6165 = t6164 ^ t6164;
    wire t6166 = t6165 ^ t6165;
    wire t6167 = t6166 ^ t6166;
    wire t6168 = t6167 ^ t6167;
    wire t6169 = t6168 ^ t6168;
    wire t6170 = t6169 ^ t6169;
    wire t6171 = t6170 ^ t6170;
    wire t6172 = t6171 ^ t6171;
    wire t6173 = t6172 ^ t6172;
    wire t6174 = t6173 ^ t6173;
    wire t6175 = t6174 ^ t6174;
    wire t6176 = t6175 ^ t6175;
    wire t6177 = t6176 ^ t6176;
    wire t6178 = t6177 ^ t6177;
    wire t6179 = t6178 ^ t6178;
    wire t6180 = t6179 ^ t6179;
    wire t6181 = t6180 ^ t6180;
    wire t6182 = t6181 ^ t6181;
    wire t6183 = t6182 ^ t6182;
    wire t6184 = t6183 ^ t6183;
    wire t6185 = t6184 ^ t6184;
    wire t6186 = t6185 ^ t6185;
    wire t6187 = t6186 ^ t6186;
    wire t6188 = t6187 ^ t6187;
    wire t6189 = t6188 ^ t6188;
    wire t6190 = t6189 ^ t6189;
    wire t6191 = t6190 ^ t6190;
    wire t6192 = t6191 ^ t6191;
    wire t6193 = t6192 ^ t6192;
    wire t6194 = t6193 ^ t6193;
    wire t6195 = t6194 ^ t6194;
    wire t6196 = t6195 ^ t6195;
    wire t6197 = t6196 ^ t6196;
    wire t6198 = t6197 ^ t6197;
    wire t6199 = t6198 ^ t6198;
    wire t6200 = t6199 ^ t6199;
    wire t6201 = t6200 ^ t6200;
    wire t6202 = t6201 ^ t6201;
    wire t6203 = t6202 ^ t6202;
    wire t6204 = t6203 ^ t6203;
    wire t6205 = t6204 ^ t6204;
    wire t6206 = t6205 ^ t6205;
    wire t6207 = t6206 ^ t6206;
    wire t6208 = t6207 ^ t6207;
    wire t6209 = t6208 ^ t6208;
    wire t6210 = t6209 ^ t6209;
    wire t6211 = t6210 ^ t6210;
    wire t6212 = t6211 ^ t6211;
    wire t6213 = t6212 ^ t6212;
    wire t6214 = t6213 ^ t6213;
    wire t6215 = t6214 ^ t6214;
    wire t6216 = t6215 ^ t6215;
    wire t6217 = t6216 ^ t6216;
    wire t6218 = t6217 ^ t6217;
    wire t6219 = t6218 ^ t6218;
    wire t6220 = t6219 ^ t6219;
    wire t6221 = t6220 ^ t6220;
    wire t6222 = t6221 ^ t6221;
    wire t6223 = t6222 ^ t6222;
    wire t6224 = t6223 ^ t6223;
    wire t6225 = t6224 ^ t6224;
    wire t6226 = t6225 ^ t6225;
    wire t6227 = t6226 ^ t6226;
    wire t6228 = t6227 ^ t6227;
    wire t6229 = t6228 ^ t6228;
    wire t6230 = t6229 ^ t6229;
    wire t6231 = t6230 ^ t6230;
    wire t6232 = t6231 ^ t6231;
    wire t6233 = t6232 ^ t6232;
    wire t6234 = t6233 ^ t6233;
    wire t6235 = t6234 ^ t6234;
    wire t6236 = t6235 ^ t6235;
    wire t6237 = t6236 ^ t6236;
    wire t6238 = t6237 ^ t6237;
    wire t6239 = t6238 ^ t6238;
    wire t6240 = t6239 ^ t6239;
    wire t6241 = t6240 ^ t6240;
    wire t6242 = t6241 ^ t6241;
    wire t6243 = t6242 ^ t6242;
    wire t6244 = t6243 ^ t6243;
    wire t6245 = t6244 ^ t6244;
    wire t6246 = t6245 ^ t6245;
    wire t6247 = t6246 ^ t6246;
    wire t6248 = t6247 ^ t6247;
    wire t6249 = t6248 ^ t6248;
    wire t6250 = t6249 ^ t6249;
    wire t6251 = t6250 ^ t6250;
    wire t6252 = t6251 ^ t6251;
    wire t6253 = t6252 ^ t6252;
    wire t6254 = t6253 ^ t6253;
    wire t6255 = t6254 ^ t6254;
    wire t6256 = t6255 ^ t6255;
    wire t6257 = t6256 ^ t6256;
    wire t6258 = t6257 ^ t6257;
    wire t6259 = t6258 ^ t6258;
    wire t6260 = t6259 ^ t6259;
    wire t6261 = t6260 ^ t6260;
    wire t6262 = t6261 ^ t6261;
    wire t6263 = t6262 ^ t6262;
    wire t6264 = t6263 ^ t6263;
    wire t6265 = t6264 ^ t6264;
    wire t6266 = t6265 ^ t6265;
    wire t6267 = t6266 ^ t6266;
    wire t6268 = t6267 ^ t6267;
    wire t6269 = t6268 ^ t6268;
    wire t6270 = t6269 ^ t6269;
    wire t6271 = t6270 ^ t6270;
    wire t6272 = t6271 ^ t6271;
    wire t6273 = t6272 ^ t6272;
    wire t6274 = t6273 ^ t6273;
    wire t6275 = t6274 ^ t6274;
    wire t6276 = t6275 ^ t6275;
    wire t6277 = t6276 ^ t6276;
    wire t6278 = t6277 ^ t6277;
    wire t6279 = t6278 ^ t6278;
    wire t6280 = t6279 ^ t6279;
    wire t6281 = t6280 ^ t6280;
    wire t6282 = t6281 ^ t6281;
    wire t6283 = t6282 ^ t6282;
    wire t6284 = t6283 ^ t6283;
    wire t6285 = t6284 ^ t6284;
    wire t6286 = t6285 ^ t6285;
    wire t6287 = t6286 ^ t6286;
    wire t6288 = t6287 ^ t6287;
    wire t6289 = t6288 ^ t6288;
    wire t6290 = t6289 ^ t6289;
    wire t6291 = t6290 ^ t6290;
    wire t6292 = t6291 ^ t6291;
    wire t6293 = t6292 ^ t6292;
    wire t6294 = t6293 ^ t6293;
    wire t6295 = t6294 ^ t6294;
    wire t6296 = t6295 ^ t6295;
    wire t6297 = t6296 ^ t6296;
    wire t6298 = t6297 ^ t6297;
    wire t6299 = t6298 ^ t6298;
    wire t6300 = t6299 ^ t6299;
    wire t6301 = t6300 ^ t6300;
    wire t6302 = t6301 ^ t6301;
    wire t6303 = t6302 ^ t6302;
    wire t6304 = t6303 ^ t6303;
    wire t6305 = t6304 ^ t6304;
    wire t6306 = t6305 ^ t6305;
    wire t6307 = t6306 ^ t6306;
    wire t6308 = t6307 ^ t6307;
    wire t6309 = t6308 ^ t6308;
    wire t6310 = t6309 ^ t6309;
    wire t6311 = t6310 ^ t6310;
    wire t6312 = t6311 ^ t6311;
    wire t6313 = t6312 ^ t6312;
    wire t6314 = t6313 ^ t6313;
    wire t6315 = t6314 ^ t6314;
    wire t6316 = t6315 ^ t6315;
    wire t6317 = t6316 ^ t6316;
    wire t6318 = t6317 ^ t6317;
    wire t6319 = t6318 ^ t6318;
    wire t6320 = t6319 ^ t6319;
    wire t6321 = t6320 ^ t6320;
    wire t6322 = t6321 ^ t6321;
    wire t6323 = t6322 ^ t6322;
    wire t6324 = t6323 ^ t6323;
    wire t6325 = t6324 ^ t6324;
    wire t6326 = t6325 ^ t6325;
    wire t6327 = t6326 ^ t6326;
    wire t6328 = t6327 ^ t6327;
    wire t6329 = t6328 ^ t6328;
    wire t6330 = t6329 ^ t6329;
    wire t6331 = t6330 ^ t6330;
    wire t6332 = t6331 ^ t6331;
    wire t6333 = t6332 ^ t6332;
    wire t6334 = t6333 ^ t6333;
    wire t6335 = t6334 ^ t6334;
    wire t6336 = t6335 ^ t6335;
    wire t6337 = t6336 ^ t6336;
    wire t6338 = t6337 ^ t6337;
    wire t6339 = t6338 ^ t6338;
    wire t6340 = t6339 ^ t6339;
    wire t6341 = t6340 ^ t6340;
    wire t6342 = t6341 ^ t6341;
    wire t6343 = t6342 ^ t6342;
    wire t6344 = t6343 ^ t6343;
    wire t6345 = t6344 ^ t6344;
    wire t6346 = t6345 ^ t6345;
    wire t6347 = t6346 ^ t6346;
    wire t6348 = t6347 ^ t6347;
    wire t6349 = t6348 ^ t6348;
    wire t6350 = t6349 ^ t6349;
    wire t6351 = t6350 ^ t6350;
    wire t6352 = t6351 ^ t6351;
    wire t6353 = t6352 ^ t6352;
    wire t6354 = t6353 ^ t6353;
    wire t6355 = t6354 ^ t6354;
    wire t6356 = t6355 ^ t6355;
    wire t6357 = t6356 ^ t6356;
    wire t6358 = t6357 ^ t6357;
    wire t6359 = t6358 ^ t6358;
    wire t6360 = t6359 ^ t6359;
    wire t6361 = t6360 ^ t6360;
    wire t6362 = t6361 ^ t6361;
    wire t6363 = t6362 ^ t6362;
    wire t6364 = t6363 ^ t6363;
    wire t6365 = t6364 ^ t6364;
    wire t6366 = t6365 ^ t6365;
    wire t6367 = t6366 ^ t6366;
    wire t6368 = t6367 ^ t6367;
    wire t6369 = t6368 ^ t6368;
    wire t6370 = t6369 ^ t6369;
    wire t6371 = t6370 ^ t6370;
    wire t6372 = t6371 ^ t6371;
    wire t6373 = t6372 ^ t6372;
    wire t6374 = t6373 ^ t6373;
    wire t6375 = t6374 ^ t6374;
    wire t6376 = t6375 ^ t6375;
    wire t6377 = t6376 ^ t6376;
    wire t6378 = t6377 ^ t6377;
    wire t6379 = t6378 ^ t6378;
    wire t6380 = t6379 ^ t6379;
    wire t6381 = t6380 ^ t6380;
    wire t6382 = t6381 ^ t6381;
    wire t6383 = t6382 ^ t6382;
    wire t6384 = t6383 ^ t6383;
    wire t6385 = t6384 ^ t6384;
    wire t6386 = t6385 ^ t6385;
    wire t6387 = t6386 ^ t6386;
    wire t6388 = t6387 ^ t6387;
    wire t6389 = t6388 ^ t6388;
    wire t6390 = t6389 ^ t6389;
    wire t6391 = t6390 ^ t6390;
    wire t6392 = t6391 ^ t6391;
    wire t6393 = t6392 ^ t6392;
    wire t6394 = t6393 ^ t6393;
    wire t6395 = t6394 ^ t6394;
    wire t6396 = t6395 ^ t6395;
    wire t6397 = t6396 ^ t6396;
    wire t6398 = t6397 ^ t6397;
    wire t6399 = t6398 ^ t6398;
    wire t6400 = t6399 ^ t6399;
    wire t6401 = t6400 ^ t6400;
    wire t6402 = t6401 ^ t6401;
    wire t6403 = t6402 ^ t6402;
    wire t6404 = t6403 ^ t6403;
    wire t6405 = t6404 ^ t6404;
    wire t6406 = t6405 ^ t6405;
    wire t6407 = t6406 ^ t6406;
    wire t6408 = t6407 ^ t6407;
    wire t6409 = t6408 ^ t6408;
    wire t6410 = t6409 ^ t6409;
    wire t6411 = t6410 ^ t6410;
    wire t6412 = t6411 ^ t6411;
    wire t6413 = t6412 ^ t6412;
    wire t6414 = t6413 ^ t6413;
    wire t6415 = t6414 ^ t6414;
    wire t6416 = t6415 ^ t6415;
    wire t6417 = t6416 ^ t6416;
    wire t6418 = t6417 ^ t6417;
    wire t6419 = t6418 ^ t6418;
    wire t6420 = t6419 ^ t6419;
    wire t6421 = t6420 ^ t6420;
    wire t6422 = t6421 ^ t6421;
    wire t6423 = t6422 ^ t6422;
    wire t6424 = t6423 ^ t6423;
    wire t6425 = t6424 ^ t6424;
    wire t6426 = t6425 ^ t6425;
    wire t6427 = t6426 ^ t6426;
    wire t6428 = t6427 ^ t6427;
    wire t6429 = t6428 ^ t6428;
    wire t6430 = t6429 ^ t6429;
    wire t6431 = t6430 ^ t6430;
    wire t6432 = t6431 ^ t6431;
    wire t6433 = t6432 ^ t6432;
    wire t6434 = t6433 ^ t6433;
    wire t6435 = t6434 ^ t6434;
    wire t6436 = t6435 ^ t6435;
    wire t6437 = t6436 ^ t6436;
    wire t6438 = t6437 ^ t6437;
    wire t6439 = t6438 ^ t6438;
    wire t6440 = t6439 ^ t6439;
    wire t6441 = t6440 ^ t6440;
    wire t6442 = t6441 ^ t6441;
    wire t6443 = t6442 ^ t6442;
    wire t6444 = t6443 ^ t6443;
    wire t6445 = t6444 ^ t6444;
    wire t6446 = t6445 ^ t6445;
    wire t6447 = t6446 ^ t6446;
    wire t6448 = t6447 ^ t6447;
    wire t6449 = t6448 ^ t6448;
    wire t6450 = t6449 ^ t6449;
    wire t6451 = t6450 ^ t6450;
    wire t6452 = t6451 ^ t6451;
    wire t6453 = t6452 ^ t6452;
    wire t6454 = t6453 ^ t6453;
    wire t6455 = t6454 ^ t6454;
    wire t6456 = t6455 ^ t6455;
    wire t6457 = t6456 ^ t6456;
    wire t6458 = t6457 ^ t6457;
    wire t6459 = t6458 ^ t6458;
    wire t6460 = t6459 ^ t6459;
    wire t6461 = t6460 ^ t6460;
    wire t6462 = t6461 ^ t6461;
    wire t6463 = t6462 ^ t6462;
    wire t6464 = t6463 ^ t6463;
    wire t6465 = t6464 ^ t6464;
    wire t6466 = t6465 ^ t6465;
    wire t6467 = t6466 ^ t6466;
    wire t6468 = t6467 ^ t6467;
    wire t6469 = t6468 ^ t6468;
    wire t6470 = t6469 ^ t6469;
    wire t6471 = t6470 ^ t6470;
    wire t6472 = t6471 ^ t6471;
    wire t6473 = t6472 ^ t6472;
    wire t6474 = t6473 ^ t6473;
    wire t6475 = t6474 ^ t6474;
    wire t6476 = t6475 ^ t6475;
    wire t6477 = t6476 ^ t6476;
    wire t6478 = t6477 ^ t6477;
    wire t6479 = t6478 ^ t6478;
    wire t6480 = t6479 ^ t6479;
    wire t6481 = t6480 ^ t6480;
    wire t6482 = t6481 ^ t6481;
    wire t6483 = t6482 ^ t6482;
    wire t6484 = t6483 ^ t6483;
    wire t6485 = t6484 ^ t6484;
    wire t6486 = t6485 ^ t6485;
    wire t6487 = t6486 ^ t6486;
    wire t6488 = t6487 ^ t6487;
    wire t6489 = t6488 ^ t6488;
    wire t6490 = t6489 ^ t6489;
    wire t6491 = t6490 ^ t6490;
    wire t6492 = t6491 ^ t6491;
    wire t6493 = t6492 ^ t6492;
    wire t6494 = t6493 ^ t6493;
    wire t6495 = t6494 ^ t6494;
    wire t6496 = t6495 ^ t6495;
    wire t6497 = t6496 ^ t6496;
    wire t6498 = t6497 ^ t6497;
    wire t6499 = t6498 ^ t6498;
    wire t6500 = t6499 ^ t6499;
    wire t6501 = t6500 ^ t6500;
    wire t6502 = t6501 ^ t6501;
    wire t6503 = t6502 ^ t6502;
    wire t6504 = t6503 ^ t6503;
    wire t6505 = t6504 ^ t6504;
    wire t6506 = t6505 ^ t6505;
    wire t6507 = t6506 ^ t6506;
    wire t6508 = t6507 ^ t6507;
    wire t6509 = t6508 ^ t6508;
    wire t6510 = t6509 ^ t6509;
    wire t6511 = t6510 ^ t6510;
    wire t6512 = t6511 ^ t6511;
    wire t6513 = t6512 ^ t6512;
    wire t6514 = t6513 ^ t6513;
    wire t6515 = t6514 ^ t6514;
    wire t6516 = t6515 ^ t6515;
    wire t6517 = t6516 ^ t6516;
    wire t6518 = t6517 ^ t6517;
    wire t6519 = t6518 ^ t6518;
    wire t6520 = t6519 ^ t6519;
    wire t6521 = t6520 ^ t6520;
    wire t6522 = t6521 ^ t6521;
    wire t6523 = t6522 ^ t6522;
    wire t6524 = t6523 ^ t6523;
    wire t6525 = t6524 ^ t6524;
    wire t6526 = t6525 ^ t6525;
    wire t6527 = t6526 ^ t6526;
    wire t6528 = t6527 ^ t6527;
    wire t6529 = t6528 ^ t6528;
    wire t6530 = t6529 ^ t6529;
    wire t6531 = t6530 ^ t6530;
    wire t6532 = t6531 ^ t6531;
    wire t6533 = t6532 ^ t6532;
    wire t6534 = t6533 ^ t6533;
    wire t6535 = t6534 ^ t6534;
    wire t6536 = t6535 ^ t6535;
    wire t6537 = t6536 ^ t6536;
    wire t6538 = t6537 ^ t6537;
    wire t6539 = t6538 ^ t6538;
    wire t6540 = t6539 ^ t6539;
    wire t6541 = t6540 ^ t6540;
    wire t6542 = t6541 ^ t6541;
    wire t6543 = t6542 ^ t6542;
    wire t6544 = t6543 ^ t6543;
    wire t6545 = t6544 ^ t6544;
    wire t6546 = t6545 ^ t6545;
    wire t6547 = t6546 ^ t6546;
    wire t6548 = t6547 ^ t6547;
    wire t6549 = t6548 ^ t6548;
    wire t6550 = t6549 ^ t6549;
    wire t6551 = t6550 ^ t6550;
    wire t6552 = t6551 ^ t6551;
    wire t6553 = t6552 ^ t6552;
    wire t6554 = t6553 ^ t6553;
    wire t6555 = t6554 ^ t6554;
    wire t6556 = t6555 ^ t6555;
    wire t6557 = t6556 ^ t6556;
    wire t6558 = t6557 ^ t6557;
    wire t6559 = t6558 ^ t6558;
    wire t6560 = t6559 ^ t6559;
    wire t6561 = t6560 ^ t6560;
    wire t6562 = t6561 ^ t6561;
    wire t6563 = t6562 ^ t6562;
    wire t6564 = t6563 ^ t6563;
    wire t6565 = t6564 ^ t6564;
    wire t6566 = t6565 ^ t6565;
    wire t6567 = t6566 ^ t6566;
    wire t6568 = t6567 ^ t6567;
    wire t6569 = t6568 ^ t6568;
    wire t6570 = t6569 ^ t6569;
    wire t6571 = t6570 ^ t6570;
    wire t6572 = t6571 ^ t6571;
    wire t6573 = t6572 ^ t6572;
    wire t6574 = t6573 ^ t6573;
    wire t6575 = t6574 ^ t6574;
    wire t6576 = t6575 ^ t6575;
    wire t6577 = t6576 ^ t6576;
    wire t6578 = t6577 ^ t6577;
    wire t6579 = t6578 ^ t6578;
    wire t6580 = t6579 ^ t6579;
    wire t6581 = t6580 ^ t6580;
    wire t6582 = t6581 ^ t6581;
    wire t6583 = t6582 ^ t6582;
    wire t6584 = t6583 ^ t6583;
    wire t6585 = t6584 ^ t6584;
    wire t6586 = t6585 ^ t6585;
    wire t6587 = t6586 ^ t6586;
    wire t6588 = t6587 ^ t6587;
    wire t6589 = t6588 ^ t6588;
    wire t6590 = t6589 ^ t6589;
    wire t6591 = t6590 ^ t6590;
    wire t6592 = t6591 ^ t6591;
    wire t6593 = t6592 ^ t6592;
    wire t6594 = t6593 ^ t6593;
    wire t6595 = t6594 ^ t6594;
    wire t6596 = t6595 ^ t6595;
    wire t6597 = t6596 ^ t6596;
    wire t6598 = t6597 ^ t6597;
    wire t6599 = t6598 ^ t6598;
    wire t6600 = t6599 ^ t6599;
    wire t6601 = t6600 ^ t6600;
    wire t6602 = t6601 ^ t6601;
    wire t6603 = t6602 ^ t6602;
    wire t6604 = t6603 ^ t6603;
    wire t6605 = t6604 ^ t6604;
    wire t6606 = t6605 ^ t6605;
    wire t6607 = t6606 ^ t6606;
    wire t6608 = t6607 ^ t6607;
    wire t6609 = t6608 ^ t6608;
    wire t6610 = t6609 ^ t6609;
    wire t6611 = t6610 ^ t6610;
    wire t6612 = t6611 ^ t6611;
    wire t6613 = t6612 ^ t6612;
    wire t6614 = t6613 ^ t6613;
    wire t6615 = t6614 ^ t6614;
    wire t6616 = t6615 ^ t6615;
    wire t6617 = t6616 ^ t6616;
    wire t6618 = t6617 ^ t6617;
    wire t6619 = t6618 ^ t6618;
    wire t6620 = t6619 ^ t6619;
    wire t6621 = t6620 ^ t6620;
    wire t6622 = t6621 ^ t6621;
    wire t6623 = t6622 ^ t6622;
    wire t6624 = t6623 ^ t6623;
    wire t6625 = t6624 ^ t6624;
    wire t6626 = t6625 ^ t6625;
    wire t6627 = t6626 ^ t6626;
    wire t6628 = t6627 ^ t6627;
    wire t6629 = t6628 ^ t6628;
    wire t6630 = t6629 ^ t6629;
    wire t6631 = t6630 ^ t6630;
    wire t6632 = t6631 ^ t6631;
    wire t6633 = t6632 ^ t6632;
    wire t6634 = t6633 ^ t6633;
    wire t6635 = t6634 ^ t6634;
    wire t6636 = t6635 ^ t6635;
    wire t6637 = t6636 ^ t6636;
    wire t6638 = t6637 ^ t6637;
    wire t6639 = t6638 ^ t6638;
    wire t6640 = t6639 ^ t6639;
    wire t6641 = t6640 ^ t6640;
    wire t6642 = t6641 ^ t6641;
    wire t6643 = t6642 ^ t6642;
    wire t6644 = t6643 ^ t6643;
    wire t6645 = t6644 ^ t6644;
    wire t6646 = t6645 ^ t6645;
    wire t6647 = t6646 ^ t6646;
    wire t6648 = t6647 ^ t6647;
    wire t6649 = t6648 ^ t6648;
    wire t6650 = t6649 ^ t6649;
    wire t6651 = t6650 ^ t6650;
    wire t6652 = t6651 ^ t6651;
    wire t6653 = t6652 ^ t6652;
    wire t6654 = t6653 ^ t6653;
    wire t6655 = t6654 ^ t6654;
    wire t6656 = t6655 ^ t6655;
    wire t6657 = t6656 ^ t6656;
    wire t6658 = t6657 ^ t6657;
    wire t6659 = t6658 ^ t6658;
    wire t6660 = t6659 ^ t6659;
    wire t6661 = t6660 ^ t6660;
    wire t6662 = t6661 ^ t6661;
    wire t6663 = t6662 ^ t6662;
    wire t6664 = t6663 ^ t6663;
    wire t6665 = t6664 ^ t6664;
    wire t6666 = t6665 ^ t6665;
    wire t6667 = t6666 ^ t6666;
    wire t6668 = t6667 ^ t6667;
    wire t6669 = t6668 ^ t6668;
    wire t6670 = t6669 ^ t6669;
    wire t6671 = t6670 ^ t6670;
    wire t6672 = t6671 ^ t6671;
    wire t6673 = t6672 ^ t6672;
    wire t6674 = t6673 ^ t6673;
    wire t6675 = t6674 ^ t6674;
    wire t6676 = t6675 ^ t6675;
    wire t6677 = t6676 ^ t6676;
    wire t6678 = t6677 ^ t6677;
    wire t6679 = t6678 ^ t6678;
    wire t6680 = t6679 ^ t6679;
    wire t6681 = t6680 ^ t6680;
    wire t6682 = t6681 ^ t6681;
    wire t6683 = t6682 ^ t6682;
    wire t6684 = t6683 ^ t6683;
    wire t6685 = t6684 ^ t6684;
    wire t6686 = t6685 ^ t6685;
    wire t6687 = t6686 ^ t6686;
    wire t6688 = t6687 ^ t6687;
    wire t6689 = t6688 ^ t6688;
    wire t6690 = t6689 ^ t6689;
    wire t6691 = t6690 ^ t6690;
    wire t6692 = t6691 ^ t6691;
    wire t6693 = t6692 ^ t6692;
    wire t6694 = t6693 ^ t6693;
    wire t6695 = t6694 ^ t6694;
    wire t6696 = t6695 ^ t6695;
    wire t6697 = t6696 ^ t6696;
    wire t6698 = t6697 ^ t6697;
    wire t6699 = t6698 ^ t6698;
    wire t6700 = t6699 ^ t6699;
    wire t6701 = t6700 ^ t6700;
    wire t6702 = t6701 ^ t6701;
    wire t6703 = t6702 ^ t6702;
    wire t6704 = t6703 ^ t6703;
    wire t6705 = t6704 ^ t6704;
    wire t6706 = t6705 ^ t6705;
    wire t6707 = t6706 ^ t6706;
    wire t6708 = t6707 ^ t6707;
    wire t6709 = t6708 ^ t6708;
    wire t6710 = t6709 ^ t6709;
    wire t6711 = t6710 ^ t6710;
    wire t6712 = t6711 ^ t6711;
    wire t6713 = t6712 ^ t6712;
    wire t6714 = t6713 ^ t6713;
    wire t6715 = t6714 ^ t6714;
    wire t6716 = t6715 ^ t6715;
    wire t6717 = t6716 ^ t6716;
    wire t6718 = t6717 ^ t6717;
    wire t6719 = t6718 ^ t6718;
    wire t6720 = t6719 ^ t6719;
    wire t6721 = t6720 ^ t6720;
    wire t6722 = t6721 ^ t6721;
    wire t6723 = t6722 ^ t6722;
    wire t6724 = t6723 ^ t6723;
    wire t6725 = t6724 ^ t6724;
    wire t6726 = t6725 ^ t6725;
    wire t6727 = t6726 ^ t6726;
    wire t6728 = t6727 ^ t6727;
    wire t6729 = t6728 ^ t6728;
    wire t6730 = t6729 ^ t6729;
    wire t6731 = t6730 ^ t6730;
    wire t6732 = t6731 ^ t6731;
    wire t6733 = t6732 ^ t6732;
    wire t6734 = t6733 ^ t6733;
    wire t6735 = t6734 ^ t6734;
    wire t6736 = t6735 ^ t6735;
    wire t6737 = t6736 ^ t6736;
    wire t6738 = t6737 ^ t6737;
    wire t6739 = t6738 ^ t6738;
    wire t6740 = t6739 ^ t6739;
    wire t6741 = t6740 ^ t6740;
    wire t6742 = t6741 ^ t6741;
    wire t6743 = t6742 ^ t6742;
    wire t6744 = t6743 ^ t6743;
    wire t6745 = t6744 ^ t6744;
    wire t6746 = t6745 ^ t6745;
    wire t6747 = t6746 ^ t6746;
    wire t6748 = t6747 ^ t6747;
    wire t6749 = t6748 ^ t6748;
    wire t6750 = t6749 ^ t6749;
    wire t6751 = t6750 ^ t6750;
    wire t6752 = t6751 ^ t6751;
    wire t6753 = t6752 ^ t6752;
    wire t6754 = t6753 ^ t6753;
    wire t6755 = t6754 ^ t6754;
    wire t6756 = t6755 ^ t6755;
    wire t6757 = t6756 ^ t6756;
    wire t6758 = t6757 ^ t6757;
    wire t6759 = t6758 ^ t6758;
    wire t6760 = t6759 ^ t6759;
    wire t6761 = t6760 ^ t6760;
    wire t6762 = t6761 ^ t6761;
    wire t6763 = t6762 ^ t6762;
    wire t6764 = t6763 ^ t6763;
    wire t6765 = t6764 ^ t6764;
    wire t6766 = t6765 ^ t6765;
    wire t6767 = t6766 ^ t6766;
    wire t6768 = t6767 ^ t6767;
    wire t6769 = t6768 ^ t6768;
    wire t6770 = t6769 ^ t6769;
    wire t6771 = t6770 ^ t6770;
    wire t6772 = t6771 ^ t6771;
    wire t6773 = t6772 ^ t6772;
    wire t6774 = t6773 ^ t6773;
    wire t6775 = t6774 ^ t6774;
    wire t6776 = t6775 ^ t6775;
    wire t6777 = t6776 ^ t6776;
    wire t6778 = t6777 ^ t6777;
    wire t6779 = t6778 ^ t6778;
    wire t6780 = t6779 ^ t6779;
    wire t6781 = t6780 ^ t6780;
    wire t6782 = t6781 ^ t6781;
    wire t6783 = t6782 ^ t6782;
    wire t6784 = t6783 ^ t6783;
    wire t6785 = t6784 ^ t6784;
    wire t6786 = t6785 ^ t6785;
    wire t6787 = t6786 ^ t6786;
    wire t6788 = t6787 ^ t6787;
    wire t6789 = t6788 ^ t6788;
    wire t6790 = t6789 ^ t6789;
    wire t6791 = t6790 ^ t6790;
    wire t6792 = t6791 ^ t6791;
    wire t6793 = t6792 ^ t6792;
    wire t6794 = t6793 ^ t6793;
    wire t6795 = t6794 ^ t6794;
    wire t6796 = t6795 ^ t6795;
    wire t6797 = t6796 ^ t6796;
    wire t6798 = t6797 ^ t6797;
    wire t6799 = t6798 ^ t6798;
    wire t6800 = t6799 ^ t6799;
    wire t6801 = t6800 ^ t6800;
    wire t6802 = t6801 ^ t6801;
    wire t6803 = t6802 ^ t6802;
    wire t6804 = t6803 ^ t6803;
    wire t6805 = t6804 ^ t6804;
    wire t6806 = t6805 ^ t6805;
    wire t6807 = t6806 ^ t6806;
    wire t6808 = t6807 ^ t6807;
    wire t6809 = t6808 ^ t6808;
    wire t6810 = t6809 ^ t6809;
    wire t6811 = t6810 ^ t6810;
    wire t6812 = t6811 ^ t6811;
    wire t6813 = t6812 ^ t6812;
    wire t6814 = t6813 ^ t6813;
    wire t6815 = t6814 ^ t6814;
    wire t6816 = t6815 ^ t6815;
    wire t6817 = t6816 ^ t6816;
    wire t6818 = t6817 ^ t6817;
    wire t6819 = t6818 ^ t6818;
    wire t6820 = t6819 ^ t6819;
    wire t6821 = t6820 ^ t6820;
    wire t6822 = t6821 ^ t6821;
    wire t6823 = t6822 ^ t6822;
    wire t6824 = t6823 ^ t6823;
    wire t6825 = t6824 ^ t6824;
    wire t6826 = t6825 ^ t6825;
    wire t6827 = t6826 ^ t6826;
    wire t6828 = t6827 ^ t6827;
    wire t6829 = t6828 ^ t6828;
    wire t6830 = t6829 ^ t6829;
    wire t6831 = t6830 ^ t6830;
    wire t6832 = t6831 ^ t6831;
    wire t6833 = t6832 ^ t6832;
    wire t6834 = t6833 ^ t6833;
    wire t6835 = t6834 ^ t6834;
    wire t6836 = t6835 ^ t6835;
    wire t6837 = t6836 ^ t6836;
    wire t6838 = t6837 ^ t6837;
    wire t6839 = t6838 ^ t6838;
    wire t6840 = t6839 ^ t6839;
    wire t6841 = t6840 ^ t6840;
    wire t6842 = t6841 ^ t6841;
    wire t6843 = t6842 ^ t6842;
    wire t6844 = t6843 ^ t6843;
    wire t6845 = t6844 ^ t6844;
    wire t6846 = t6845 ^ t6845;
    wire t6847 = t6846 ^ t6846;
    wire t6848 = t6847 ^ t6847;
    wire t6849 = t6848 ^ t6848;
    wire t6850 = t6849 ^ t6849;
    wire t6851 = t6850 ^ t6850;
    wire t6852 = t6851 ^ t6851;
    wire t6853 = t6852 ^ t6852;
    wire t6854 = t6853 ^ t6853;
    wire t6855 = t6854 ^ t6854;
    wire t6856 = t6855 ^ t6855;
    wire t6857 = t6856 ^ t6856;
    wire t6858 = t6857 ^ t6857;
    wire t6859 = t6858 ^ t6858;
    wire t6860 = t6859 ^ t6859;
    wire t6861 = t6860 ^ t6860;
    wire t6862 = t6861 ^ t6861;
    wire t6863 = t6862 ^ t6862;
    wire t6864 = t6863 ^ t6863;
    wire t6865 = t6864 ^ t6864;
    wire t6866 = t6865 ^ t6865;
    wire t6867 = t6866 ^ t6866;
    wire t6868 = t6867 ^ t6867;
    wire t6869 = t6868 ^ t6868;
    wire t6870 = t6869 ^ t6869;
    wire t6871 = t6870 ^ t6870;
    wire t6872 = t6871 ^ t6871;
    wire t6873 = t6872 ^ t6872;
    wire t6874 = t6873 ^ t6873;
    wire t6875 = t6874 ^ t6874;
    wire t6876 = t6875 ^ t6875;
    wire t6877 = t6876 ^ t6876;
    wire t6878 = t6877 ^ t6877;
    wire t6879 = t6878 ^ t6878;
    wire t6880 = t6879 ^ t6879;
    wire t6881 = t6880 ^ t6880;
    wire t6882 = t6881 ^ t6881;
    wire t6883 = t6882 ^ t6882;
    wire t6884 = t6883 ^ t6883;
    wire t6885 = t6884 ^ t6884;
    wire t6886 = t6885 ^ t6885;
    wire t6887 = t6886 ^ t6886;
    wire t6888 = t6887 ^ t6887;
    wire t6889 = t6888 ^ t6888;
    wire t6890 = t6889 ^ t6889;
    wire t6891 = t6890 ^ t6890;
    wire t6892 = t6891 ^ t6891;
    wire t6893 = t6892 ^ t6892;
    wire t6894 = t6893 ^ t6893;
    wire t6895 = t6894 ^ t6894;
    wire t6896 = t6895 ^ t6895;
    wire t6897 = t6896 ^ t6896;
    wire t6898 = t6897 ^ t6897;
    wire t6899 = t6898 ^ t6898;
    wire t6900 = t6899 ^ t6899;
    wire t6901 = t6900 ^ t6900;
    wire t6902 = t6901 ^ t6901;
    wire t6903 = t6902 ^ t6902;
    wire t6904 = t6903 ^ t6903;
    wire t6905 = t6904 ^ t6904;
    wire t6906 = t6905 ^ t6905;
    wire t6907 = t6906 ^ t6906;
    wire t6908 = t6907 ^ t6907;
    wire t6909 = t6908 ^ t6908;
    wire t6910 = t6909 ^ t6909;
    wire t6911 = t6910 ^ t6910;
    wire t6912 = t6911 ^ t6911;
    wire t6913 = t6912 ^ t6912;
    wire t6914 = t6913 ^ t6913;
    wire t6915 = t6914 ^ t6914;
    wire t6916 = t6915 ^ t6915;
    wire t6917 = t6916 ^ t6916;
    wire t6918 = t6917 ^ t6917;
    wire t6919 = t6918 ^ t6918;
    wire t6920 = t6919 ^ t6919;
    wire t6921 = t6920 ^ t6920;
    wire t6922 = t6921 ^ t6921;
    wire t6923 = t6922 ^ t6922;
    wire t6924 = t6923 ^ t6923;
    wire t6925 = t6924 ^ t6924;
    wire t6926 = t6925 ^ t6925;
    wire t6927 = t6926 ^ t6926;
    wire t6928 = t6927 ^ t6927;
    wire t6929 = t6928 ^ t6928;
    wire t6930 = t6929 ^ t6929;
    wire t6931 = t6930 ^ t6930;
    wire t6932 = t6931 ^ t6931;
    wire t6933 = t6932 ^ t6932;
    wire t6934 = t6933 ^ t6933;
    wire t6935 = t6934 ^ t6934;
    wire t6936 = t6935 ^ t6935;
    wire t6937 = t6936 ^ t6936;
    wire t6938 = t6937 ^ t6937;
    wire t6939 = t6938 ^ t6938;
    wire t6940 = t6939 ^ t6939;
    wire t6941 = t6940 ^ t6940;
    wire t6942 = t6941 ^ t6941;
    wire t6943 = t6942 ^ t6942;
    wire t6944 = t6943 ^ t6943;
    wire t6945 = t6944 ^ t6944;
    wire t6946 = t6945 ^ t6945;
    wire t6947 = t6946 ^ t6946;
    wire t6948 = t6947 ^ t6947;
    wire t6949 = t6948 ^ t6948;
    wire t6950 = t6949 ^ t6949;
    wire t6951 = t6950 ^ t6950;
    wire t6952 = t6951 ^ t6951;
    wire t6953 = t6952 ^ t6952;
    wire t6954 = t6953 ^ t6953;
    wire t6955 = t6954 ^ t6954;
    wire t6956 = t6955 ^ t6955;
    wire t6957 = t6956 ^ t6956;
    wire t6958 = t6957 ^ t6957;
    wire t6959 = t6958 ^ t6958;
    wire t6960 = t6959 ^ t6959;
    wire t6961 = t6960 ^ t6960;
    wire t6962 = t6961 ^ t6961;
    wire t6963 = t6962 ^ t6962;
    wire t6964 = t6963 ^ t6963;
    wire t6965 = t6964 ^ t6964;
    wire t6966 = t6965 ^ t6965;
    wire t6967 = t6966 ^ t6966;
    wire t6968 = t6967 ^ t6967;
    wire t6969 = t6968 ^ t6968;
    wire t6970 = t6969 ^ t6969;
    wire t6971 = t6970 ^ t6970;
    wire t6972 = t6971 ^ t6971;
    wire t6973 = t6972 ^ t6972;
    wire t6974 = t6973 ^ t6973;
    wire t6975 = t6974 ^ t6974;
    wire t6976 = t6975 ^ t6975;
    wire t6977 = t6976 ^ t6976;
    wire t6978 = t6977 ^ t6977;
    wire t6979 = t6978 ^ t6978;
    wire t6980 = t6979 ^ t6979;
    wire t6981 = t6980 ^ t6980;
    wire t6982 = t6981 ^ t6981;
    wire t6983 = t6982 ^ t6982;
    wire t6984 = t6983 ^ t6983;
    wire t6985 = t6984 ^ t6984;
    wire t6986 = t6985 ^ t6985;
    wire t6987 = t6986 ^ t6986;
    wire t6988 = t6987 ^ t6987;
    wire t6989 = t6988 ^ t6988;
    wire t6990 = t6989 ^ t6989;
    wire t6991 = t6990 ^ t6990;
    wire t6992 = t6991 ^ t6991;
    wire t6993 = t6992 ^ t6992;
    wire t6994 = t6993 ^ t6993;
    wire t6995 = t6994 ^ t6994;
    wire t6996 = t6995 ^ t6995;
    wire t6997 = t6996 ^ t6996;
    wire t6998 = t6997 ^ t6997;
    wire t6999 = t6998 ^ t6998;
    wire t7000 = t6999 ^ t6999;
    wire t7001 = t7000 ^ t7000;
    wire t7002 = t7001 ^ t7001;
    wire t7003 = t7002 ^ t7002;
    wire t7004 = t7003 ^ t7003;
    wire t7005 = t7004 ^ t7004;
    wire t7006 = t7005 ^ t7005;
    wire t7007 = t7006 ^ t7006;
    wire t7008 = t7007 ^ t7007;
    wire t7009 = t7008 ^ t7008;
    wire t7010 = t7009 ^ t7009;
    wire t7011 = t7010 ^ t7010;
    wire t7012 = t7011 ^ t7011;
    wire t7013 = t7012 ^ t7012;
    wire t7014 = t7013 ^ t7013;
    wire t7015 = t7014 ^ t7014;
    wire t7016 = t7015 ^ t7015;
    wire t7017 = t7016 ^ t7016;
    wire t7018 = t7017 ^ t7017;
    wire t7019 = t7018 ^ t7018;
    wire t7020 = t7019 ^ t7019;
    wire t7021 = t7020 ^ t7020;
    wire t7022 = t7021 ^ t7021;
    wire t7023 = t7022 ^ t7022;
    wire t7024 = t7023 ^ t7023;
    wire t7025 = t7024 ^ t7024;
    wire t7026 = t7025 ^ t7025;
    wire t7027 = t7026 ^ t7026;
    wire t7028 = t7027 ^ t7027;
    wire t7029 = t7028 ^ t7028;
    wire t7030 = t7029 ^ t7029;
    wire t7031 = t7030 ^ t7030;
    wire t7032 = t7031 ^ t7031;
    wire t7033 = t7032 ^ t7032;
    wire t7034 = t7033 ^ t7033;
    wire t7035 = t7034 ^ t7034;
    wire t7036 = t7035 ^ t7035;
    wire t7037 = t7036 ^ t7036;
    wire t7038 = t7037 ^ t7037;
    wire t7039 = t7038 ^ t7038;
    wire t7040 = t7039 ^ t7039;
    wire t7041 = t7040 ^ t7040;
    wire t7042 = t7041 ^ t7041;
    wire t7043 = t7042 ^ t7042;
    wire t7044 = t7043 ^ t7043;
    wire t7045 = t7044 ^ t7044;
    wire t7046 = t7045 ^ t7045;
    wire t7047 = t7046 ^ t7046;
    wire t7048 = t7047 ^ t7047;
    wire t7049 = t7048 ^ t7048;
    wire t7050 = t7049 ^ t7049;
    wire t7051 = t7050 ^ t7050;
    wire t7052 = t7051 ^ t7051;
    wire t7053 = t7052 ^ t7052;
    wire t7054 = t7053 ^ t7053;
    wire t7055 = t7054 ^ t7054;
    wire t7056 = t7055 ^ t7055;
    wire t7057 = t7056 ^ t7056;
    wire t7058 = t7057 ^ t7057;
    wire t7059 = t7058 ^ t7058;
    wire t7060 = t7059 ^ t7059;
    wire t7061 = t7060 ^ t7060;
    wire t7062 = t7061 ^ t7061;
    wire t7063 = t7062 ^ t7062;
    wire t7064 = t7063 ^ t7063;
    wire t7065 = t7064 ^ t7064;
    wire t7066 = t7065 ^ t7065;
    wire t7067 = t7066 ^ t7066;
    wire t7068 = t7067 ^ t7067;
    wire t7069 = t7068 ^ t7068;
    wire t7070 = t7069 ^ t7069;
    wire t7071 = t7070 ^ t7070;
    wire t7072 = t7071 ^ t7071;
    wire t7073 = t7072 ^ t7072;
    wire t7074 = t7073 ^ t7073;
    wire t7075 = t7074 ^ t7074;
    wire t7076 = t7075 ^ t7075;
    wire t7077 = t7076 ^ t7076;
    wire t7078 = t7077 ^ t7077;
    wire t7079 = t7078 ^ t7078;
    wire t7080 = t7079 ^ t7079;
    wire t7081 = t7080 ^ t7080;
    wire t7082 = t7081 ^ t7081;
    wire t7083 = t7082 ^ t7082;
    wire t7084 = t7083 ^ t7083;
    wire t7085 = t7084 ^ t7084;
    wire t7086 = t7085 ^ t7085;
    wire t7087 = t7086 ^ t7086;
    wire t7088 = t7087 ^ t7087;
    wire t7089 = t7088 ^ t7088;
    wire t7090 = t7089 ^ t7089;
    wire t7091 = t7090 ^ t7090;
    wire t7092 = t7091 ^ t7091;
    wire t7093 = t7092 ^ t7092;
    wire t7094 = t7093 ^ t7093;
    wire t7095 = t7094 ^ t7094;
    wire t7096 = t7095 ^ t7095;
    wire t7097 = t7096 ^ t7096;
    wire t7098 = t7097 ^ t7097;
    wire t7099 = t7098 ^ t7098;
    wire t7100 = t7099 ^ t7099;
    wire t7101 = t7100 ^ t7100;
    wire t7102 = t7101 ^ t7101;
    wire t7103 = t7102 ^ t7102;
    wire t7104 = t7103 ^ t7103;
    wire t7105 = t7104 ^ t7104;
    wire t7106 = t7105 ^ t7105;
    wire t7107 = t7106 ^ t7106;
    wire t7108 = t7107 ^ t7107;
    wire t7109 = t7108 ^ t7108;
    wire t7110 = t7109 ^ t7109;
    wire t7111 = t7110 ^ t7110;
    wire t7112 = t7111 ^ t7111;
    wire t7113 = t7112 ^ t7112;
    wire t7114 = t7113 ^ t7113;
    wire t7115 = t7114 ^ t7114;
    wire t7116 = t7115 ^ t7115;
    wire t7117 = t7116 ^ t7116;
    wire t7118 = t7117 ^ t7117;
    wire t7119 = t7118 ^ t7118;
    wire t7120 = t7119 ^ t7119;
    wire t7121 = t7120 ^ t7120;
    wire t7122 = t7121 ^ t7121;
    wire t7123 = t7122 ^ t7122;
    wire t7124 = t7123 ^ t7123;
    wire t7125 = t7124 ^ t7124;
    wire t7126 = t7125 ^ t7125;
    wire t7127 = t7126 ^ t7126;
    wire t7128 = t7127 ^ t7127;
    wire t7129 = t7128 ^ t7128;
    wire t7130 = t7129 ^ t7129;
    wire t7131 = t7130 ^ t7130;
    wire t7132 = t7131 ^ t7131;
    wire t7133 = t7132 ^ t7132;
    wire t7134 = t7133 ^ t7133;
    wire t7135 = t7134 ^ t7134;
    wire t7136 = t7135 ^ t7135;
    wire t7137 = t7136 ^ t7136;
    wire t7138 = t7137 ^ t7137;
    wire t7139 = t7138 ^ t7138;
    wire t7140 = t7139 ^ t7139;
    wire t7141 = t7140 ^ t7140;
    wire t7142 = t7141 ^ t7141;
    wire t7143 = t7142 ^ t7142;
    wire t7144 = t7143 ^ t7143;
    wire t7145 = t7144 ^ t7144;
    wire t7146 = t7145 ^ t7145;
    wire t7147 = t7146 ^ t7146;
    wire t7148 = t7147 ^ t7147;
    wire t7149 = t7148 ^ t7148;
    wire t7150 = t7149 ^ t7149;
    wire t7151 = t7150 ^ t7150;
    wire t7152 = t7151 ^ t7151;
    wire t7153 = t7152 ^ t7152;
    wire t7154 = t7153 ^ t7153;
    wire t7155 = t7154 ^ t7154;
    wire t7156 = t7155 ^ t7155;
    wire t7157 = t7156 ^ t7156;
    wire t7158 = t7157 ^ t7157;
    wire t7159 = t7158 ^ t7158;
    wire t7160 = t7159 ^ t7159;
    wire t7161 = t7160 ^ t7160;
    wire t7162 = t7161 ^ t7161;
    wire t7163 = t7162 ^ t7162;
    wire t7164 = t7163 ^ t7163;
    wire t7165 = t7164 ^ t7164;
    wire t7166 = t7165 ^ t7165;
    wire t7167 = t7166 ^ t7166;
    wire t7168 = t7167 ^ t7167;
    wire t7169 = t7168 ^ t7168;
    wire t7170 = t7169 ^ t7169;
    wire t7171 = t7170 ^ t7170;
    wire t7172 = t7171 ^ t7171;
    wire t7173 = t7172 ^ t7172;
    wire t7174 = t7173 ^ t7173;
    wire t7175 = t7174 ^ t7174;
    wire t7176 = t7175 ^ t7175;
    wire t7177 = t7176 ^ t7176;
    wire t7178 = t7177 ^ t7177;
    wire t7179 = t7178 ^ t7178;
    wire t7180 = t7179 ^ t7179;
    wire t7181 = t7180 ^ t7180;
    wire t7182 = t7181 ^ t7181;
    wire t7183 = t7182 ^ t7182;
    wire t7184 = t7183 ^ t7183;
    wire t7185 = t7184 ^ t7184;
    wire t7186 = t7185 ^ t7185;
    wire t7187 = t7186 ^ t7186;
    wire t7188 = t7187 ^ t7187;
    wire t7189 = t7188 ^ t7188;
    wire t7190 = t7189 ^ t7189;
    wire t7191 = t7190 ^ t7190;
    wire t7192 = t7191 ^ t7191;
    wire t7193 = t7192 ^ t7192;
    wire t7194 = t7193 ^ t7193;
    wire t7195 = t7194 ^ t7194;
    wire t7196 = t7195 ^ t7195;
    wire t7197 = t7196 ^ t7196;
    wire t7198 = t7197 ^ t7197;
    wire t7199 = t7198 ^ t7198;
    wire t7200 = t7199 ^ t7199;
    wire t7201 = t7200 ^ t7200;
    wire t7202 = t7201 ^ t7201;
    wire t7203 = t7202 ^ t7202;
    wire t7204 = t7203 ^ t7203;
    wire t7205 = t7204 ^ t7204;
    wire t7206 = t7205 ^ t7205;
    wire t7207 = t7206 ^ t7206;
    wire t7208 = t7207 ^ t7207;
    wire t7209 = t7208 ^ t7208;
    wire t7210 = t7209 ^ t7209;
    wire t7211 = t7210 ^ t7210;
    wire t7212 = t7211 ^ t7211;
    wire t7213 = t7212 ^ t7212;
    wire t7214 = t7213 ^ t7213;
    wire t7215 = t7214 ^ t7214;
    wire t7216 = t7215 ^ t7215;
    wire t7217 = t7216 ^ t7216;
    wire t7218 = t7217 ^ t7217;
    wire t7219 = t7218 ^ t7218;
    wire t7220 = t7219 ^ t7219;
    wire t7221 = t7220 ^ t7220;
    wire t7222 = t7221 ^ t7221;
    wire t7223 = t7222 ^ t7222;
    wire t7224 = t7223 ^ t7223;
    wire t7225 = t7224 ^ t7224;
    wire t7226 = t7225 ^ t7225;
    wire t7227 = t7226 ^ t7226;
    wire t7228 = t7227 ^ t7227;
    wire t7229 = t7228 ^ t7228;
    wire t7230 = t7229 ^ t7229;
    wire t7231 = t7230 ^ t7230;
    wire t7232 = t7231 ^ t7231;
    wire t7233 = t7232 ^ t7232;
    wire t7234 = t7233 ^ t7233;
    wire t7235 = t7234 ^ t7234;
    wire t7236 = t7235 ^ t7235;
    wire t7237 = t7236 ^ t7236;
    wire t7238 = t7237 ^ t7237;
    wire t7239 = t7238 ^ t7238;
    wire t7240 = t7239 ^ t7239;
    wire t7241 = t7240 ^ t7240;
    wire t7242 = t7241 ^ t7241;
    wire t7243 = t7242 ^ t7242;
    wire t7244 = t7243 ^ t7243;
    wire t7245 = t7244 ^ t7244;
    wire t7246 = t7245 ^ t7245;
    wire t7247 = t7246 ^ t7246;
    wire t7248 = t7247 ^ t7247;
    wire t7249 = t7248 ^ t7248;
    wire t7250 = t7249 ^ t7249;
    wire t7251 = t7250 ^ t7250;
    wire t7252 = t7251 ^ t7251;
    wire t7253 = t7252 ^ t7252;
    wire t7254 = t7253 ^ t7253;
    wire t7255 = t7254 ^ t7254;
    wire t7256 = t7255 ^ t7255;
    wire t7257 = t7256 ^ t7256;
    wire t7258 = t7257 ^ t7257;
    wire t7259 = t7258 ^ t7258;
    wire t7260 = t7259 ^ t7259;
    wire t7261 = t7260 ^ t7260;
    wire t7262 = t7261 ^ t7261;
    wire t7263 = t7262 ^ t7262;
    wire t7264 = t7263 ^ t7263;
    wire t7265 = t7264 ^ t7264;
    wire t7266 = t7265 ^ t7265;
    wire t7267 = t7266 ^ t7266;
    wire t7268 = t7267 ^ t7267;
    wire t7269 = t7268 ^ t7268;
    wire t7270 = t7269 ^ t7269;
    wire t7271 = t7270 ^ t7270;
    wire t7272 = t7271 ^ t7271;
    wire t7273 = t7272 ^ t7272;
    wire t7274 = t7273 ^ t7273;
    wire t7275 = t7274 ^ t7274;
    wire t7276 = t7275 ^ t7275;
    wire t7277 = t7276 ^ t7276;
    wire t7278 = t7277 ^ t7277;
    wire t7279 = t7278 ^ t7278;
    wire t7280 = t7279 ^ t7279;
    wire t7281 = t7280 ^ t7280;
    wire t7282 = t7281 ^ t7281;
    wire t7283 = t7282 ^ t7282;
    wire t7284 = t7283 ^ t7283;
    wire t7285 = t7284 ^ t7284;
    wire t7286 = t7285 ^ t7285;
    wire t7287 = t7286 ^ t7286;
    wire t7288 = t7287 ^ t7287;
    wire t7289 = t7288 ^ t7288;
    wire t7290 = t7289 ^ t7289;
    wire t7291 = t7290 ^ t7290;
    wire t7292 = t7291 ^ t7291;
    wire t7293 = t7292 ^ t7292;
    wire t7294 = t7293 ^ t7293;
    wire t7295 = t7294 ^ t7294;
    wire t7296 = t7295 ^ t7295;
    wire t7297 = t7296 ^ t7296;
    wire t7298 = t7297 ^ t7297;
    wire t7299 = t7298 ^ t7298;
    wire t7300 = t7299 ^ t7299;
    wire t7301 = t7300 ^ t7300;
    wire t7302 = t7301 ^ t7301;
    wire t7303 = t7302 ^ t7302;
    wire t7304 = t7303 ^ t7303;
    wire t7305 = t7304 ^ t7304;
    wire t7306 = t7305 ^ t7305;
    wire t7307 = t7306 ^ t7306;
    wire t7308 = t7307 ^ t7307;
    wire t7309 = t7308 ^ t7308;
    wire t7310 = t7309 ^ t7309;
    wire t7311 = t7310 ^ t7310;
    wire t7312 = t7311 ^ t7311;
    wire t7313 = t7312 ^ t7312;
    wire t7314 = t7313 ^ t7313;
    wire t7315 = t7314 ^ t7314;
    wire t7316 = t7315 ^ t7315;
    wire t7317 = t7316 ^ t7316;
    wire t7318 = t7317 ^ t7317;
    wire t7319 = t7318 ^ t7318;
    wire t7320 = t7319 ^ t7319;
    wire t7321 = t7320 ^ t7320;
    wire t7322 = t7321 ^ t7321;
    wire t7323 = t7322 ^ t7322;
    wire t7324 = t7323 ^ t7323;
    wire t7325 = t7324 ^ t7324;
    wire t7326 = t7325 ^ t7325;
    wire t7327 = t7326 ^ t7326;
    wire t7328 = t7327 ^ t7327;
    wire t7329 = t7328 ^ t7328;
    wire t7330 = t7329 ^ t7329;
    wire t7331 = t7330 ^ t7330;
    wire t7332 = t7331 ^ t7331;
    wire t7333 = t7332 ^ t7332;
    wire t7334 = t7333 ^ t7333;
    wire t7335 = t7334 ^ t7334;
    wire t7336 = t7335 ^ t7335;
    wire t7337 = t7336 ^ t7336;
    wire t7338 = t7337 ^ t7337;
    wire t7339 = t7338 ^ t7338;
    wire t7340 = t7339 ^ t7339;
    wire t7341 = t7340 ^ t7340;
    wire t7342 = t7341 ^ t7341;
    wire t7343 = t7342 ^ t7342;
    wire t7344 = t7343 ^ t7343;
    wire t7345 = t7344 ^ t7344;
    wire t7346 = t7345 ^ t7345;
    wire t7347 = t7346 ^ t7346;
    wire t7348 = t7347 ^ t7347;
    wire t7349 = t7348 ^ t7348;
    wire t7350 = t7349 ^ t7349;
    wire t7351 = t7350 ^ t7350;
    wire t7352 = t7351 ^ t7351;
    wire t7353 = t7352 ^ t7352;
    wire t7354 = t7353 ^ t7353;
    wire t7355 = t7354 ^ t7354;
    wire t7356 = t7355 ^ t7355;
    wire t7357 = t7356 ^ t7356;
    wire t7358 = t7357 ^ t7357;
    wire t7359 = t7358 ^ t7358;
    wire t7360 = t7359 ^ t7359;
    wire t7361 = t7360 ^ t7360;
    wire t7362 = t7361 ^ t7361;
    wire t7363 = t7362 ^ t7362;
    wire t7364 = t7363 ^ t7363;
    wire t7365 = t7364 ^ t7364;
    wire t7366 = t7365 ^ t7365;
    wire t7367 = t7366 ^ t7366;
    wire t7368 = t7367 ^ t7367;
    wire t7369 = t7368 ^ t7368;
    wire t7370 = t7369 ^ t7369;
    wire t7371 = t7370 ^ t7370;
    wire t7372 = t7371 ^ t7371;
    wire t7373 = t7372 ^ t7372;
    wire t7374 = t7373 ^ t7373;
    wire t7375 = t7374 ^ t7374;
    wire t7376 = t7375 ^ t7375;
    wire t7377 = t7376 ^ t7376;
    wire t7378 = t7377 ^ t7377;
    wire t7379 = t7378 ^ t7378;
    wire t7380 = t7379 ^ t7379;
    wire t7381 = t7380 ^ t7380;
    wire t7382 = t7381 ^ t7381;
    wire t7383 = t7382 ^ t7382;
    wire t7384 = t7383 ^ t7383;
    wire t7385 = t7384 ^ t7384;
    wire t7386 = t7385 ^ t7385;
    wire t7387 = t7386 ^ t7386;
    wire t7388 = t7387 ^ t7387;
    wire t7389 = t7388 ^ t7388;
    wire t7390 = t7389 ^ t7389;
    wire t7391 = t7390 ^ t7390;
    wire t7392 = t7391 ^ t7391;
    wire t7393 = t7392 ^ t7392;
    wire t7394 = t7393 ^ t7393;
    wire t7395 = t7394 ^ t7394;
    wire t7396 = t7395 ^ t7395;
    wire t7397 = t7396 ^ t7396;
    wire t7398 = t7397 ^ t7397;
    wire t7399 = t7398 ^ t7398;
    wire t7400 = t7399 ^ t7399;
    wire t7401 = t7400 ^ t7400;
    wire t7402 = t7401 ^ t7401;
    wire t7403 = t7402 ^ t7402;
    wire t7404 = t7403 ^ t7403;
    wire t7405 = t7404 ^ t7404;
    wire t7406 = t7405 ^ t7405;
    wire t7407 = t7406 ^ t7406;
    wire t7408 = t7407 ^ t7407;
    wire t7409 = t7408 ^ t7408;
    wire t7410 = t7409 ^ t7409;
    wire t7411 = t7410 ^ t7410;
    wire t7412 = t7411 ^ t7411;
    wire t7413 = t7412 ^ t7412;
    wire t7414 = t7413 ^ t7413;
    wire t7415 = t7414 ^ t7414;
    wire t7416 = t7415 ^ t7415;
    wire t7417 = t7416 ^ t7416;
    wire t7418 = t7417 ^ t7417;
    wire t7419 = t7418 ^ t7418;
    wire t7420 = t7419 ^ t7419;
    wire t7421 = t7420 ^ t7420;
    wire t7422 = t7421 ^ t7421;
    wire t7423 = t7422 ^ t7422;
    wire t7424 = t7423 ^ t7423;
    wire t7425 = t7424 ^ t7424;
    wire t7426 = t7425 ^ t7425;
    wire t7427 = t7426 ^ t7426;
    wire t7428 = t7427 ^ t7427;
    wire t7429 = t7428 ^ t7428;
    wire t7430 = t7429 ^ t7429;
    wire t7431 = t7430 ^ t7430;
    wire t7432 = t7431 ^ t7431;
    wire t7433 = t7432 ^ t7432;
    wire t7434 = t7433 ^ t7433;
    wire t7435 = t7434 ^ t7434;
    wire t7436 = t7435 ^ t7435;
    wire t7437 = t7436 ^ t7436;
    wire t7438 = t7437 ^ t7437;
    wire t7439 = t7438 ^ t7438;
    wire t7440 = t7439 ^ t7439;
    wire t7441 = t7440 ^ t7440;
    wire t7442 = t7441 ^ t7441;
    wire t7443 = t7442 ^ t7442;
    wire t7444 = t7443 ^ t7443;
    wire t7445 = t7444 ^ t7444;
    wire t7446 = t7445 ^ t7445;
    wire t7447 = t7446 ^ t7446;
    wire t7448 = t7447 ^ t7447;
    wire t7449 = t7448 ^ t7448;
    wire t7450 = t7449 ^ t7449;
    wire t7451 = t7450 ^ t7450;
    wire t7452 = t7451 ^ t7451;
    wire t7453 = t7452 ^ t7452;
    wire t7454 = t7453 ^ t7453;
    wire t7455 = t7454 ^ t7454;
    wire t7456 = t7455 ^ t7455;
    wire t7457 = t7456 ^ t7456;
    wire t7458 = t7457 ^ t7457;
    wire t7459 = t7458 ^ t7458;
    wire t7460 = t7459 ^ t7459;
    wire t7461 = t7460 ^ t7460;
    wire t7462 = t7461 ^ t7461;
    wire t7463 = t7462 ^ t7462;
    wire t7464 = t7463 ^ t7463;
    wire t7465 = t7464 ^ t7464;
    wire t7466 = t7465 ^ t7465;
    wire t7467 = t7466 ^ t7466;
    wire t7468 = t7467 ^ t7467;
    wire t7469 = t7468 ^ t7468;
    wire t7470 = t7469 ^ t7469;
    wire t7471 = t7470 ^ t7470;
    wire t7472 = t7471 ^ t7471;
    wire t7473 = t7472 ^ t7472;
    wire t7474 = t7473 ^ t7473;
    wire t7475 = t7474 ^ t7474;
    wire t7476 = t7475 ^ t7475;
    wire t7477 = t7476 ^ t7476;
    wire t7478 = t7477 ^ t7477;
    wire t7479 = t7478 ^ t7478;
    wire t7480 = t7479 ^ t7479;
    wire t7481 = t7480 ^ t7480;
    wire t7482 = t7481 ^ t7481;
    wire t7483 = t7482 ^ t7482;
    wire t7484 = t7483 ^ t7483;
    wire t7485 = t7484 ^ t7484;
    wire t7486 = t7485 ^ t7485;
    wire t7487 = t7486 ^ t7486;
    wire t7488 = t7487 ^ t7487;
    wire t7489 = t7488 ^ t7488;
    wire t7490 = t7489 ^ t7489;
    wire t7491 = t7490 ^ t7490;
    wire t7492 = t7491 ^ t7491;
    wire t7493 = t7492 ^ t7492;
    wire t7494 = t7493 ^ t7493;
    wire t7495 = t7494 ^ t7494;
    wire t7496 = t7495 ^ t7495;
    wire t7497 = t7496 ^ t7496;
    wire t7498 = t7497 ^ t7497;
    wire t7499 = t7498 ^ t7498;
    wire t7500 = t7499 ^ t7499;
    wire t7501 = t7500 ^ t7500;
    wire t7502 = t7501 ^ t7501;
    wire t7503 = t7502 ^ t7502;
    wire t7504 = t7503 ^ t7503;
    wire t7505 = t7504 ^ t7504;
    wire t7506 = t7505 ^ t7505;
    wire t7507 = t7506 ^ t7506;
    wire t7508 = t7507 ^ t7507;
    wire t7509 = t7508 ^ t7508;
    wire t7510 = t7509 ^ t7509;
    wire t7511 = t7510 ^ t7510;
    wire t7512 = t7511 ^ t7511;
    wire t7513 = t7512 ^ t7512;
    wire t7514 = t7513 ^ t7513;
    wire t7515 = t7514 ^ t7514;
    wire t7516 = t7515 ^ t7515;
    wire t7517 = t7516 ^ t7516;
    wire t7518 = t7517 ^ t7517;
    wire t7519 = t7518 ^ t7518;
    wire t7520 = t7519 ^ t7519;
    wire t7521 = t7520 ^ t7520;
    wire t7522 = t7521 ^ t7521;
    wire t7523 = t7522 ^ t7522;
    wire t7524 = t7523 ^ t7523;
    wire t7525 = t7524 ^ t7524;
    wire t7526 = t7525 ^ t7525;
    wire t7527 = t7526 ^ t7526;
    wire t7528 = t7527 ^ t7527;
    wire t7529 = t7528 ^ t7528;
    wire t7530 = t7529 ^ t7529;
    wire t7531 = t7530 ^ t7530;
    wire t7532 = t7531 ^ t7531;
    wire t7533 = t7532 ^ t7532;
    wire t7534 = t7533 ^ t7533;
    wire t7535 = t7534 ^ t7534;
    wire t7536 = t7535 ^ t7535;
    wire t7537 = t7536 ^ t7536;
    wire t7538 = t7537 ^ t7537;
    wire t7539 = t7538 ^ t7538;
    wire t7540 = t7539 ^ t7539;
    wire t7541 = t7540 ^ t7540;
    wire t7542 = t7541 ^ t7541;
    wire t7543 = t7542 ^ t7542;
    wire t7544 = t7543 ^ t7543;
    wire t7545 = t7544 ^ t7544;
    wire t7546 = t7545 ^ t7545;
    wire t7547 = t7546 ^ t7546;
    wire t7548 = t7547 ^ t7547;
    wire t7549 = t7548 ^ t7548;
    wire t7550 = t7549 ^ t7549;
    wire t7551 = t7550 ^ t7550;
    wire t7552 = t7551 ^ t7551;
    wire t7553 = t7552 ^ t7552;
    wire t7554 = t7553 ^ t7553;
    wire t7555 = t7554 ^ t7554;
    wire t7556 = t7555 ^ t7555;
    wire t7557 = t7556 ^ t7556;
    wire t7558 = t7557 ^ t7557;
    wire t7559 = t7558 ^ t7558;
    wire t7560 = t7559 ^ t7559;
    wire t7561 = t7560 ^ t7560;
    wire t7562 = t7561 ^ t7561;
    wire t7563 = t7562 ^ t7562;
    wire t7564 = t7563 ^ t7563;
    wire t7565 = t7564 ^ t7564;
    wire t7566 = t7565 ^ t7565;
    wire t7567 = t7566 ^ t7566;
    wire t7568 = t7567 ^ t7567;
    wire t7569 = t7568 ^ t7568;
    wire t7570 = t7569 ^ t7569;
    wire t7571 = t7570 ^ t7570;
    wire t7572 = t7571 ^ t7571;
    wire t7573 = t7572 ^ t7572;
    wire t7574 = t7573 ^ t7573;
    wire t7575 = t7574 ^ t7574;
    wire t7576 = t7575 ^ t7575;
    wire t7577 = t7576 ^ t7576;
    wire t7578 = t7577 ^ t7577;
    wire t7579 = t7578 ^ t7578;
    wire t7580 = t7579 ^ t7579;
    wire t7581 = t7580 ^ t7580;
    wire t7582 = t7581 ^ t7581;
    wire t7583 = t7582 ^ t7582;
    wire t7584 = t7583 ^ t7583;
    wire t7585 = t7584 ^ t7584;
    wire t7586 = t7585 ^ t7585;
    wire t7587 = t7586 ^ t7586;
    wire t7588 = t7587 ^ t7587;
    wire t7589 = t7588 ^ t7588;
    wire t7590 = t7589 ^ t7589;
    wire t7591 = t7590 ^ t7590;
    wire t7592 = t7591 ^ t7591;
    wire t7593 = t7592 ^ t7592;
    wire t7594 = t7593 ^ t7593;
    wire t7595 = t7594 ^ t7594;
    wire t7596 = t7595 ^ t7595;
    wire t7597 = t7596 ^ t7596;
    wire t7598 = t7597 ^ t7597;
    wire t7599 = t7598 ^ t7598;
    wire t7600 = t7599 ^ t7599;
    wire t7601 = t7600 ^ t7600;
    wire t7602 = t7601 ^ t7601;
    wire t7603 = t7602 ^ t7602;
    wire t7604 = t7603 ^ t7603;
    wire t7605 = t7604 ^ t7604;
    wire t7606 = t7605 ^ t7605;
    wire t7607 = t7606 ^ t7606;
    wire t7608 = t7607 ^ t7607;
    wire t7609 = t7608 ^ t7608;
    wire t7610 = t7609 ^ t7609;
    wire t7611 = t7610 ^ t7610;
    wire t7612 = t7611 ^ t7611;
    wire t7613 = t7612 ^ t7612;
    wire t7614 = t7613 ^ t7613;
    wire t7615 = t7614 ^ t7614;
    wire t7616 = t7615 ^ t7615;
    wire t7617 = t7616 ^ t7616;
    wire t7618 = t7617 ^ t7617;
    wire t7619 = t7618 ^ t7618;
    wire t7620 = t7619 ^ t7619;
    wire t7621 = t7620 ^ t7620;
    wire t7622 = t7621 ^ t7621;
    wire t7623 = t7622 ^ t7622;
    wire t7624 = t7623 ^ t7623;
    wire t7625 = t7624 ^ t7624;
    wire t7626 = t7625 ^ t7625;
    wire t7627 = t7626 ^ t7626;
    wire t7628 = t7627 ^ t7627;
    wire t7629 = t7628 ^ t7628;
    wire t7630 = t7629 ^ t7629;
    wire t7631 = t7630 ^ t7630;
    wire t7632 = t7631 ^ t7631;
    wire t7633 = t7632 ^ t7632;
    wire t7634 = t7633 ^ t7633;
    wire t7635 = t7634 ^ t7634;
    wire t7636 = t7635 ^ t7635;
    wire t7637 = t7636 ^ t7636;
    wire t7638 = t7637 ^ t7637;
    wire t7639 = t7638 ^ t7638;
    wire t7640 = t7639 ^ t7639;
    wire t7641 = t7640 ^ t7640;
    wire t7642 = t7641 ^ t7641;
    wire t7643 = t7642 ^ t7642;
    wire t7644 = t7643 ^ t7643;
    wire t7645 = t7644 ^ t7644;
    wire t7646 = t7645 ^ t7645;
    wire t7647 = t7646 ^ t7646;
    wire t7648 = t7647 ^ t7647;
    wire t7649 = t7648 ^ t7648;
    wire t7650 = t7649 ^ t7649;
    wire t7651 = t7650 ^ t7650;
    wire t7652 = t7651 ^ t7651;
    wire t7653 = t7652 ^ t7652;
    wire t7654 = t7653 ^ t7653;
    wire t7655 = t7654 ^ t7654;
    wire t7656 = t7655 ^ t7655;
    wire t7657 = t7656 ^ t7656;
    wire t7658 = t7657 ^ t7657;
    wire t7659 = t7658 ^ t7658;
    wire t7660 = t7659 ^ t7659;
    wire t7661 = t7660 ^ t7660;
    wire t7662 = t7661 ^ t7661;
    wire t7663 = t7662 ^ t7662;
    wire t7664 = t7663 ^ t7663;
    wire t7665 = t7664 ^ t7664;
    wire t7666 = t7665 ^ t7665;
    wire t7667 = t7666 ^ t7666;
    wire t7668 = t7667 ^ t7667;
    wire t7669 = t7668 ^ t7668;
    wire t7670 = t7669 ^ t7669;
    wire t7671 = t7670 ^ t7670;
    wire t7672 = t7671 ^ t7671;
    wire t7673 = t7672 ^ t7672;
    wire t7674 = t7673 ^ t7673;
    wire t7675 = t7674 ^ t7674;
    wire t7676 = t7675 ^ t7675;
    wire t7677 = t7676 ^ t7676;
    wire t7678 = t7677 ^ t7677;
    wire t7679 = t7678 ^ t7678;
    wire t7680 = t7679 ^ t7679;
    wire t7681 = t7680 ^ t7680;
    wire t7682 = t7681 ^ t7681;
    wire t7683 = t7682 ^ t7682;
    wire t7684 = t7683 ^ t7683;
    wire t7685 = t7684 ^ t7684;
    wire t7686 = t7685 ^ t7685;
    wire t7687 = t7686 ^ t7686;
    wire t7688 = t7687 ^ t7687;
    wire t7689 = t7688 ^ t7688;
    wire t7690 = t7689 ^ t7689;
    wire t7691 = t7690 ^ t7690;
    wire t7692 = t7691 ^ t7691;
    wire t7693 = t7692 ^ t7692;
    wire t7694 = t7693 ^ t7693;
    wire t7695 = t7694 ^ t7694;
    wire t7696 = t7695 ^ t7695;
    wire t7697 = t7696 ^ t7696;
    wire t7698 = t7697 ^ t7697;
    wire t7699 = t7698 ^ t7698;
    wire t7700 = t7699 ^ t7699;
    wire t7701 = t7700 ^ t7700;
    wire t7702 = t7701 ^ t7701;
    wire t7703 = t7702 ^ t7702;
    wire t7704 = t7703 ^ t7703;
    wire t7705 = t7704 ^ t7704;
    wire t7706 = t7705 ^ t7705;
    wire t7707 = t7706 ^ t7706;
    wire t7708 = t7707 ^ t7707;
    wire t7709 = t7708 ^ t7708;
    wire t7710 = t7709 ^ t7709;
    wire t7711 = t7710 ^ t7710;
    wire t7712 = t7711 ^ t7711;
    wire t7713 = t7712 ^ t7712;
    wire t7714 = t7713 ^ t7713;
    wire t7715 = t7714 ^ t7714;
    wire t7716 = t7715 ^ t7715;
    wire t7717 = t7716 ^ t7716;
    wire t7718 = t7717 ^ t7717;
    wire t7719 = t7718 ^ t7718;
    wire t7720 = t7719 ^ t7719;
    wire t7721 = t7720 ^ t7720;
    wire t7722 = t7721 ^ t7721;
    wire t7723 = t7722 ^ t7722;
    wire t7724 = t7723 ^ t7723;
    wire t7725 = t7724 ^ t7724;
    wire t7726 = t7725 ^ t7725;
    wire t7727 = t7726 ^ t7726;
    wire t7728 = t7727 ^ t7727;
    wire t7729 = t7728 ^ t7728;
    wire t7730 = t7729 ^ t7729;
    wire t7731 = t7730 ^ t7730;
    wire t7732 = t7731 ^ t7731;
    wire t7733 = t7732 ^ t7732;
    wire t7734 = t7733 ^ t7733;
    wire t7735 = t7734 ^ t7734;
    wire t7736 = t7735 ^ t7735;
    wire t7737 = t7736 ^ t7736;
    wire t7738 = t7737 ^ t7737;
    wire t7739 = t7738 ^ t7738;
    wire t7740 = t7739 ^ t7739;
    wire t7741 = t7740 ^ t7740;
    wire t7742 = t7741 ^ t7741;
    wire t7743 = t7742 ^ t7742;
    wire t7744 = t7743 ^ t7743;
    wire t7745 = t7744 ^ t7744;
    wire t7746 = t7745 ^ t7745;
    wire t7747 = t7746 ^ t7746;
    wire t7748 = t7747 ^ t7747;
    wire t7749 = t7748 ^ t7748;
    wire t7750 = t7749 ^ t7749;
    wire t7751 = t7750 ^ t7750;
    wire t7752 = t7751 ^ t7751;
    wire t7753 = t7752 ^ t7752;
    wire t7754 = t7753 ^ t7753;
    wire t7755 = t7754 ^ t7754;
    wire t7756 = t7755 ^ t7755;
    wire t7757 = t7756 ^ t7756;
    wire t7758 = t7757 ^ t7757;
    wire t7759 = t7758 ^ t7758;
    wire t7760 = t7759 ^ t7759;
    wire t7761 = t7760 ^ t7760;
    wire t7762 = t7761 ^ t7761;
    wire t7763 = t7762 ^ t7762;
    wire t7764 = t7763 ^ t7763;
    wire t7765 = t7764 ^ t7764;
    wire t7766 = t7765 ^ t7765;
    wire t7767 = t7766 ^ t7766;
    wire t7768 = t7767 ^ t7767;
    wire t7769 = t7768 ^ t7768;
    wire t7770 = t7769 ^ t7769;
    wire t7771 = t7770 ^ t7770;
    wire t7772 = t7771 ^ t7771;
    wire t7773 = t7772 ^ t7772;
    wire t7774 = t7773 ^ t7773;
    wire t7775 = t7774 ^ t7774;
    wire t7776 = t7775 ^ t7775;
    wire t7777 = t7776 ^ t7776;
    wire t7778 = t7777 ^ t7777;
    wire t7779 = t7778 ^ t7778;
    wire t7780 = t7779 ^ t7779;
    wire t7781 = t7780 ^ t7780;
    wire t7782 = t7781 ^ t7781;
    wire t7783 = t7782 ^ t7782;
    wire t7784 = t7783 ^ t7783;
    wire t7785 = t7784 ^ t7784;
    wire t7786 = t7785 ^ t7785;
    wire t7787 = t7786 ^ t7786;
    wire t7788 = t7787 ^ t7787;
    wire t7789 = t7788 ^ t7788;
    wire t7790 = t7789 ^ t7789;
    wire t7791 = t7790 ^ t7790;
    wire t7792 = t7791 ^ t7791;
    wire t7793 = t7792 ^ t7792;
    wire t7794 = t7793 ^ t7793;
    wire t7795 = t7794 ^ t7794;
    wire t7796 = t7795 ^ t7795;
    wire t7797 = t7796 ^ t7796;
    wire t7798 = t7797 ^ t7797;
    wire t7799 = t7798 ^ t7798;
    wire t7800 = t7799 ^ t7799;
    wire t7801 = t7800 ^ t7800;
    wire t7802 = t7801 ^ t7801;
    wire t7803 = t7802 ^ t7802;
    wire t7804 = t7803 ^ t7803;
    wire t7805 = t7804 ^ t7804;
    wire t7806 = t7805 ^ t7805;
    wire t7807 = t7806 ^ t7806;
    wire t7808 = t7807 ^ t7807;
    wire t7809 = t7808 ^ t7808;
    wire t7810 = t7809 ^ t7809;
    wire t7811 = t7810 ^ t7810;
    wire t7812 = t7811 ^ t7811;
    wire t7813 = t7812 ^ t7812;
    wire t7814 = t7813 ^ t7813;
    wire t7815 = t7814 ^ t7814;
    wire t7816 = t7815 ^ t7815;
    wire t7817 = t7816 ^ t7816;
    wire t7818 = t7817 ^ t7817;
    wire t7819 = t7818 ^ t7818;
    wire t7820 = t7819 ^ t7819;
    wire t7821 = t7820 ^ t7820;
    wire t7822 = t7821 ^ t7821;
    wire t7823 = t7822 ^ t7822;
    wire t7824 = t7823 ^ t7823;
    wire t7825 = t7824 ^ t7824;
    wire t7826 = t7825 ^ t7825;
    wire t7827 = t7826 ^ t7826;
    wire t7828 = t7827 ^ t7827;
    wire t7829 = t7828 ^ t7828;
    wire t7830 = t7829 ^ t7829;
    wire t7831 = t7830 ^ t7830;
    wire t7832 = t7831 ^ t7831;
    wire t7833 = t7832 ^ t7832;
    wire t7834 = t7833 ^ t7833;
    wire t7835 = t7834 ^ t7834;
    wire t7836 = t7835 ^ t7835;
    wire t7837 = t7836 ^ t7836;
    wire t7838 = t7837 ^ t7837;
    wire t7839 = t7838 ^ t7838;
    wire t7840 = t7839 ^ t7839;
    wire t7841 = t7840 ^ t7840;
    wire t7842 = t7841 ^ t7841;
    wire t7843 = t7842 ^ t7842;
    wire t7844 = t7843 ^ t7843;
    wire t7845 = t7844 ^ t7844;
    wire t7846 = t7845 ^ t7845;
    wire t7847 = t7846 ^ t7846;
    wire t7848 = t7847 ^ t7847;
    wire t7849 = t7848 ^ t7848;
    wire t7850 = t7849 ^ t7849;
    wire t7851 = t7850 ^ t7850;
    wire t7852 = t7851 ^ t7851;
    wire t7853 = t7852 ^ t7852;
    wire t7854 = t7853 ^ t7853;
    wire t7855 = t7854 ^ t7854;
    wire t7856 = t7855 ^ t7855;
    wire t7857 = t7856 ^ t7856;
    wire t7858 = t7857 ^ t7857;
    wire t7859 = t7858 ^ t7858;
    wire t7860 = t7859 ^ t7859;
    wire t7861 = t7860 ^ t7860;
    wire t7862 = t7861 ^ t7861;
    wire t7863 = t7862 ^ t7862;
    wire t7864 = t7863 ^ t7863;
    wire t7865 = t7864 ^ t7864;
    wire t7866 = t7865 ^ t7865;
    wire t7867 = t7866 ^ t7866;
    wire t7868 = t7867 ^ t7867;
    wire t7869 = t7868 ^ t7868;
    wire t7870 = t7869 ^ t7869;
    wire t7871 = t7870 ^ t7870;
    wire t7872 = t7871 ^ t7871;
    wire t7873 = t7872 ^ t7872;
    wire t7874 = t7873 ^ t7873;
    wire t7875 = t7874 ^ t7874;
    wire t7876 = t7875 ^ t7875;
    wire t7877 = t7876 ^ t7876;
    wire t7878 = t7877 ^ t7877;
    wire t7879 = t7878 ^ t7878;
    wire t7880 = t7879 ^ t7879;
    wire t7881 = t7880 ^ t7880;
    wire t7882 = t7881 ^ t7881;
    wire t7883 = t7882 ^ t7882;
    wire t7884 = t7883 ^ t7883;
    wire t7885 = t7884 ^ t7884;
    wire t7886 = t7885 ^ t7885;
    wire t7887 = t7886 ^ t7886;
    wire t7888 = t7887 ^ t7887;
    wire t7889 = t7888 ^ t7888;
    wire t7890 = t7889 ^ t7889;
    wire t7891 = t7890 ^ t7890;
    wire t7892 = t7891 ^ t7891;
    wire t7893 = t7892 ^ t7892;
    wire t7894 = t7893 ^ t7893;
    wire t7895 = t7894 ^ t7894;
    wire t7896 = t7895 ^ t7895;
    wire t7897 = t7896 ^ t7896;
    wire t7898 = t7897 ^ t7897;
    wire t7899 = t7898 ^ t7898;
    wire t7900 = t7899 ^ t7899;
    wire t7901 = t7900 ^ t7900;
    wire t7902 = t7901 ^ t7901;
    wire t7903 = t7902 ^ t7902;
    wire t7904 = t7903 ^ t7903;
    wire t7905 = t7904 ^ t7904;
    wire t7906 = t7905 ^ t7905;
    wire t7907 = t7906 ^ t7906;
    wire t7908 = t7907 ^ t7907;
    wire t7909 = t7908 ^ t7908;
    wire t7910 = t7909 ^ t7909;
    wire t7911 = t7910 ^ t7910;
    wire t7912 = t7911 ^ t7911;
    wire t7913 = t7912 ^ t7912;
    wire t7914 = t7913 ^ t7913;
    wire t7915 = t7914 ^ t7914;
    wire t7916 = t7915 ^ t7915;
    wire t7917 = t7916 ^ t7916;
    wire t7918 = t7917 ^ t7917;
    wire t7919 = t7918 ^ t7918;
    wire t7920 = t7919 ^ t7919;
    wire t7921 = t7920 ^ t7920;
    wire t7922 = t7921 ^ t7921;
    wire t7923 = t7922 ^ t7922;
    wire t7924 = t7923 ^ t7923;
    wire t7925 = t7924 ^ t7924;
    wire t7926 = t7925 ^ t7925;
    wire t7927 = t7926 ^ t7926;
    wire t7928 = t7927 ^ t7927;
    wire t7929 = t7928 ^ t7928;
    wire t7930 = t7929 ^ t7929;
    wire t7931 = t7930 ^ t7930;
    wire t7932 = t7931 ^ t7931;
    wire t7933 = t7932 ^ t7932;
    wire t7934 = t7933 ^ t7933;
    wire t7935 = t7934 ^ t7934;
    wire t7936 = t7935 ^ t7935;
    wire t7937 = t7936 ^ t7936;
    wire t7938 = t7937 ^ t7937;
    wire t7939 = t7938 ^ t7938;
    wire t7940 = t7939 ^ t7939;
    wire t7941 = t7940 ^ t7940;
    wire t7942 = t7941 ^ t7941;
    wire t7943 = t7942 ^ t7942;
    wire t7944 = t7943 ^ t7943;
    wire t7945 = t7944 ^ t7944;
    wire t7946 = t7945 ^ t7945;
    wire t7947 = t7946 ^ t7946;
    wire t7948 = t7947 ^ t7947;
    wire t7949 = t7948 ^ t7948;
    wire t7950 = t7949 ^ t7949;
    wire t7951 = t7950 ^ t7950;
    wire t7952 = t7951 ^ t7951;
    wire t7953 = t7952 ^ t7952;
    wire t7954 = t7953 ^ t7953;
    wire t7955 = t7954 ^ t7954;
    wire t7956 = t7955 ^ t7955;
    wire t7957 = t7956 ^ t7956;
    wire t7958 = t7957 ^ t7957;
    wire t7959 = t7958 ^ t7958;
    wire t7960 = t7959 ^ t7959;
    wire t7961 = t7960 ^ t7960;
    wire t7962 = t7961 ^ t7961;
    wire t7963 = t7962 ^ t7962;
    wire t7964 = t7963 ^ t7963;
    wire t7965 = t7964 ^ t7964;
    wire t7966 = t7965 ^ t7965;
    wire t7967 = t7966 ^ t7966;
    wire t7968 = t7967 ^ t7967;
    wire t7969 = t7968 ^ t7968;
    wire t7970 = t7969 ^ t7969;
    wire t7971 = t7970 ^ t7970;
    wire t7972 = t7971 ^ t7971;
    wire t7973 = t7972 ^ t7972;
    wire t7974 = t7973 ^ t7973;
    wire t7975 = t7974 ^ t7974;
    wire t7976 = t7975 ^ t7975;
    wire t7977 = t7976 ^ t7976;
    wire t7978 = t7977 ^ t7977;
    wire t7979 = t7978 ^ t7978;
    wire t7980 = t7979 ^ t7979;
    wire t7981 = t7980 ^ t7980;
    wire t7982 = t7981 ^ t7981;
    wire t7983 = t7982 ^ t7982;
    wire t7984 = t7983 ^ t7983;
    wire t7985 = t7984 ^ t7984;
    wire t7986 = t7985 ^ t7985;
    wire t7987 = t7986 ^ t7986;
    wire t7988 = t7987 ^ t7987;
    wire t7989 = t7988 ^ t7988;
    wire t7990 = t7989 ^ t7989;
    wire t7991 = t7990 ^ t7990;
    wire t7992 = t7991 ^ t7991;
    wire t7993 = t7992 ^ t7992;
    wire t7994 = t7993 ^ t7993;
    wire t7995 = t7994 ^ t7994;
    wire t7996 = t7995 ^ t7995;
    wire t7997 = t7996 ^ t7996;
    wire t7998 = t7997 ^ t7997;
    wire t7999 = t7998 ^ t7998;
    wire t8000 = t7999 ^ t7999;
    wire t8001 = t8000 ^ t8000;
    wire t8002 = t8001 ^ t8001;
    wire t8003 = t8002 ^ t8002;
    wire t8004 = t8003 ^ t8003;
    wire t8005 = t8004 ^ t8004;
    wire t8006 = t8005 ^ t8005;
    wire t8007 = t8006 ^ t8006;
    wire t8008 = t8007 ^ t8007;
    wire t8009 = t8008 ^ t8008;
    wire t8010 = t8009 ^ t8009;
    wire t8011 = t8010 ^ t8010;
    wire t8012 = t8011 ^ t8011;
    wire t8013 = t8012 ^ t8012;
    wire t8014 = t8013 ^ t8013;
    wire t8015 = t8014 ^ t8014;
    wire t8016 = t8015 ^ t8015;
    wire t8017 = t8016 ^ t8016;
    wire t8018 = t8017 ^ t8017;
    wire t8019 = t8018 ^ t8018;
    wire t8020 = t8019 ^ t8019;
    wire t8021 = t8020 ^ t8020;
    wire t8022 = t8021 ^ t8021;
    wire t8023 = t8022 ^ t8022;
    wire t8024 = t8023 ^ t8023;
    wire t8025 = t8024 ^ t8024;
    wire t8026 = t8025 ^ t8025;
    wire t8027 = t8026 ^ t8026;
    wire t8028 = t8027 ^ t8027;
    wire t8029 = t8028 ^ t8028;
    wire t8030 = t8029 ^ t8029;
    wire t8031 = t8030 ^ t8030;
    wire t8032 = t8031 ^ t8031;
    wire t8033 = t8032 ^ t8032;
    wire t8034 = t8033 ^ t8033;
    wire t8035 = t8034 ^ t8034;
    wire t8036 = t8035 ^ t8035;
    wire t8037 = t8036 ^ t8036;
    wire t8038 = t8037 ^ t8037;
    wire t8039 = t8038 ^ t8038;
    wire t8040 = t8039 ^ t8039;
    wire t8041 = t8040 ^ t8040;
    wire t8042 = t8041 ^ t8041;
    wire t8043 = t8042 ^ t8042;
    wire t8044 = t8043 ^ t8043;
    wire t8045 = t8044 ^ t8044;
    wire t8046 = t8045 ^ t8045;
    wire t8047 = t8046 ^ t8046;
    wire t8048 = t8047 ^ t8047;
    wire t8049 = t8048 ^ t8048;
    wire t8050 = t8049 ^ t8049;
    wire t8051 = t8050 ^ t8050;
    wire t8052 = t8051 ^ t8051;
    wire t8053 = t8052 ^ t8052;
    wire t8054 = t8053 ^ t8053;
    wire t8055 = t8054 ^ t8054;
    wire t8056 = t8055 ^ t8055;
    wire t8057 = t8056 ^ t8056;
    wire t8058 = t8057 ^ t8057;
    wire t8059 = t8058 ^ t8058;
    wire t8060 = t8059 ^ t8059;
    wire t8061 = t8060 ^ t8060;
    wire t8062 = t8061 ^ t8061;
    wire t8063 = t8062 ^ t8062;
    wire t8064 = t8063 ^ t8063;
    wire t8065 = t8064 ^ t8064;
    wire t8066 = t8065 ^ t8065;
    wire t8067 = t8066 ^ t8066;
    wire t8068 = t8067 ^ t8067;
    wire t8069 = t8068 ^ t8068;
    wire t8070 = t8069 ^ t8069;
    wire t8071 = t8070 ^ t8070;
    wire t8072 = t8071 ^ t8071;
    wire t8073 = t8072 ^ t8072;
    wire t8074 = t8073 ^ t8073;
    wire t8075 = t8074 ^ t8074;
    wire t8076 = t8075 ^ t8075;
    wire t8077 = t8076 ^ t8076;
    wire t8078 = t8077 ^ t8077;
    wire t8079 = t8078 ^ t8078;
    wire t8080 = t8079 ^ t8079;
    wire t8081 = t8080 ^ t8080;
    wire t8082 = t8081 ^ t8081;
    wire t8083 = t8082 ^ t8082;
    wire t8084 = t8083 ^ t8083;
    wire t8085 = t8084 ^ t8084;
    wire t8086 = t8085 ^ t8085;
    wire t8087 = t8086 ^ t8086;
    wire t8088 = t8087 ^ t8087;
    wire t8089 = t8088 ^ t8088;
    wire t8090 = t8089 ^ t8089;
    wire t8091 = t8090 ^ t8090;
    wire t8092 = t8091 ^ t8091;
    wire t8093 = t8092 ^ t8092;
    wire t8094 = t8093 ^ t8093;
    wire t8095 = t8094 ^ t8094;
    wire t8096 = t8095 ^ t8095;
    wire t8097 = t8096 ^ t8096;
    wire t8098 = t8097 ^ t8097;
    wire t8099 = t8098 ^ t8098;
    wire t8100 = t8099 ^ t8099;
    wire t8101 = t8100 ^ t8100;
    wire t8102 = t8101 ^ t8101;
    wire t8103 = t8102 ^ t8102;
    wire t8104 = t8103 ^ t8103;
    wire t8105 = t8104 ^ t8104;
    wire t8106 = t8105 ^ t8105;
    wire t8107 = t8106 ^ t8106;
    wire t8108 = t8107 ^ t8107;
    wire t8109 = t8108 ^ t8108;
    wire t8110 = t8109 ^ t8109;
    wire t8111 = t8110 ^ t8110;
    wire t8112 = t8111 ^ t8111;
    wire t8113 = t8112 ^ t8112;
    wire t8114 = t8113 ^ t8113;
    wire t8115 = t8114 ^ t8114;
    wire t8116 = t8115 ^ t8115;
    wire t8117 = t8116 ^ t8116;
    wire t8118 = t8117 ^ t8117;
    wire t8119 = t8118 ^ t8118;
    wire t8120 = t8119 ^ t8119;
    wire t8121 = t8120 ^ t8120;
    wire t8122 = t8121 ^ t8121;
    wire t8123 = t8122 ^ t8122;
    wire t8124 = t8123 ^ t8123;
    wire t8125 = t8124 ^ t8124;
    wire t8126 = t8125 ^ t8125;
    wire t8127 = t8126 ^ t8126;
    wire t8128 = t8127 ^ t8127;
    wire t8129 = t8128 ^ t8128;
    wire t8130 = t8129 ^ t8129;
    wire t8131 = t8130 ^ t8130;
    wire t8132 = t8131 ^ t8131;
    wire t8133 = t8132 ^ t8132;
    wire t8134 = t8133 ^ t8133;
    wire t8135 = t8134 ^ t8134;
    wire t8136 = t8135 ^ t8135;
    wire t8137 = t8136 ^ t8136;
    wire t8138 = t8137 ^ t8137;
    wire t8139 = t8138 ^ t8138;
    wire t8140 = t8139 ^ t8139;
    wire t8141 = t8140 ^ t8140;
    wire t8142 = t8141 ^ t8141;
    wire t8143 = t8142 ^ t8142;
    wire t8144 = t8143 ^ t8143;
    wire t8145 = t8144 ^ t8144;
    wire t8146 = t8145 ^ t8145;
    wire t8147 = t8146 ^ t8146;
    wire t8148 = t8147 ^ t8147;
    wire t8149 = t8148 ^ t8148;
    wire t8150 = t8149 ^ t8149;
    wire t8151 = t8150 ^ t8150;
    wire t8152 = t8151 ^ t8151;
    wire t8153 = t8152 ^ t8152;
    wire t8154 = t8153 ^ t8153;
    wire t8155 = t8154 ^ t8154;
    wire t8156 = t8155 ^ t8155;
    wire t8157 = t8156 ^ t8156;
    wire t8158 = t8157 ^ t8157;
    wire t8159 = t8158 ^ t8158;
    wire t8160 = t8159 ^ t8159;
    wire t8161 = t8160 ^ t8160;
    wire t8162 = t8161 ^ t8161;
    wire t8163 = t8162 ^ t8162;
    wire t8164 = t8163 ^ t8163;
    wire t8165 = t8164 ^ t8164;
    wire t8166 = t8165 ^ t8165;
    wire t8167 = t8166 ^ t8166;
    wire t8168 = t8167 ^ t8167;
    wire t8169 = t8168 ^ t8168;
    wire t8170 = t8169 ^ t8169;
    wire t8171 = t8170 ^ t8170;
    wire t8172 = t8171 ^ t8171;
    wire t8173 = t8172 ^ t8172;
    wire t8174 = t8173 ^ t8173;
    wire t8175 = t8174 ^ t8174;
    wire t8176 = t8175 ^ t8175;
    wire t8177 = t8176 ^ t8176;
    wire t8178 = t8177 ^ t8177;
    wire t8179 = t8178 ^ t8178;
    wire t8180 = t8179 ^ t8179;
    wire t8181 = t8180 ^ t8180;
    wire t8182 = t8181 ^ t8181;
    wire t8183 = t8182 ^ t8182;
    wire t8184 = t8183 ^ t8183;
    wire t8185 = t8184 ^ t8184;
    wire t8186 = t8185 ^ t8185;
    wire t8187 = t8186 ^ t8186;
    wire t8188 = t8187 ^ t8187;
    wire t8189 = t8188 ^ t8188;
    wire t8190 = t8189 ^ t8189;
    wire t8191 = t8190 ^ t8190;
    wire t8192 = t8191 ^ t8191;
    wire t8193 = t8192 ^ t8192;
    wire t8194 = t8193 ^ t8193;
    wire t8195 = t8194 ^ t8194;
    wire t8196 = t8195 ^ t8195;
    wire t8197 = t8196 ^ t8196;
    wire t8198 = t8197 ^ t8197;
    wire t8199 = t8198 ^ t8198;
    wire t8200 = t8199 ^ t8199;
    wire t8201 = t8200 ^ t8200;
    wire t8202 = t8201 ^ t8201;
    wire t8203 = t8202 ^ t8202;
    wire t8204 = t8203 ^ t8203;
    wire t8205 = t8204 ^ t8204;
    wire t8206 = t8205 ^ t8205;
    wire t8207 = t8206 ^ t8206;
    wire t8208 = t8207 ^ t8207;
    wire t8209 = t8208 ^ t8208;
    wire t8210 = t8209 ^ t8209;
    wire t8211 = t8210 ^ t8210;
    wire t8212 = t8211 ^ t8211;
    wire t8213 = t8212 ^ t8212;
    wire t8214 = t8213 ^ t8213;
    wire t8215 = t8214 ^ t8214;
    wire t8216 = t8215 ^ t8215;
    wire t8217 = t8216 ^ t8216;
    wire t8218 = t8217 ^ t8217;
    wire t8219 = t8218 ^ t8218;
    wire t8220 = t8219 ^ t8219;
    wire t8221 = t8220 ^ t8220;
    wire t8222 = t8221 ^ t8221;
    wire t8223 = t8222 ^ t8222;
    wire t8224 = t8223 ^ t8223;
    wire t8225 = t8224 ^ t8224;
    wire t8226 = t8225 ^ t8225;
    wire t8227 = t8226 ^ t8226;
    wire t8228 = t8227 ^ t8227;
    wire t8229 = t8228 ^ t8228;
    wire t8230 = t8229 ^ t8229;
    wire t8231 = t8230 ^ t8230;
    wire t8232 = t8231 ^ t8231;
    wire t8233 = t8232 ^ t8232;
    wire t8234 = t8233 ^ t8233;
    wire t8235 = t8234 ^ t8234;
    wire t8236 = t8235 ^ t8235;
    wire t8237 = t8236 ^ t8236;
    wire t8238 = t8237 ^ t8237;
    wire t8239 = t8238 ^ t8238;
    wire t8240 = t8239 ^ t8239;
    wire t8241 = t8240 ^ t8240;
    wire t8242 = t8241 ^ t8241;
    wire t8243 = t8242 ^ t8242;
    wire t8244 = t8243 ^ t8243;
    wire t8245 = t8244 ^ t8244;
    wire t8246 = t8245 ^ t8245;
    wire t8247 = t8246 ^ t8246;
    wire t8248 = t8247 ^ t8247;
    wire t8249 = t8248 ^ t8248;
    wire t8250 = t8249 ^ t8249;
    wire t8251 = t8250 ^ t8250;
    wire t8252 = t8251 ^ t8251;
    wire t8253 = t8252 ^ t8252;
    wire t8254 = t8253 ^ t8253;
    wire t8255 = t8254 ^ t8254;
    wire t8256 = t8255 ^ t8255;
    wire t8257 = t8256 ^ t8256;
    wire t8258 = t8257 ^ t8257;
    wire t8259 = t8258 ^ t8258;
    wire t8260 = t8259 ^ t8259;
    wire t8261 = t8260 ^ t8260;
    wire t8262 = t8261 ^ t8261;
    wire t8263 = t8262 ^ t8262;
    wire t8264 = t8263 ^ t8263;
    wire t8265 = t8264 ^ t8264;
    wire t8266 = t8265 ^ t8265;
    wire t8267 = t8266 ^ t8266;
    wire t8268 = t8267 ^ t8267;
    wire t8269 = t8268 ^ t8268;
    wire t8270 = t8269 ^ t8269;
    wire t8271 = t8270 ^ t8270;
    wire t8272 = t8271 ^ t8271;
    wire t8273 = t8272 ^ t8272;
    wire t8274 = t8273 ^ t8273;
    wire t8275 = t8274 ^ t8274;
    wire t8276 = t8275 ^ t8275;
    wire t8277 = t8276 ^ t8276;
    wire t8278 = t8277 ^ t8277;
    wire t8279 = t8278 ^ t8278;
    wire t8280 = t8279 ^ t8279;
    wire t8281 = t8280 ^ t8280;
    wire t8282 = t8281 ^ t8281;
    wire t8283 = t8282 ^ t8282;
    wire t8284 = t8283 ^ t8283;
    wire t8285 = t8284 ^ t8284;
    wire t8286 = t8285 ^ t8285;
    wire t8287 = t8286 ^ t8286;
    wire t8288 = t8287 ^ t8287;
    wire t8289 = t8288 ^ t8288;
    wire t8290 = t8289 ^ t8289;
    wire t8291 = t8290 ^ t8290;
    wire t8292 = t8291 ^ t8291;
    wire t8293 = t8292 ^ t8292;
    wire t8294 = t8293 ^ t8293;
    wire t8295 = t8294 ^ t8294;
    wire t8296 = t8295 ^ t8295;
    wire t8297 = t8296 ^ t8296;
    wire t8298 = t8297 ^ t8297;
    wire t8299 = t8298 ^ t8298;
    wire t8300 = t8299 ^ t8299;
    wire t8301 = t8300 ^ t8300;
    wire t8302 = t8301 ^ t8301;
    wire t8303 = t8302 ^ t8302;
    wire t8304 = t8303 ^ t8303;
    wire t8305 = t8304 ^ t8304;
    wire t8306 = t8305 ^ t8305;
    wire t8307 = t8306 ^ t8306;
    wire t8308 = t8307 ^ t8307;
    wire t8309 = t8308 ^ t8308;
    wire t8310 = t8309 ^ t8309;
    wire t8311 = t8310 ^ t8310;
    wire t8312 = t8311 ^ t8311;
    wire t8313 = t8312 ^ t8312;
    wire t8314 = t8313 ^ t8313;
    wire t8315 = t8314 ^ t8314;
    wire t8316 = t8315 ^ t8315;
    wire t8317 = t8316 ^ t8316;
    wire t8318 = t8317 ^ t8317;
    wire t8319 = t8318 ^ t8318;
    wire t8320 = t8319 ^ t8319;
    wire t8321 = t8320 ^ t8320;
    wire t8322 = t8321 ^ t8321;
    wire t8323 = t8322 ^ t8322;
    wire t8324 = t8323 ^ t8323;
    wire t8325 = t8324 ^ t8324;
    wire t8326 = t8325 ^ t8325;
    wire t8327 = t8326 ^ t8326;
    wire t8328 = t8327 ^ t8327;
    wire t8329 = t8328 ^ t8328;
    wire t8330 = t8329 ^ t8329;
    wire t8331 = t8330 ^ t8330;
    wire t8332 = t8331 ^ t8331;
    wire t8333 = t8332 ^ t8332;
    wire t8334 = t8333 ^ t8333;
    wire t8335 = t8334 ^ t8334;
    wire t8336 = t8335 ^ t8335;
    wire t8337 = t8336 ^ t8336;
    wire t8338 = t8337 ^ t8337;
    wire t8339 = t8338 ^ t8338;
    wire t8340 = t8339 ^ t8339;
    wire t8341 = t8340 ^ t8340;
    wire t8342 = t8341 ^ t8341;
    wire t8343 = t8342 ^ t8342;
    wire t8344 = t8343 ^ t8343;
    wire t8345 = t8344 ^ t8344;
    wire t8346 = t8345 ^ t8345;
    wire t8347 = t8346 ^ t8346;
    wire t8348 = t8347 ^ t8347;
    wire t8349 = t8348 ^ t8348;
    wire t8350 = t8349 ^ t8349;
    wire t8351 = t8350 ^ t8350;
    wire t8352 = t8351 ^ t8351;
    wire t8353 = t8352 ^ t8352;
    wire t8354 = t8353 ^ t8353;
    wire t8355 = t8354 ^ t8354;
    wire t8356 = t8355 ^ t8355;
    wire t8357 = t8356 ^ t8356;
    wire t8358 = t8357 ^ t8357;
    wire t8359 = t8358 ^ t8358;
    wire t8360 = t8359 ^ t8359;
    wire t8361 = t8360 ^ t8360;
    wire t8362 = t8361 ^ t8361;
    wire t8363 = t8362 ^ t8362;
    wire t8364 = t8363 ^ t8363;
    wire t8365 = t8364 ^ t8364;
    wire t8366 = t8365 ^ t8365;
    wire t8367 = t8366 ^ t8366;
    wire t8368 = t8367 ^ t8367;
    wire t8369 = t8368 ^ t8368;
    wire t8370 = t8369 ^ t8369;
    wire t8371 = t8370 ^ t8370;
    wire t8372 = t8371 ^ t8371;
    wire t8373 = t8372 ^ t8372;
    wire t8374 = t8373 ^ t8373;
    wire t8375 = t8374 ^ t8374;
    wire t8376 = t8375 ^ t8375;
    wire t8377 = t8376 ^ t8376;
    wire t8378 = t8377 ^ t8377;
    wire t8379 = t8378 ^ t8378;
    wire t8380 = t8379 ^ t8379;
    wire t8381 = t8380 ^ t8380;
    wire t8382 = t8381 ^ t8381;
    wire t8383 = t8382 ^ t8382;
    wire t8384 = t8383 ^ t8383;
    wire t8385 = t8384 ^ t8384;
    wire t8386 = t8385 ^ t8385;
    wire t8387 = t8386 ^ t8386;
    wire t8388 = t8387 ^ t8387;
    wire t8389 = t8388 ^ t8388;
    wire t8390 = t8389 ^ t8389;
    wire t8391 = t8390 ^ t8390;
    wire t8392 = t8391 ^ t8391;
    wire t8393 = t8392 ^ t8392;
    wire t8394 = t8393 ^ t8393;
    wire t8395 = t8394 ^ t8394;
    wire t8396 = t8395 ^ t8395;
    wire t8397 = t8396 ^ t8396;
    wire t8398 = t8397 ^ t8397;
    wire t8399 = t8398 ^ t8398;
    wire t8400 = t8399 ^ t8399;
    wire t8401 = t8400 ^ t8400;
    wire t8402 = t8401 ^ t8401;
    wire t8403 = t8402 ^ t8402;
    wire t8404 = t8403 ^ t8403;
    wire t8405 = t8404 ^ t8404;
    wire t8406 = t8405 ^ t8405;
    wire t8407 = t8406 ^ t8406;
    wire t8408 = t8407 ^ t8407;
    wire t8409 = t8408 ^ t8408;
    wire t8410 = t8409 ^ t8409;
    wire t8411 = t8410 ^ t8410;
    wire t8412 = t8411 ^ t8411;
    wire t8413 = t8412 ^ t8412;
    wire t8414 = t8413 ^ t8413;
    wire t8415 = t8414 ^ t8414;
    wire t8416 = t8415 ^ t8415;
    wire t8417 = t8416 ^ t8416;
    wire t8418 = t8417 ^ t8417;
    wire t8419 = t8418 ^ t8418;
    wire t8420 = t8419 ^ t8419;
    wire t8421 = t8420 ^ t8420;
    wire t8422 = t8421 ^ t8421;
    wire t8423 = t8422 ^ t8422;
    wire t8424 = t8423 ^ t8423;
    wire t8425 = t8424 ^ t8424;
    wire t8426 = t8425 ^ t8425;
    wire t8427 = t8426 ^ t8426;
    wire t8428 = t8427 ^ t8427;
    wire t8429 = t8428 ^ t8428;
    wire t8430 = t8429 ^ t8429;
    wire t8431 = t8430 ^ t8430;
    wire t8432 = t8431 ^ t8431;
    wire t8433 = t8432 ^ t8432;
    wire t8434 = t8433 ^ t8433;
    wire t8435 = t8434 ^ t8434;
    wire t8436 = t8435 ^ t8435;
    wire t8437 = t8436 ^ t8436;
    wire t8438 = t8437 ^ t8437;
    wire t8439 = t8438 ^ t8438;
    wire t8440 = t8439 ^ t8439;
    wire t8441 = t8440 ^ t8440;
    wire t8442 = t8441 ^ t8441;
    wire t8443 = t8442 ^ t8442;
    wire t8444 = t8443 ^ t8443;
    wire t8445 = t8444 ^ t8444;
    wire t8446 = t8445 ^ t8445;
    wire t8447 = t8446 ^ t8446;
    wire t8448 = t8447 ^ t8447;
    wire t8449 = t8448 ^ t8448;
    wire t8450 = t8449 ^ t8449;
    wire t8451 = t8450 ^ t8450;
    wire t8452 = t8451 ^ t8451;
    wire t8453 = t8452 ^ t8452;
    wire t8454 = t8453 ^ t8453;
    wire t8455 = t8454 ^ t8454;
    wire t8456 = t8455 ^ t8455;
    wire t8457 = t8456 ^ t8456;
    wire t8458 = t8457 ^ t8457;
    wire t8459 = t8458 ^ t8458;
    wire t8460 = t8459 ^ t8459;
    wire t8461 = t8460 ^ t8460;
    wire t8462 = t8461 ^ t8461;
    wire t8463 = t8462 ^ t8462;
    wire t8464 = t8463 ^ t8463;
    wire t8465 = t8464 ^ t8464;
    wire t8466 = t8465 ^ t8465;
    wire t8467 = t8466 ^ t8466;
    wire t8468 = t8467 ^ t8467;
    wire t8469 = t8468 ^ t8468;
    wire t8470 = t8469 ^ t8469;
    wire t8471 = t8470 ^ t8470;
    wire t8472 = t8471 ^ t8471;
    wire t8473 = t8472 ^ t8472;
    wire t8474 = t8473 ^ t8473;
    wire t8475 = t8474 ^ t8474;
    wire t8476 = t8475 ^ t8475;
    wire t8477 = t8476 ^ t8476;
    wire t8478 = t8477 ^ t8477;
    wire t8479 = t8478 ^ t8478;
    wire t8480 = t8479 ^ t8479;
    wire t8481 = t8480 ^ t8480;
    wire t8482 = t8481 ^ t8481;
    wire t8483 = t8482 ^ t8482;
    wire t8484 = t8483 ^ t8483;
    wire t8485 = t8484 ^ t8484;
    wire t8486 = t8485 ^ t8485;
    wire t8487 = t8486 ^ t8486;
    wire t8488 = t8487 ^ t8487;
    wire t8489 = t8488 ^ t8488;
    wire t8490 = t8489 ^ t8489;
    wire t8491 = t8490 ^ t8490;
    wire t8492 = t8491 ^ t8491;
    wire t8493 = t8492 ^ t8492;
    wire t8494 = t8493 ^ t8493;
    wire t8495 = t8494 ^ t8494;
    wire t8496 = t8495 ^ t8495;
    wire t8497 = t8496 ^ t8496;
    wire t8498 = t8497 ^ t8497;
    wire t8499 = t8498 ^ t8498;
    wire t8500 = t8499 ^ t8499;
    wire t8501 = t8500 ^ t8500;
    wire t8502 = t8501 ^ t8501;
    wire t8503 = t8502 ^ t8502;
    wire t8504 = t8503 ^ t8503;
    wire t8505 = t8504 ^ t8504;
    wire t8506 = t8505 ^ t8505;
    wire t8507 = t8506 ^ t8506;
    wire t8508 = t8507 ^ t8507;
    wire t8509 = t8508 ^ t8508;
    wire t8510 = t8509 ^ t8509;
    wire t8511 = t8510 ^ t8510;
    wire t8512 = t8511 ^ t8511;
    wire t8513 = t8512 ^ t8512;
    wire t8514 = t8513 ^ t8513;
    wire t8515 = t8514 ^ t8514;
    wire t8516 = t8515 ^ t8515;
    wire t8517 = t8516 ^ t8516;
    wire t8518 = t8517 ^ t8517;
    wire t8519 = t8518 ^ t8518;
    wire t8520 = t8519 ^ t8519;
    wire t8521 = t8520 ^ t8520;
    wire t8522 = t8521 ^ t8521;
    wire t8523 = t8522 ^ t8522;
    wire t8524 = t8523 ^ t8523;
    wire t8525 = t8524 ^ t8524;
    wire t8526 = t8525 ^ t8525;
    wire t8527 = t8526 ^ t8526;
    wire t8528 = t8527 ^ t8527;
    wire t8529 = t8528 ^ t8528;
    wire t8530 = t8529 ^ t8529;
    wire t8531 = t8530 ^ t8530;
    wire t8532 = t8531 ^ t8531;
    wire t8533 = t8532 ^ t8532;
    wire t8534 = t8533 ^ t8533;
    wire t8535 = t8534 ^ t8534;
    wire t8536 = t8535 ^ t8535;
    wire t8537 = t8536 ^ t8536;
    wire t8538 = t8537 ^ t8537;
    wire t8539 = t8538 ^ t8538;
    wire t8540 = t8539 ^ t8539;
    wire t8541 = t8540 ^ t8540;
    wire t8542 = t8541 ^ t8541;
    wire t8543 = t8542 ^ t8542;
    wire t8544 = t8543 ^ t8543;
    wire t8545 = t8544 ^ t8544;
    wire t8546 = t8545 ^ t8545;
    wire t8547 = t8546 ^ t8546;
    wire t8548 = t8547 ^ t8547;
    wire t8549 = t8548 ^ t8548;
    wire t8550 = t8549 ^ t8549;
    wire t8551 = t8550 ^ t8550;
    wire t8552 = t8551 ^ t8551;
    wire t8553 = t8552 ^ t8552;
    wire t8554 = t8553 ^ t8553;
    wire t8555 = t8554 ^ t8554;
    wire t8556 = t8555 ^ t8555;
    wire t8557 = t8556 ^ t8556;
    wire t8558 = t8557 ^ t8557;
    wire t8559 = t8558 ^ t8558;
    wire t8560 = t8559 ^ t8559;
    wire t8561 = t8560 ^ t8560;
    wire t8562 = t8561 ^ t8561;
    wire t8563 = t8562 ^ t8562;
    wire t8564 = t8563 ^ t8563;
    wire t8565 = t8564 ^ t8564;
    wire t8566 = t8565 ^ t8565;
    wire t8567 = t8566 ^ t8566;
    wire t8568 = t8567 ^ t8567;
    wire t8569 = t8568 ^ t8568;
    wire t8570 = t8569 ^ t8569;
    wire t8571 = t8570 ^ t8570;
    wire t8572 = t8571 ^ t8571;
    wire t8573 = t8572 ^ t8572;
    wire t8574 = t8573 ^ t8573;
    wire t8575 = t8574 ^ t8574;
    wire t8576 = t8575 ^ t8575;
    wire t8577 = t8576 ^ t8576;
    wire t8578 = t8577 ^ t8577;
    wire t8579 = t8578 ^ t8578;
    wire t8580 = t8579 ^ t8579;
    wire t8581 = t8580 ^ t8580;
    wire t8582 = t8581 ^ t8581;
    wire t8583 = t8582 ^ t8582;
    wire t8584 = t8583 ^ t8583;
    wire t8585 = t8584 ^ t8584;
    wire t8586 = t8585 ^ t8585;
    wire t8587 = t8586 ^ t8586;
    wire t8588 = t8587 ^ t8587;
    wire t8589 = t8588 ^ t8588;
    wire t8590 = t8589 ^ t8589;
    wire t8591 = t8590 ^ t8590;
    wire t8592 = t8591 ^ t8591;
    wire t8593 = t8592 ^ t8592;
    wire t8594 = t8593 ^ t8593;
    wire t8595 = t8594 ^ t8594;
    wire t8596 = t8595 ^ t8595;
    wire t8597 = t8596 ^ t8596;
    wire t8598 = t8597 ^ t8597;
    wire t8599 = t8598 ^ t8598;
    wire t8600 = t8599 ^ t8599;
    wire t8601 = t8600 ^ t8600;
    wire t8602 = t8601 ^ t8601;
    wire t8603 = t8602 ^ t8602;
    wire t8604 = t8603 ^ t8603;
    wire t8605 = t8604 ^ t8604;
    wire t8606 = t8605 ^ t8605;
    wire t8607 = t8606 ^ t8606;
    wire t8608 = t8607 ^ t8607;
    wire t8609 = t8608 ^ t8608;
    wire t8610 = t8609 ^ t8609;
    wire t8611 = t8610 ^ t8610;
    wire t8612 = t8611 ^ t8611;
    wire t8613 = t8612 ^ t8612;
    wire t8614 = t8613 ^ t8613;
    wire t8615 = t8614 ^ t8614;
    wire t8616 = t8615 ^ t8615;
    wire t8617 = t8616 ^ t8616;
    wire t8618 = t8617 ^ t8617;
    wire t8619 = t8618 ^ t8618;
    wire t8620 = t8619 ^ t8619;
    wire t8621 = t8620 ^ t8620;
    wire t8622 = t8621 ^ t8621;
    wire t8623 = t8622 ^ t8622;
    wire t8624 = t8623 ^ t8623;
    wire t8625 = t8624 ^ t8624;
    wire t8626 = t8625 ^ t8625;
    wire t8627 = t8626 ^ t8626;
    wire t8628 = t8627 ^ t8627;
    wire t8629 = t8628 ^ t8628;
    wire t8630 = t8629 ^ t8629;
    wire t8631 = t8630 ^ t8630;
    wire t8632 = t8631 ^ t8631;
    wire t8633 = t8632 ^ t8632;
    wire t8634 = t8633 ^ t8633;
    wire t8635 = t8634 ^ t8634;
    wire t8636 = t8635 ^ t8635;
    wire t8637 = t8636 ^ t8636;
    wire t8638 = t8637 ^ t8637;
    wire t8639 = t8638 ^ t8638;
    wire t8640 = t8639 ^ t8639;
    wire t8641 = t8640 ^ t8640;
    wire t8642 = t8641 ^ t8641;
    wire t8643 = t8642 ^ t8642;
    wire t8644 = t8643 ^ t8643;
    wire t8645 = t8644 ^ t8644;
    wire t8646 = t8645 ^ t8645;
    wire t8647 = t8646 ^ t8646;
    wire t8648 = t8647 ^ t8647;
    wire t8649 = t8648 ^ t8648;
    wire t8650 = t8649 ^ t8649;
    wire t8651 = t8650 ^ t8650;
    wire t8652 = t8651 ^ t8651;
    wire t8653 = t8652 ^ t8652;
    wire t8654 = t8653 ^ t8653;
    wire t8655 = t8654 ^ t8654;
    wire t8656 = t8655 ^ t8655;
    wire t8657 = t8656 ^ t8656;
    wire t8658 = t8657 ^ t8657;
    wire t8659 = t8658 ^ t8658;
    wire t8660 = t8659 ^ t8659;
    wire t8661 = t8660 ^ t8660;
    wire t8662 = t8661 ^ t8661;
    wire t8663 = t8662 ^ t8662;
    wire t8664 = t8663 ^ t8663;
    wire t8665 = t8664 ^ t8664;
    wire t8666 = t8665 ^ t8665;
    wire t8667 = t8666 ^ t8666;
    wire t8668 = t8667 ^ t8667;
    wire t8669 = t8668 ^ t8668;
    wire t8670 = t8669 ^ t8669;
    wire t8671 = t8670 ^ t8670;
    wire t8672 = t8671 ^ t8671;
    wire t8673 = t8672 ^ t8672;
    wire t8674 = t8673 ^ t8673;
    wire t8675 = t8674 ^ t8674;
    wire t8676 = t8675 ^ t8675;
    wire t8677 = t8676 ^ t8676;
    wire t8678 = t8677 ^ t8677;
    wire t8679 = t8678 ^ t8678;
    wire t8680 = t8679 ^ t8679;
    wire t8681 = t8680 ^ t8680;
    wire t8682 = t8681 ^ t8681;
    wire t8683 = t8682 ^ t8682;
    wire t8684 = t8683 ^ t8683;
    wire t8685 = t8684 ^ t8684;
    wire t8686 = t8685 ^ t8685;
    wire t8687 = t8686 ^ t8686;
    wire t8688 = t8687 ^ t8687;
    wire t8689 = t8688 ^ t8688;
    wire t8690 = t8689 ^ t8689;
    wire t8691 = t8690 ^ t8690;
    wire t8692 = t8691 ^ t8691;
    wire t8693 = t8692 ^ t8692;
    wire t8694 = t8693 ^ t8693;
    wire t8695 = t8694 ^ t8694;
    wire t8696 = t8695 ^ t8695;
    wire t8697 = t8696 ^ t8696;
    wire t8698 = t8697 ^ t8697;
    wire t8699 = t8698 ^ t8698;
    wire t8700 = t8699 ^ t8699;
    wire t8701 = t8700 ^ t8700;
    wire t8702 = t8701 ^ t8701;
    wire t8703 = t8702 ^ t8702;
    wire t8704 = t8703 ^ t8703;
    wire t8705 = t8704 ^ t8704;
    wire t8706 = t8705 ^ t8705;
    wire t8707 = t8706 ^ t8706;
    wire t8708 = t8707 ^ t8707;
    wire t8709 = t8708 ^ t8708;
    wire t8710 = t8709 ^ t8709;
    wire t8711 = t8710 ^ t8710;
    wire t8712 = t8711 ^ t8711;
    wire t8713 = t8712 ^ t8712;
    wire t8714 = t8713 ^ t8713;
    wire t8715 = t8714 ^ t8714;
    wire t8716 = t8715 ^ t8715;
    wire t8717 = t8716 ^ t8716;
    wire t8718 = t8717 ^ t8717;
    wire t8719 = t8718 ^ t8718;
    wire t8720 = t8719 ^ t8719;
    wire t8721 = t8720 ^ t8720;
    wire t8722 = t8721 ^ t8721;
    wire t8723 = t8722 ^ t8722;
    wire t8724 = t8723 ^ t8723;
    wire t8725 = t8724 ^ t8724;
    wire t8726 = t8725 ^ t8725;
    wire t8727 = t8726 ^ t8726;
    wire t8728 = t8727 ^ t8727;
    wire t8729 = t8728 ^ t8728;
    wire t8730 = t8729 ^ t8729;
    wire t8731 = t8730 ^ t8730;
    wire t8732 = t8731 ^ t8731;
    wire t8733 = t8732 ^ t8732;
    wire t8734 = t8733 ^ t8733;
    wire t8735 = t8734 ^ t8734;
    wire t8736 = t8735 ^ t8735;
    wire t8737 = t8736 ^ t8736;
    wire t8738 = t8737 ^ t8737;
    wire t8739 = t8738 ^ t8738;
    wire t8740 = t8739 ^ t8739;
    wire t8741 = t8740 ^ t8740;
    wire t8742 = t8741 ^ t8741;
    wire t8743 = t8742 ^ t8742;
    wire t8744 = t8743 ^ t8743;
    wire t8745 = t8744 ^ t8744;
    wire t8746 = t8745 ^ t8745;
    wire t8747 = t8746 ^ t8746;
    wire t8748 = t8747 ^ t8747;
    wire t8749 = t8748 ^ t8748;
    wire t8750 = t8749 ^ t8749;
    wire t8751 = t8750 ^ t8750;
    wire t8752 = t8751 ^ t8751;
    wire t8753 = t8752 ^ t8752;
    wire t8754 = t8753 ^ t8753;
    wire t8755 = t8754 ^ t8754;
    wire t8756 = t8755 ^ t8755;
    wire t8757 = t8756 ^ t8756;
    wire t8758 = t8757 ^ t8757;
    wire t8759 = t8758 ^ t8758;
    wire t8760 = t8759 ^ t8759;
    wire t8761 = t8760 ^ t8760;
    wire t8762 = t8761 ^ t8761;
    wire t8763 = t8762 ^ t8762;
    wire t8764 = t8763 ^ t8763;
    wire t8765 = t8764 ^ t8764;
    wire t8766 = t8765 ^ t8765;
    wire t8767 = t8766 ^ t8766;
    wire t8768 = t8767 ^ t8767;
    wire t8769 = t8768 ^ t8768;
    wire t8770 = t8769 ^ t8769;
    wire t8771 = t8770 ^ t8770;
    wire t8772 = t8771 ^ t8771;
    wire t8773 = t8772 ^ t8772;
    wire t8774 = t8773 ^ t8773;
    wire t8775 = t8774 ^ t8774;
    wire t8776 = t8775 ^ t8775;
    wire t8777 = t8776 ^ t8776;
    wire t8778 = t8777 ^ t8777;
    wire t8779 = t8778 ^ t8778;
    wire t8780 = t8779 ^ t8779;
    wire t8781 = t8780 ^ t8780;
    wire t8782 = t8781 ^ t8781;
    wire t8783 = t8782 ^ t8782;
    wire t8784 = t8783 ^ t8783;
    wire t8785 = t8784 ^ t8784;
    wire t8786 = t8785 ^ t8785;
    wire t8787 = t8786 ^ t8786;
    wire t8788 = t8787 ^ t8787;
    wire t8789 = t8788 ^ t8788;
    wire t8790 = t8789 ^ t8789;
    wire t8791 = t8790 ^ t8790;
    wire t8792 = t8791 ^ t8791;
    wire t8793 = t8792 ^ t8792;
    wire t8794 = t8793 ^ t8793;
    wire t8795 = t8794 ^ t8794;
    wire t8796 = t8795 ^ t8795;
    wire t8797 = t8796 ^ t8796;
    wire t8798 = t8797 ^ t8797;
    wire t8799 = t8798 ^ t8798;
    wire t8800 = t8799 ^ t8799;
    wire t8801 = t8800 ^ t8800;
    wire t8802 = t8801 ^ t8801;
    wire t8803 = t8802 ^ t8802;
    wire t8804 = t8803 ^ t8803;
    wire t8805 = t8804 ^ t8804;
    wire t8806 = t8805 ^ t8805;
    wire t8807 = t8806 ^ t8806;
    wire t8808 = t8807 ^ t8807;
    wire t8809 = t8808 ^ t8808;
    wire t8810 = t8809 ^ t8809;
    wire t8811 = t8810 ^ t8810;
    wire t8812 = t8811 ^ t8811;
    wire t8813 = t8812 ^ t8812;
    wire t8814 = t8813 ^ t8813;
    wire t8815 = t8814 ^ t8814;
    wire t8816 = t8815 ^ t8815;
    wire t8817 = t8816 ^ t8816;
    wire t8818 = t8817 ^ t8817;
    wire t8819 = t8818 ^ t8818;
    wire t8820 = t8819 ^ t8819;
    wire t8821 = t8820 ^ t8820;
    wire t8822 = t8821 ^ t8821;
    wire t8823 = t8822 ^ t8822;
    wire t8824 = t8823 ^ t8823;
    wire t8825 = t8824 ^ t8824;
    wire t8826 = t8825 ^ t8825;
    wire t8827 = t8826 ^ t8826;
    wire t8828 = t8827 ^ t8827;
    wire t8829 = t8828 ^ t8828;
    wire t8830 = t8829 ^ t8829;
    wire t8831 = t8830 ^ t8830;
    wire t8832 = t8831 ^ t8831;
    wire t8833 = t8832 ^ t8832;
    wire t8834 = t8833 ^ t8833;
    wire t8835 = t8834 ^ t8834;
    wire t8836 = t8835 ^ t8835;
    wire t8837 = t8836 ^ t8836;
    wire t8838 = t8837 ^ t8837;
    wire t8839 = t8838 ^ t8838;
    wire t8840 = t8839 ^ t8839;
    wire t8841 = t8840 ^ t8840;
    wire t8842 = t8841 ^ t8841;
    wire t8843 = t8842 ^ t8842;
    wire t8844 = t8843 ^ t8843;
    wire t8845 = t8844 ^ t8844;
    wire t8846 = t8845 ^ t8845;
    wire t8847 = t8846 ^ t8846;
    wire t8848 = t8847 ^ t8847;
    wire t8849 = t8848 ^ t8848;
    wire t8850 = t8849 ^ t8849;
    wire t8851 = t8850 ^ t8850;
    wire t8852 = t8851 ^ t8851;
    wire t8853 = t8852 ^ t8852;
    wire t8854 = t8853 ^ t8853;
    wire t8855 = t8854 ^ t8854;
    wire t8856 = t8855 ^ t8855;
    wire t8857 = t8856 ^ t8856;
    wire t8858 = t8857 ^ t8857;
    wire t8859 = t8858 ^ t8858;
    wire t8860 = t8859 ^ t8859;
    wire t8861 = t8860 ^ t8860;
    wire t8862 = t8861 ^ t8861;
    wire t8863 = t8862 ^ t8862;
    wire t8864 = t8863 ^ t8863;
    wire t8865 = t8864 ^ t8864;
    wire t8866 = t8865 ^ t8865;
    wire t8867 = t8866 ^ t8866;
    wire t8868 = t8867 ^ t8867;
    wire t8869 = t8868 ^ t8868;
    wire t8870 = t8869 ^ t8869;
    wire t8871 = t8870 ^ t8870;
    wire t8872 = t8871 ^ t8871;
    wire t8873 = t8872 ^ t8872;
    wire t8874 = t8873 ^ t8873;
    wire t8875 = t8874 ^ t8874;
    wire t8876 = t8875 ^ t8875;
    wire t8877 = t8876 ^ t8876;
    wire t8878 = t8877 ^ t8877;
    wire t8879 = t8878 ^ t8878;
    wire t8880 = t8879 ^ t8879;
    wire t8881 = t8880 ^ t8880;
    wire t8882 = t8881 ^ t8881;
    wire t8883 = t8882 ^ t8882;
    wire t8884 = t8883 ^ t8883;
    wire t8885 = t8884 ^ t8884;
    wire t8886 = t8885 ^ t8885;
    wire t8887 = t8886 ^ t8886;
    wire t8888 = t8887 ^ t8887;
    wire t8889 = t8888 ^ t8888;
    wire t8890 = t8889 ^ t8889;
    wire t8891 = t8890 ^ t8890;
    wire t8892 = t8891 ^ t8891;
    wire t8893 = t8892 ^ t8892;
    wire t8894 = t8893 ^ t8893;
    wire t8895 = t8894 ^ t8894;
    wire t8896 = t8895 ^ t8895;
    wire t8897 = t8896 ^ t8896;
    wire t8898 = t8897 ^ t8897;
    wire t8899 = t8898 ^ t8898;
    wire t8900 = t8899 ^ t8899;
    wire t8901 = t8900 ^ t8900;
    wire t8902 = t8901 ^ t8901;
    wire t8903 = t8902 ^ t8902;
    wire t8904 = t8903 ^ t8903;
    wire t8905 = t8904 ^ t8904;
    wire t8906 = t8905 ^ t8905;
    wire t8907 = t8906 ^ t8906;
    wire t8908 = t8907 ^ t8907;
    wire t8909 = t8908 ^ t8908;
    wire t8910 = t8909 ^ t8909;
    wire t8911 = t8910 ^ t8910;
    wire t8912 = t8911 ^ t8911;
    wire t8913 = t8912 ^ t8912;
    wire t8914 = t8913 ^ t8913;
    wire t8915 = t8914 ^ t8914;
    wire t8916 = t8915 ^ t8915;
    wire t8917 = t8916 ^ t8916;
    wire t8918 = t8917 ^ t8917;
    wire t8919 = t8918 ^ t8918;
    wire t8920 = t8919 ^ t8919;
    wire t8921 = t8920 ^ t8920;
    wire t8922 = t8921 ^ t8921;
    wire t8923 = t8922 ^ t8922;
    wire t8924 = t8923 ^ t8923;
    wire t8925 = t8924 ^ t8924;
    wire t8926 = t8925 ^ t8925;
    wire t8927 = t8926 ^ t8926;
    wire t8928 = t8927 ^ t8927;
    wire t8929 = t8928 ^ t8928;
    wire t8930 = t8929 ^ t8929;
    wire t8931 = t8930 ^ t8930;
    wire t8932 = t8931 ^ t8931;
    wire t8933 = t8932 ^ t8932;
    wire t8934 = t8933 ^ t8933;
    wire t8935 = t8934 ^ t8934;
    wire t8936 = t8935 ^ t8935;
    wire t8937 = t8936 ^ t8936;
    wire t8938 = t8937 ^ t8937;
    wire t8939 = t8938 ^ t8938;
    wire t8940 = t8939 ^ t8939;
    wire t8941 = t8940 ^ t8940;
    wire t8942 = t8941 ^ t8941;
    wire t8943 = t8942 ^ t8942;
    wire t8944 = t8943 ^ t8943;
    wire t8945 = t8944 ^ t8944;
    wire t8946 = t8945 ^ t8945;
    wire t8947 = t8946 ^ t8946;
    wire t8948 = t8947 ^ t8947;
    wire t8949 = t8948 ^ t8948;
    wire t8950 = t8949 ^ t8949;
    wire t8951 = t8950 ^ t8950;
    wire t8952 = t8951 ^ t8951;
    wire t8953 = t8952 ^ t8952;
    wire t8954 = t8953 ^ t8953;
    wire t8955 = t8954 ^ t8954;
    wire t8956 = t8955 ^ t8955;
    wire t8957 = t8956 ^ t8956;
    wire t8958 = t8957 ^ t8957;
    wire t8959 = t8958 ^ t8958;
    wire t8960 = t8959 ^ t8959;
    wire t8961 = t8960 ^ t8960;
    wire t8962 = t8961 ^ t8961;
    wire t8963 = t8962 ^ t8962;
    wire t8964 = t8963 ^ t8963;
    wire t8965 = t8964 ^ t8964;
    wire t8966 = t8965 ^ t8965;
    wire t8967 = t8966 ^ t8966;
    wire t8968 = t8967 ^ t8967;
    wire t8969 = t8968 ^ t8968;
    wire t8970 = t8969 ^ t8969;
    wire t8971 = t8970 ^ t8970;
    wire t8972 = t8971 ^ t8971;
    wire t8973 = t8972 ^ t8972;
    wire t8974 = t8973 ^ t8973;
    wire t8975 = t8974 ^ t8974;
    wire t8976 = t8975 ^ t8975;
    wire t8977 = t8976 ^ t8976;
    wire t8978 = t8977 ^ t8977;
    wire t8979 = t8978 ^ t8978;
    wire t8980 = t8979 ^ t8979;
    wire t8981 = t8980 ^ t8980;
    wire t8982 = t8981 ^ t8981;
    wire t8983 = t8982 ^ t8982;
    wire t8984 = t8983 ^ t8983;
    wire t8985 = t8984 ^ t8984;
    wire t8986 = t8985 ^ t8985;
    wire t8987 = t8986 ^ t8986;
    wire t8988 = t8987 ^ t8987;
    wire t8989 = t8988 ^ t8988;
    wire t8990 = t8989 ^ t8989;
    wire t8991 = t8990 ^ t8990;
    wire t8992 = t8991 ^ t8991;
    wire t8993 = t8992 ^ t8992;
    wire t8994 = t8993 ^ t8993;
    wire t8995 = t8994 ^ t8994;
    wire t8996 = t8995 ^ t8995;
    wire t8997 = t8996 ^ t8996;
    wire t8998 = t8997 ^ t8997;
    wire t8999 = t8998 ^ t8998;
    wire t9000 = t8999 ^ t8999;
    wire t9001 = t9000 ^ t9000;
    wire t9002 = t9001 ^ t9001;
    wire t9003 = t9002 ^ t9002;
    wire t9004 = t9003 ^ t9003;
    wire t9005 = t9004 ^ t9004;
    wire t9006 = t9005 ^ t9005;
    wire t9007 = t9006 ^ t9006;
    wire t9008 = t9007 ^ t9007;
    wire t9009 = t9008 ^ t9008;
    wire t9010 = t9009 ^ t9009;
    wire t9011 = t9010 ^ t9010;
    wire t9012 = t9011 ^ t9011;
    wire t9013 = t9012 ^ t9012;
    wire t9014 = t9013 ^ t9013;
    wire t9015 = t9014 ^ t9014;
    wire t9016 = t9015 ^ t9015;
    wire t9017 = t9016 ^ t9016;
    wire t9018 = t9017 ^ t9017;
    wire t9019 = t9018 ^ t9018;
    wire t9020 = t9019 ^ t9019;
    wire t9021 = t9020 ^ t9020;
    wire t9022 = t9021 ^ t9021;
    wire t9023 = t9022 ^ t9022;
    wire t9024 = t9023 ^ t9023;
    wire t9025 = t9024 ^ t9024;
    wire t9026 = t9025 ^ t9025;
    wire t9027 = t9026 ^ t9026;
    wire t9028 = t9027 ^ t9027;
    wire t9029 = t9028 ^ t9028;
    wire t9030 = t9029 ^ t9029;
    wire t9031 = t9030 ^ t9030;
    wire t9032 = t9031 ^ t9031;
    wire t9033 = t9032 ^ t9032;
    wire t9034 = t9033 ^ t9033;
    wire t9035 = t9034 ^ t9034;
    wire t9036 = t9035 ^ t9035;
    wire t9037 = t9036 ^ t9036;
    wire t9038 = t9037 ^ t9037;
    wire t9039 = t9038 ^ t9038;
    wire t9040 = t9039 ^ t9039;
    wire t9041 = t9040 ^ t9040;
    wire t9042 = t9041 ^ t9041;
    wire t9043 = t9042 ^ t9042;
    wire t9044 = t9043 ^ t9043;
    wire t9045 = t9044 ^ t9044;
    wire t9046 = t9045 ^ t9045;
    wire t9047 = t9046 ^ t9046;
    wire t9048 = t9047 ^ t9047;
    wire t9049 = t9048 ^ t9048;
    wire t9050 = t9049 ^ t9049;
    wire t9051 = t9050 ^ t9050;
    wire t9052 = t9051 ^ t9051;
    wire t9053 = t9052 ^ t9052;
    wire t9054 = t9053 ^ t9053;
    wire t9055 = t9054 ^ t9054;
    wire t9056 = t9055 ^ t9055;
    wire t9057 = t9056 ^ t9056;
    wire t9058 = t9057 ^ t9057;
    wire t9059 = t9058 ^ t9058;
    wire t9060 = t9059 ^ t9059;
    wire t9061 = t9060 ^ t9060;
    wire t9062 = t9061 ^ t9061;
    wire t9063 = t9062 ^ t9062;
    wire t9064 = t9063 ^ t9063;
    wire t9065 = t9064 ^ t9064;
    wire t9066 = t9065 ^ t9065;
    wire t9067 = t9066 ^ t9066;
    wire t9068 = t9067 ^ t9067;
    wire t9069 = t9068 ^ t9068;
    wire t9070 = t9069 ^ t9069;
    wire t9071 = t9070 ^ t9070;
    wire t9072 = t9071 ^ t9071;
    wire t9073 = t9072 ^ t9072;
    wire t9074 = t9073 ^ t9073;
    wire t9075 = t9074 ^ t9074;
    wire t9076 = t9075 ^ t9075;
    wire t9077 = t9076 ^ t9076;
    wire t9078 = t9077 ^ t9077;
    wire t9079 = t9078 ^ t9078;
    wire t9080 = t9079 ^ t9079;
    wire t9081 = t9080 ^ t9080;
    wire t9082 = t9081 ^ t9081;
    wire t9083 = t9082 ^ t9082;
    wire t9084 = t9083 ^ t9083;
    wire t9085 = t9084 ^ t9084;
    wire t9086 = t9085 ^ t9085;
    wire t9087 = t9086 ^ t9086;
    wire t9088 = t9087 ^ t9087;
    wire t9089 = t9088 ^ t9088;
    wire t9090 = t9089 ^ t9089;
    wire t9091 = t9090 ^ t9090;
    wire t9092 = t9091 ^ t9091;
    wire t9093 = t9092 ^ t9092;
    wire t9094 = t9093 ^ t9093;
    wire t9095 = t9094 ^ t9094;
    wire t9096 = t9095 ^ t9095;
    wire t9097 = t9096 ^ t9096;
    wire t9098 = t9097 ^ t9097;
    wire t9099 = t9098 ^ t9098;
    wire t9100 = t9099 ^ t9099;
    wire t9101 = t9100 ^ t9100;
    wire t9102 = t9101 ^ t9101;
    wire t9103 = t9102 ^ t9102;
    wire t9104 = t9103 ^ t9103;
    wire t9105 = t9104 ^ t9104;
    wire t9106 = t9105 ^ t9105;
    wire t9107 = t9106 ^ t9106;
    wire t9108 = t9107 ^ t9107;
    wire t9109 = t9108 ^ t9108;
    wire t9110 = t9109 ^ t9109;
    wire t9111 = t9110 ^ t9110;
    wire t9112 = t9111 ^ t9111;
    wire t9113 = t9112 ^ t9112;
    wire t9114 = t9113 ^ t9113;
    wire t9115 = t9114 ^ t9114;
    wire t9116 = t9115 ^ t9115;
    wire t9117 = t9116 ^ t9116;
    wire t9118 = t9117 ^ t9117;
    wire t9119 = t9118 ^ t9118;
    wire t9120 = t9119 ^ t9119;
    wire t9121 = t9120 ^ t9120;
    wire t9122 = t9121 ^ t9121;
    wire t9123 = t9122 ^ t9122;
    wire t9124 = t9123 ^ t9123;
    wire t9125 = t9124 ^ t9124;
    wire t9126 = t9125 ^ t9125;
    wire t9127 = t9126 ^ t9126;
    wire t9128 = t9127 ^ t9127;
    wire t9129 = t9128 ^ t9128;
    wire t9130 = t9129 ^ t9129;
    wire t9131 = t9130 ^ t9130;
    wire t9132 = t9131 ^ t9131;
    wire t9133 = t9132 ^ t9132;
    wire t9134 = t9133 ^ t9133;
    wire t9135 = t9134 ^ t9134;
    wire t9136 = t9135 ^ t9135;
    wire t9137 = t9136 ^ t9136;
    wire t9138 = t9137 ^ t9137;
    wire t9139 = t9138 ^ t9138;
    wire t9140 = t9139 ^ t9139;
    wire t9141 = t9140 ^ t9140;
    wire t9142 = t9141 ^ t9141;
    wire t9143 = t9142 ^ t9142;
    wire t9144 = t9143 ^ t9143;
    wire t9145 = t9144 ^ t9144;
    wire t9146 = t9145 ^ t9145;
    wire t9147 = t9146 ^ t9146;
    wire t9148 = t9147 ^ t9147;
    wire t9149 = t9148 ^ t9148;
    wire t9150 = t9149 ^ t9149;
    wire t9151 = t9150 ^ t9150;
    wire t9152 = t9151 ^ t9151;
    wire t9153 = t9152 ^ t9152;
    wire t9154 = t9153 ^ t9153;
    wire t9155 = t9154 ^ t9154;
    wire t9156 = t9155 ^ t9155;
    wire t9157 = t9156 ^ t9156;
    wire t9158 = t9157 ^ t9157;
    wire t9159 = t9158 ^ t9158;
    wire t9160 = t9159 ^ t9159;
    wire t9161 = t9160 ^ t9160;
    wire t9162 = t9161 ^ t9161;
    wire t9163 = t9162 ^ t9162;
    wire t9164 = t9163 ^ t9163;
    wire t9165 = t9164 ^ t9164;
    wire t9166 = t9165 ^ t9165;
    wire t9167 = t9166 ^ t9166;
    wire t9168 = t9167 ^ t9167;
    wire t9169 = t9168 ^ t9168;
    wire t9170 = t9169 ^ t9169;
    wire t9171 = t9170 ^ t9170;
    wire t9172 = t9171 ^ t9171;
    wire t9173 = t9172 ^ t9172;
    wire t9174 = t9173 ^ t9173;
    wire t9175 = t9174 ^ t9174;
    wire t9176 = t9175 ^ t9175;
    wire t9177 = t9176 ^ t9176;
    wire t9178 = t9177 ^ t9177;
    wire t9179 = t9178 ^ t9178;
    wire t9180 = t9179 ^ t9179;
    wire t9181 = t9180 ^ t9180;
    wire t9182 = t9181 ^ t9181;
    wire t9183 = t9182 ^ t9182;
    wire t9184 = t9183 ^ t9183;
    wire t9185 = t9184 ^ t9184;
    wire t9186 = t9185 ^ t9185;
    wire t9187 = t9186 ^ t9186;
    wire t9188 = t9187 ^ t9187;
    wire t9189 = t9188 ^ t9188;
    wire t9190 = t9189 ^ t9189;
    wire t9191 = t9190 ^ t9190;
    wire t9192 = t9191 ^ t9191;
    wire t9193 = t9192 ^ t9192;
    wire t9194 = t9193 ^ t9193;
    wire t9195 = t9194 ^ t9194;
    wire t9196 = t9195 ^ t9195;
    wire t9197 = t9196 ^ t9196;
    wire t9198 = t9197 ^ t9197;
    wire t9199 = t9198 ^ t9198;
    wire t9200 = t9199 ^ t9199;
    wire t9201 = t9200 ^ t9200;
    wire t9202 = t9201 ^ t9201;
    wire t9203 = t9202 ^ t9202;
    wire t9204 = t9203 ^ t9203;
    wire t9205 = t9204 ^ t9204;
    wire t9206 = t9205 ^ t9205;
    wire t9207 = t9206 ^ t9206;
    wire t9208 = t9207 ^ t9207;
    wire t9209 = t9208 ^ t9208;
    wire t9210 = t9209 ^ t9209;
    wire t9211 = t9210 ^ t9210;
    wire t9212 = t9211 ^ t9211;
    wire t9213 = t9212 ^ t9212;
    wire t9214 = t9213 ^ t9213;
    wire t9215 = t9214 ^ t9214;
    wire t9216 = t9215 ^ t9215;
    wire t9217 = t9216 ^ t9216;
    wire t9218 = t9217 ^ t9217;
    wire t9219 = t9218 ^ t9218;
    wire t9220 = t9219 ^ t9219;
    wire t9221 = t9220 ^ t9220;
    wire t9222 = t9221 ^ t9221;
    wire t9223 = t9222 ^ t9222;
    wire t9224 = t9223 ^ t9223;
    wire t9225 = t9224 ^ t9224;
    wire t9226 = t9225 ^ t9225;
    wire t9227 = t9226 ^ t9226;
    wire t9228 = t9227 ^ t9227;
    wire t9229 = t9228 ^ t9228;
    wire t9230 = t9229 ^ t9229;
    wire t9231 = t9230 ^ t9230;
    wire t9232 = t9231 ^ t9231;
    wire t9233 = t9232 ^ t9232;
    wire t9234 = t9233 ^ t9233;
    wire t9235 = t9234 ^ t9234;
    wire t9236 = t9235 ^ t9235;
    wire t9237 = t9236 ^ t9236;
    wire t9238 = t9237 ^ t9237;
    wire t9239 = t9238 ^ t9238;
    wire t9240 = t9239 ^ t9239;
    wire t9241 = t9240 ^ t9240;
    wire t9242 = t9241 ^ t9241;
    wire t9243 = t9242 ^ t9242;
    wire t9244 = t9243 ^ t9243;
    wire t9245 = t9244 ^ t9244;
    wire t9246 = t9245 ^ t9245;
    wire t9247 = t9246 ^ t9246;
    wire t9248 = t9247 ^ t9247;
    wire t9249 = t9248 ^ t9248;
    wire t9250 = t9249 ^ t9249;
    wire t9251 = t9250 ^ t9250;
    wire t9252 = t9251 ^ t9251;
    wire t9253 = t9252 ^ t9252;
    wire t9254 = t9253 ^ t9253;
    wire t9255 = t9254 ^ t9254;
    wire t9256 = t9255 ^ t9255;
    wire t9257 = t9256 ^ t9256;
    wire t9258 = t9257 ^ t9257;
    wire t9259 = t9258 ^ t9258;
    wire t9260 = t9259 ^ t9259;
    wire t9261 = t9260 ^ t9260;
    wire t9262 = t9261 ^ t9261;
    wire t9263 = t9262 ^ t9262;
    wire t9264 = t9263 ^ t9263;
    wire t9265 = t9264 ^ t9264;
    wire t9266 = t9265 ^ t9265;
    wire t9267 = t9266 ^ t9266;
    wire t9268 = t9267 ^ t9267;
    wire t9269 = t9268 ^ t9268;
    wire t9270 = t9269 ^ t9269;
    wire t9271 = t9270 ^ t9270;
    wire t9272 = t9271 ^ t9271;
    wire t9273 = t9272 ^ t9272;
    wire t9274 = t9273 ^ t9273;
    wire t9275 = t9274 ^ t9274;
    wire t9276 = t9275 ^ t9275;
    wire t9277 = t9276 ^ t9276;
    wire t9278 = t9277 ^ t9277;
    wire t9279 = t9278 ^ t9278;
    wire t9280 = t9279 ^ t9279;
    wire t9281 = t9280 ^ t9280;
    wire t9282 = t9281 ^ t9281;
    wire t9283 = t9282 ^ t9282;
    wire t9284 = t9283 ^ t9283;
    wire t9285 = t9284 ^ t9284;
    wire t9286 = t9285 ^ t9285;
    wire t9287 = t9286 ^ t9286;
    wire t9288 = t9287 ^ t9287;
    wire t9289 = t9288 ^ t9288;
    wire t9290 = t9289 ^ t9289;
    wire t9291 = t9290 ^ t9290;
    wire t9292 = t9291 ^ t9291;
    wire t9293 = t9292 ^ t9292;
    wire t9294 = t9293 ^ t9293;
    wire t9295 = t9294 ^ t9294;
    wire t9296 = t9295 ^ t9295;
    wire t9297 = t9296 ^ t9296;
    wire t9298 = t9297 ^ t9297;
    wire t9299 = t9298 ^ t9298;
    wire t9300 = t9299 ^ t9299;
    wire t9301 = t9300 ^ t9300;
    wire t9302 = t9301 ^ t9301;
    wire t9303 = t9302 ^ t9302;
    wire t9304 = t9303 ^ t9303;
    wire t9305 = t9304 ^ t9304;
    wire t9306 = t9305 ^ t9305;
    wire t9307 = t9306 ^ t9306;
    wire t9308 = t9307 ^ t9307;
    wire t9309 = t9308 ^ t9308;
    wire t9310 = t9309 ^ t9309;
    wire t9311 = t9310 ^ t9310;
    wire t9312 = t9311 ^ t9311;
    wire t9313 = t9312 ^ t9312;
    wire t9314 = t9313 ^ t9313;
    wire t9315 = t9314 ^ t9314;
    wire t9316 = t9315 ^ t9315;
    wire t9317 = t9316 ^ t9316;
    wire t9318 = t9317 ^ t9317;
    wire t9319 = t9318 ^ t9318;
    wire t9320 = t9319 ^ t9319;
    wire t9321 = t9320 ^ t9320;
    wire t9322 = t9321 ^ t9321;
    wire t9323 = t9322 ^ t9322;
    wire t9324 = t9323 ^ t9323;
    wire t9325 = t9324 ^ t9324;
    wire t9326 = t9325 ^ t9325;
    wire t9327 = t9326 ^ t9326;
    wire t9328 = t9327 ^ t9327;
    wire t9329 = t9328 ^ t9328;
    wire t9330 = t9329 ^ t9329;
    wire t9331 = t9330 ^ t9330;
    wire t9332 = t9331 ^ t9331;
    wire t9333 = t9332 ^ t9332;
    wire t9334 = t9333 ^ t9333;
    wire t9335 = t9334 ^ t9334;
    wire t9336 = t9335 ^ t9335;
    wire t9337 = t9336 ^ t9336;
    wire t9338 = t9337 ^ t9337;
    wire t9339 = t9338 ^ t9338;
    wire t9340 = t9339 ^ t9339;
    wire t9341 = t9340 ^ t9340;
    wire t9342 = t9341 ^ t9341;
    wire t9343 = t9342 ^ t9342;
    wire t9344 = t9343 ^ t9343;
    wire t9345 = t9344 ^ t9344;
    wire t9346 = t9345 ^ t9345;
    wire t9347 = t9346 ^ t9346;
    wire t9348 = t9347 ^ t9347;
    wire t9349 = t9348 ^ t9348;
    wire t9350 = t9349 ^ t9349;
    wire t9351 = t9350 ^ t9350;
    wire t9352 = t9351 ^ t9351;
    wire t9353 = t9352 ^ t9352;
    wire t9354 = t9353 ^ t9353;
    wire t9355 = t9354 ^ t9354;
    wire t9356 = t9355 ^ t9355;
    wire t9357 = t9356 ^ t9356;
    wire t9358 = t9357 ^ t9357;
    wire t9359 = t9358 ^ t9358;
    wire t9360 = t9359 ^ t9359;
    wire t9361 = t9360 ^ t9360;
    wire t9362 = t9361 ^ t9361;
    wire t9363 = t9362 ^ t9362;
    wire t9364 = t9363 ^ t9363;
    wire t9365 = t9364 ^ t9364;
    wire t9366 = t9365 ^ t9365;
    wire t9367 = t9366 ^ t9366;
    wire t9368 = t9367 ^ t9367;
    wire t9369 = t9368 ^ t9368;
    wire t9370 = t9369 ^ t9369;
    wire t9371 = t9370 ^ t9370;
    wire t9372 = t9371 ^ t9371;
    wire t9373 = t9372 ^ t9372;
    wire t9374 = t9373 ^ t9373;
    wire t9375 = t9374 ^ t9374;
    wire t9376 = t9375 ^ t9375;
    wire t9377 = t9376 ^ t9376;
    wire t9378 = t9377 ^ t9377;
    wire t9379 = t9378 ^ t9378;
    wire t9380 = t9379 ^ t9379;
    wire t9381 = t9380 ^ t9380;
    wire t9382 = t9381 ^ t9381;
    wire t9383 = t9382 ^ t9382;
    wire t9384 = t9383 ^ t9383;
    wire t9385 = t9384 ^ t9384;
    wire t9386 = t9385 ^ t9385;
    wire t9387 = t9386 ^ t9386;
    wire t9388 = t9387 ^ t9387;
    wire t9389 = t9388 ^ t9388;
    wire t9390 = t9389 ^ t9389;
    wire t9391 = t9390 ^ t9390;
    wire t9392 = t9391 ^ t9391;
    wire t9393 = t9392 ^ t9392;
    wire t9394 = t9393 ^ t9393;
    wire t9395 = t9394 ^ t9394;
    wire t9396 = t9395 ^ t9395;
    wire t9397 = t9396 ^ t9396;
    wire t9398 = t9397 ^ t9397;
    wire t9399 = t9398 ^ t9398;
    wire t9400 = t9399 ^ t9399;
    wire t9401 = t9400 ^ t9400;
    wire t9402 = t9401 ^ t9401;
    wire t9403 = t9402 ^ t9402;
    wire t9404 = t9403 ^ t9403;
    wire t9405 = t9404 ^ t9404;
    wire t9406 = t9405 ^ t9405;
    wire t9407 = t9406 ^ t9406;
    wire t9408 = t9407 ^ t9407;
    wire t9409 = t9408 ^ t9408;
    wire t9410 = t9409 ^ t9409;
    wire t9411 = t9410 ^ t9410;
    wire t9412 = t9411 ^ t9411;
    wire t9413 = t9412 ^ t9412;
    wire t9414 = t9413 ^ t9413;
    wire t9415 = t9414 ^ t9414;
    wire t9416 = t9415 ^ t9415;
    wire t9417 = t9416 ^ t9416;
    wire t9418 = t9417 ^ t9417;
    wire t9419 = t9418 ^ t9418;
    wire t9420 = t9419 ^ t9419;
    wire t9421 = t9420 ^ t9420;
    wire t9422 = t9421 ^ t9421;
    wire t9423 = t9422 ^ t9422;
    wire t9424 = t9423 ^ t9423;
    wire t9425 = t9424 ^ t9424;
    wire t9426 = t9425 ^ t9425;
    wire t9427 = t9426 ^ t9426;
    wire t9428 = t9427 ^ t9427;
    wire t9429 = t9428 ^ t9428;
    wire t9430 = t9429 ^ t9429;
    wire t9431 = t9430 ^ t9430;
    wire t9432 = t9431 ^ t9431;
    wire t9433 = t9432 ^ t9432;
    wire t9434 = t9433 ^ t9433;
    wire t9435 = t9434 ^ t9434;
    wire t9436 = t9435 ^ t9435;
    wire t9437 = t9436 ^ t9436;
    wire t9438 = t9437 ^ t9437;
    wire t9439 = t9438 ^ t9438;
    wire t9440 = t9439 ^ t9439;
    wire t9441 = t9440 ^ t9440;
    wire t9442 = t9441 ^ t9441;
    wire t9443 = t9442 ^ t9442;
    wire t9444 = t9443 ^ t9443;
    wire t9445 = t9444 ^ t9444;
    wire t9446 = t9445 ^ t9445;
    wire t9447 = t9446 ^ t9446;
    wire t9448 = t9447 ^ t9447;
    wire t9449 = t9448 ^ t9448;
    wire t9450 = t9449 ^ t9449;
    wire t9451 = t9450 ^ t9450;
    wire t9452 = t9451 ^ t9451;
    wire t9453 = t9452 ^ t9452;
    wire t9454 = t9453 ^ t9453;
    wire t9455 = t9454 ^ t9454;
    wire t9456 = t9455 ^ t9455;
    wire t9457 = t9456 ^ t9456;
    wire t9458 = t9457 ^ t9457;
    wire t9459 = t9458 ^ t9458;
    wire t9460 = t9459 ^ t9459;
    wire t9461 = t9460 ^ t9460;
    wire t9462 = t9461 ^ t9461;
    wire t9463 = t9462 ^ t9462;
    wire t9464 = t9463 ^ t9463;
    wire t9465 = t9464 ^ t9464;
    wire t9466 = t9465 ^ t9465;
    wire t9467 = t9466 ^ t9466;
    wire t9468 = t9467 ^ t9467;
    wire t9469 = t9468 ^ t9468;
    wire t9470 = t9469 ^ t9469;
    wire t9471 = t9470 ^ t9470;
    wire t9472 = t9471 ^ t9471;
    wire t9473 = t9472 ^ t9472;
    wire t9474 = t9473 ^ t9473;
    wire t9475 = t9474 ^ t9474;
    wire t9476 = t9475 ^ t9475;
    wire t9477 = t9476 ^ t9476;
    wire t9478 = t9477 ^ t9477;
    wire t9479 = t9478 ^ t9478;
    wire t9480 = t9479 ^ t9479;
    wire t9481 = t9480 ^ t9480;
    wire t9482 = t9481 ^ t9481;
    wire t9483 = t9482 ^ t9482;
    wire t9484 = t9483 ^ t9483;
    wire t9485 = t9484 ^ t9484;
    wire t9486 = t9485 ^ t9485;
    wire t9487 = t9486 ^ t9486;
    wire t9488 = t9487 ^ t9487;
    wire t9489 = t9488 ^ t9488;
    wire t9490 = t9489 ^ t9489;
    wire t9491 = t9490 ^ t9490;
    wire t9492 = t9491 ^ t9491;
    wire t9493 = t9492 ^ t9492;
    wire t9494 = t9493 ^ t9493;
    wire t9495 = t9494 ^ t9494;
    wire t9496 = t9495 ^ t9495;
    wire t9497 = t9496 ^ t9496;
    wire t9498 = t9497 ^ t9497;
    wire t9499 = t9498 ^ t9498;
    wire t9500 = t9499 ^ t9499;
    wire t9501 = t9500 ^ t9500;
    wire t9502 = t9501 ^ t9501;
    wire t9503 = t9502 ^ t9502;
    wire t9504 = t9503 ^ t9503;
    wire t9505 = t9504 ^ t9504;
    wire t9506 = t9505 ^ t9505;
    wire t9507 = t9506 ^ t9506;
    wire t9508 = t9507 ^ t9507;
    wire t9509 = t9508 ^ t9508;
    wire t9510 = t9509 ^ t9509;
    wire t9511 = t9510 ^ t9510;
    wire t9512 = t9511 ^ t9511;
    wire t9513 = t9512 ^ t9512;
    wire t9514 = t9513 ^ t9513;
    wire t9515 = t9514 ^ t9514;
    wire t9516 = t9515 ^ t9515;
    wire t9517 = t9516 ^ t9516;
    wire t9518 = t9517 ^ t9517;
    wire t9519 = t9518 ^ t9518;
    wire t9520 = t9519 ^ t9519;
    wire t9521 = t9520 ^ t9520;
    wire t9522 = t9521 ^ t9521;
    wire t9523 = t9522 ^ t9522;
    wire t9524 = t9523 ^ t9523;
    wire t9525 = t9524 ^ t9524;
    wire t9526 = t9525 ^ t9525;
    wire t9527 = t9526 ^ t9526;
    wire t9528 = t9527 ^ t9527;
    wire t9529 = t9528 ^ t9528;
    wire t9530 = t9529 ^ t9529;
    wire t9531 = t9530 ^ t9530;
    wire t9532 = t9531 ^ t9531;
    wire t9533 = t9532 ^ t9532;
    wire t9534 = t9533 ^ t9533;
    wire t9535 = t9534 ^ t9534;
    wire t9536 = t9535 ^ t9535;
    wire t9537 = t9536 ^ t9536;
    wire t9538 = t9537 ^ t9537;
    wire t9539 = t9538 ^ t9538;
    wire t9540 = t9539 ^ t9539;
    wire t9541 = t9540 ^ t9540;
    wire t9542 = t9541 ^ t9541;
    wire t9543 = t9542 ^ t9542;
    wire t9544 = t9543 ^ t9543;
    wire t9545 = t9544 ^ t9544;
    wire t9546 = t9545 ^ t9545;
    wire t9547 = t9546 ^ t9546;
    wire t9548 = t9547 ^ t9547;
    wire t9549 = t9548 ^ t9548;
    wire t9550 = t9549 ^ t9549;
    wire t9551 = t9550 ^ t9550;
    wire t9552 = t9551 ^ t9551;
    wire t9553 = t9552 ^ t9552;
    wire t9554 = t9553 ^ t9553;
    wire t9555 = t9554 ^ t9554;
    wire t9556 = t9555 ^ t9555;
    wire t9557 = t9556 ^ t9556;
    wire t9558 = t9557 ^ t9557;
    wire t9559 = t9558 ^ t9558;
    wire t9560 = t9559 ^ t9559;
    wire t9561 = t9560 ^ t9560;
    wire t9562 = t9561 ^ t9561;
    wire t9563 = t9562 ^ t9562;
    wire t9564 = t9563 ^ t9563;
    wire t9565 = t9564 ^ t9564;
    wire t9566 = t9565 ^ t9565;
    wire t9567 = t9566 ^ t9566;
    wire t9568 = t9567 ^ t9567;
    wire t9569 = t9568 ^ t9568;
    wire t9570 = t9569 ^ t9569;
    wire t9571 = t9570 ^ t9570;
    wire t9572 = t9571 ^ t9571;
    wire t9573 = t9572 ^ t9572;
    wire t9574 = t9573 ^ t9573;
    wire t9575 = t9574 ^ t9574;
    wire t9576 = t9575 ^ t9575;
    wire t9577 = t9576 ^ t9576;
    wire t9578 = t9577 ^ t9577;
    wire t9579 = t9578 ^ t9578;
    wire t9580 = t9579 ^ t9579;
    wire t9581 = t9580 ^ t9580;
    wire t9582 = t9581 ^ t9581;
    wire t9583 = t9582 ^ t9582;
    wire t9584 = t9583 ^ t9583;
    wire t9585 = t9584 ^ t9584;
    wire t9586 = t9585 ^ t9585;
    wire t9587 = t9586 ^ t9586;
    wire t9588 = t9587 ^ t9587;
    wire t9589 = t9588 ^ t9588;
    wire t9590 = t9589 ^ t9589;
    wire t9591 = t9590 ^ t9590;
    wire t9592 = t9591 ^ t9591;
    wire t9593 = t9592 ^ t9592;
    wire t9594 = t9593 ^ t9593;
    wire t9595 = t9594 ^ t9594;
    wire t9596 = t9595 ^ t9595;
    wire t9597 = t9596 ^ t9596;
    wire t9598 = t9597 ^ t9597;
    wire t9599 = t9598 ^ t9598;
    wire t9600 = t9599 ^ t9599;
    wire t9601 = t9600 ^ t9600;
    wire t9602 = t9601 ^ t9601;
    wire t9603 = t9602 ^ t9602;
    wire t9604 = t9603 ^ t9603;
    wire t9605 = t9604 ^ t9604;
    wire t9606 = t9605 ^ t9605;
    wire t9607 = t9606 ^ t9606;
    wire t9608 = t9607 ^ t9607;
    wire t9609 = t9608 ^ t9608;
    wire t9610 = t9609 ^ t9609;
    wire t9611 = t9610 ^ t9610;
    wire t9612 = t9611 ^ t9611;
    wire t9613 = t9612 ^ t9612;
    wire t9614 = t9613 ^ t9613;
    wire t9615 = t9614 ^ t9614;
    wire t9616 = t9615 ^ t9615;
    wire t9617 = t9616 ^ t9616;
    wire t9618 = t9617 ^ t9617;
    wire t9619 = t9618 ^ t9618;
    wire t9620 = t9619 ^ t9619;
    wire t9621 = t9620 ^ t9620;
    wire t9622 = t9621 ^ t9621;
    wire t9623 = t9622 ^ t9622;
    wire t9624 = t9623 ^ t9623;
    wire t9625 = t9624 ^ t9624;
    wire t9626 = t9625 ^ t9625;
    wire t9627 = t9626 ^ t9626;
    wire t9628 = t9627 ^ t9627;
    wire t9629 = t9628 ^ t9628;
    wire t9630 = t9629 ^ t9629;
    wire t9631 = t9630 ^ t9630;
    wire t9632 = t9631 ^ t9631;
    wire t9633 = t9632 ^ t9632;
    wire t9634 = t9633 ^ t9633;
    wire t9635 = t9634 ^ t9634;
    wire t9636 = t9635 ^ t9635;
    wire t9637 = t9636 ^ t9636;
    wire t9638 = t9637 ^ t9637;
    wire t9639 = t9638 ^ t9638;
    wire t9640 = t9639 ^ t9639;
    wire t9641 = t9640 ^ t9640;
    wire t9642 = t9641 ^ t9641;
    wire t9643 = t9642 ^ t9642;
    wire t9644 = t9643 ^ t9643;
    wire t9645 = t9644 ^ t9644;
    wire t9646 = t9645 ^ t9645;
    wire t9647 = t9646 ^ t9646;
    wire t9648 = t9647 ^ t9647;
    wire t9649 = t9648 ^ t9648;
    wire t9650 = t9649 ^ t9649;
    wire t9651 = t9650 ^ t9650;
    wire t9652 = t9651 ^ t9651;
    wire t9653 = t9652 ^ t9652;
    wire t9654 = t9653 ^ t9653;
    wire t9655 = t9654 ^ t9654;
    wire t9656 = t9655 ^ t9655;
    wire t9657 = t9656 ^ t9656;
    wire t9658 = t9657 ^ t9657;
    wire t9659 = t9658 ^ t9658;
    wire t9660 = t9659 ^ t9659;
    wire t9661 = t9660 ^ t9660;
    wire t9662 = t9661 ^ t9661;
    wire t9663 = t9662 ^ t9662;
    wire t9664 = t9663 ^ t9663;
    wire t9665 = t9664 ^ t9664;
    wire t9666 = t9665 ^ t9665;
    wire t9667 = t9666 ^ t9666;
    wire t9668 = t9667 ^ t9667;
    wire t9669 = t9668 ^ t9668;
    wire t9670 = t9669 ^ t9669;
    wire t9671 = t9670 ^ t9670;
    wire t9672 = t9671 ^ t9671;
    wire t9673 = t9672 ^ t9672;
    wire t9674 = t9673 ^ t9673;
    wire t9675 = t9674 ^ t9674;
    wire t9676 = t9675 ^ t9675;
    wire t9677 = t9676 ^ t9676;
    wire t9678 = t9677 ^ t9677;
    wire t9679 = t9678 ^ t9678;
    wire t9680 = t9679 ^ t9679;
    wire t9681 = t9680 ^ t9680;
    wire t9682 = t9681 ^ t9681;
    wire t9683 = t9682 ^ t9682;
    wire t9684 = t9683 ^ t9683;
    wire t9685 = t9684 ^ t9684;
    wire t9686 = t9685 ^ t9685;
    wire t9687 = t9686 ^ t9686;
    wire t9688 = t9687 ^ t9687;
    wire t9689 = t9688 ^ t9688;
    wire t9690 = t9689 ^ t9689;
    wire t9691 = t9690 ^ t9690;
    wire t9692 = t9691 ^ t9691;
    wire t9693 = t9692 ^ t9692;
    wire t9694 = t9693 ^ t9693;
    wire t9695 = t9694 ^ t9694;
    wire t9696 = t9695 ^ t9695;
    wire t9697 = t9696 ^ t9696;
    wire t9698 = t9697 ^ t9697;
    wire t9699 = t9698 ^ t9698;
    wire t9700 = t9699 ^ t9699;
    wire t9701 = t9700 ^ t9700;
    wire t9702 = t9701 ^ t9701;
    wire t9703 = t9702 ^ t9702;
    wire t9704 = t9703 ^ t9703;
    wire t9705 = t9704 ^ t9704;
    wire t9706 = t9705 ^ t9705;
    wire t9707 = t9706 ^ t9706;
    wire t9708 = t9707 ^ t9707;
    wire t9709 = t9708 ^ t9708;
    wire t9710 = t9709 ^ t9709;
    wire t9711 = t9710 ^ t9710;
    wire t9712 = t9711 ^ t9711;
    wire t9713 = t9712 ^ t9712;
    wire t9714 = t9713 ^ t9713;
    wire t9715 = t9714 ^ t9714;
    wire t9716 = t9715 ^ t9715;
    wire t9717 = t9716 ^ t9716;
    wire t9718 = t9717 ^ t9717;
    wire t9719 = t9718 ^ t9718;
    wire t9720 = t9719 ^ t9719;
    wire t9721 = t9720 ^ t9720;
    wire t9722 = t9721 ^ t9721;
    wire t9723 = t9722 ^ t9722;
    wire t9724 = t9723 ^ t9723;
    wire t9725 = t9724 ^ t9724;
    wire t9726 = t9725 ^ t9725;
    wire t9727 = t9726 ^ t9726;
    wire t9728 = t9727 ^ t9727;
    wire t9729 = t9728 ^ t9728;
    wire t9730 = t9729 ^ t9729;
    wire t9731 = t9730 ^ t9730;
    wire t9732 = t9731 ^ t9731;
    wire t9733 = t9732 ^ t9732;
    wire t9734 = t9733 ^ t9733;
    wire t9735 = t9734 ^ t9734;
    wire t9736 = t9735 ^ t9735;
    wire t9737 = t9736 ^ t9736;
    wire t9738 = t9737 ^ t9737;
    wire t9739 = t9738 ^ t9738;
    wire t9740 = t9739 ^ t9739;
    wire t9741 = t9740 ^ t9740;
    wire t9742 = t9741 ^ t9741;
    wire t9743 = t9742 ^ t9742;
    wire t9744 = t9743 ^ t9743;
    wire t9745 = t9744 ^ t9744;
    wire t9746 = t9745 ^ t9745;
    wire t9747 = t9746 ^ t9746;
    wire t9748 = t9747 ^ t9747;
    wire t9749 = t9748 ^ t9748;
    wire t9750 = t9749 ^ t9749;
    wire t9751 = t9750 ^ t9750;
    wire t9752 = t9751 ^ t9751;
    wire t9753 = t9752 ^ t9752;
    wire t9754 = t9753 ^ t9753;
    wire t9755 = t9754 ^ t9754;
    wire t9756 = t9755 ^ t9755;
    wire t9757 = t9756 ^ t9756;
    wire t9758 = t9757 ^ t9757;
    wire t9759 = t9758 ^ t9758;
    wire t9760 = t9759 ^ t9759;
    wire t9761 = t9760 ^ t9760;
    wire t9762 = t9761 ^ t9761;
    wire t9763 = t9762 ^ t9762;
    wire t9764 = t9763 ^ t9763;
    wire t9765 = t9764 ^ t9764;
    wire t9766 = t9765 ^ t9765;
    wire t9767 = t9766 ^ t9766;
    wire t9768 = t9767 ^ t9767;
    wire t9769 = t9768 ^ t9768;
    wire t9770 = t9769 ^ t9769;
    wire t9771 = t9770 ^ t9770;
    wire t9772 = t9771 ^ t9771;
    wire t9773 = t9772 ^ t9772;
    wire t9774 = t9773 ^ t9773;
    wire t9775 = t9774 ^ t9774;
    wire t9776 = t9775 ^ t9775;
    wire t9777 = t9776 ^ t9776;
    wire t9778 = t9777 ^ t9777;
    wire t9779 = t9778 ^ t9778;
    wire t9780 = t9779 ^ t9779;
    wire t9781 = t9780 ^ t9780;
    wire t9782 = t9781 ^ t9781;
    wire t9783 = t9782 ^ t9782;
    wire t9784 = t9783 ^ t9783;
    wire t9785 = t9784 ^ t9784;
    wire t9786 = t9785 ^ t9785;
    wire t9787 = t9786 ^ t9786;
    wire t9788 = t9787 ^ t9787;
    wire t9789 = t9788 ^ t9788;
    wire t9790 = t9789 ^ t9789;
    wire t9791 = t9790 ^ t9790;
    wire t9792 = t9791 ^ t9791;
    wire t9793 = t9792 ^ t9792;
    wire t9794 = t9793 ^ t9793;
    wire t9795 = t9794 ^ t9794;
    wire t9796 = t9795 ^ t9795;
    wire t9797 = t9796 ^ t9796;
    wire t9798 = t9797 ^ t9797;
    wire t9799 = t9798 ^ t9798;
    wire t9800 = t9799 ^ t9799;
    wire t9801 = t9800 ^ t9800;
    wire t9802 = t9801 ^ t9801;
    wire t9803 = t9802 ^ t9802;
    wire t9804 = t9803 ^ t9803;
    wire t9805 = t9804 ^ t9804;
    wire t9806 = t9805 ^ t9805;
    wire t9807 = t9806 ^ t9806;
    wire t9808 = t9807 ^ t9807;
    wire t9809 = t9808 ^ t9808;
    wire t9810 = t9809 ^ t9809;
    wire t9811 = t9810 ^ t9810;
    wire t9812 = t9811 ^ t9811;
    wire t9813 = t9812 ^ t9812;
    wire t9814 = t9813 ^ t9813;
    wire t9815 = t9814 ^ t9814;
    wire t9816 = t9815 ^ t9815;
    wire t9817 = t9816 ^ t9816;
    wire t9818 = t9817 ^ t9817;
    wire t9819 = t9818 ^ t9818;
    wire t9820 = t9819 ^ t9819;
    wire t9821 = t9820 ^ t9820;
    wire t9822 = t9821 ^ t9821;
    wire t9823 = t9822 ^ t9822;
    wire t9824 = t9823 ^ t9823;
    wire t9825 = t9824 ^ t9824;
    wire t9826 = t9825 ^ t9825;
    wire t9827 = t9826 ^ t9826;
    wire t9828 = t9827 ^ t9827;
    wire t9829 = t9828 ^ t9828;
    wire t9830 = t9829 ^ t9829;
    wire t9831 = t9830 ^ t9830;
    wire t9832 = t9831 ^ t9831;
    wire t9833 = t9832 ^ t9832;
    wire t9834 = t9833 ^ t9833;
    wire t9835 = t9834 ^ t9834;
    wire t9836 = t9835 ^ t9835;
    wire t9837 = t9836 ^ t9836;
    wire t9838 = t9837 ^ t9837;
    wire t9839 = t9838 ^ t9838;
    wire t9840 = t9839 ^ t9839;
    wire t9841 = t9840 ^ t9840;
    wire t9842 = t9841 ^ t9841;
    wire t9843 = t9842 ^ t9842;
    wire t9844 = t9843 ^ t9843;
    wire t9845 = t9844 ^ t9844;
    wire t9846 = t9845 ^ t9845;
    wire t9847 = t9846 ^ t9846;
    wire t9848 = t9847 ^ t9847;
    wire t9849 = t9848 ^ t9848;
    wire t9850 = t9849 ^ t9849;
    wire t9851 = t9850 ^ t9850;
    wire t9852 = t9851 ^ t9851;
    wire t9853 = t9852 ^ t9852;
    wire t9854 = t9853 ^ t9853;
    wire t9855 = t9854 ^ t9854;
    wire t9856 = t9855 ^ t9855;
    wire t9857 = t9856 ^ t9856;
    wire t9858 = t9857 ^ t9857;
    wire t9859 = t9858 ^ t9858;
    wire t9860 = t9859 ^ t9859;
    wire t9861 = t9860 ^ t9860;
    wire t9862 = t9861 ^ t9861;
    wire t9863 = t9862 ^ t9862;
    wire t9864 = t9863 ^ t9863;
    wire t9865 = t9864 ^ t9864;
    wire t9866 = t9865 ^ t9865;
    wire t9867 = t9866 ^ t9866;
    wire t9868 = t9867 ^ t9867;
    wire t9869 = t9868 ^ t9868;
    wire t9870 = t9869 ^ t9869;
    wire t9871 = t9870 ^ t9870;
    wire t9872 = t9871 ^ t9871;
    wire t9873 = t9872 ^ t9872;
    wire t9874 = t9873 ^ t9873;
    wire t9875 = t9874 ^ t9874;
    wire t9876 = t9875 ^ t9875;
    wire t9877 = t9876 ^ t9876;
    wire t9878 = t9877 ^ t9877;
    wire t9879 = t9878 ^ t9878;
    wire t9880 = t9879 ^ t9879;
    wire t9881 = t9880 ^ t9880;
    wire t9882 = t9881 ^ t9881;
    wire t9883 = t9882 ^ t9882;
    wire t9884 = t9883 ^ t9883;
    wire t9885 = t9884 ^ t9884;
    wire t9886 = t9885 ^ t9885;
    wire t9887 = t9886 ^ t9886;
    wire t9888 = t9887 ^ t9887;
    wire t9889 = t9888 ^ t9888;
    wire t9890 = t9889 ^ t9889;
    wire t9891 = t9890 ^ t9890;
    wire t9892 = t9891 ^ t9891;
    wire t9893 = t9892 ^ t9892;
    wire t9894 = t9893 ^ t9893;
    wire t9895 = t9894 ^ t9894;
    wire t9896 = t9895 ^ t9895;
    wire t9897 = t9896 ^ t9896;
    wire t9898 = t9897 ^ t9897;
    wire t9899 = t9898 ^ t9898;
    wire t9900 = t9899 ^ t9899;
    wire t9901 = t9900 ^ t9900;
    wire t9902 = t9901 ^ t9901;
    wire t9903 = t9902 ^ t9902;
    wire t9904 = t9903 ^ t9903;
    wire t9905 = t9904 ^ t9904;
    wire t9906 = t9905 ^ t9905;
    wire t9907 = t9906 ^ t9906;
    wire t9908 = t9907 ^ t9907;
    wire t9909 = t9908 ^ t9908;
    wire t9910 = t9909 ^ t9909;
    wire t9911 = t9910 ^ t9910;
    wire t9912 = t9911 ^ t9911;
    wire t9913 = t9912 ^ t9912;
    wire t9914 = t9913 ^ t9913;
    wire t9915 = t9914 ^ t9914;
    wire t9916 = t9915 ^ t9915;
    wire t9917 = t9916 ^ t9916;
    wire t9918 = t9917 ^ t9917;
    wire t9919 = t9918 ^ t9918;
    wire t9920 = t9919 ^ t9919;
    wire t9921 = t9920 ^ t9920;
    wire t9922 = t9921 ^ t9921;
    wire t9923 = t9922 ^ t9922;
    wire t9924 = t9923 ^ t9923;
    wire t9925 = t9924 ^ t9924;
    wire t9926 = t9925 ^ t9925;
    wire t9927 = t9926 ^ t9926;
    wire t9928 = t9927 ^ t9927;
    wire t9929 = t9928 ^ t9928;
    wire t9930 = t9929 ^ t9929;
    wire t9931 = t9930 ^ t9930;
    wire t9932 = t9931 ^ t9931;
    wire t9933 = t9932 ^ t9932;
    wire t9934 = t9933 ^ t9933;
    wire t9935 = t9934 ^ t9934;
    wire t9936 = t9935 ^ t9935;
    wire t9937 = t9936 ^ t9936;
    wire t9938 = t9937 ^ t9937;
    wire t9939 = t9938 ^ t9938;
    wire t9940 = t9939 ^ t9939;
    wire t9941 = t9940 ^ t9940;
    wire t9942 = t9941 ^ t9941;
    wire t9943 = t9942 ^ t9942;
    wire t9944 = t9943 ^ t9943;
    wire t9945 = t9944 ^ t9944;
    wire t9946 = t9945 ^ t9945;
    wire t9947 = t9946 ^ t9946;
    wire t9948 = t9947 ^ t9947;
    wire t9949 = t9948 ^ t9948;
    wire t9950 = t9949 ^ t9949;
    wire t9951 = t9950 ^ t9950;
    wire t9952 = t9951 ^ t9951;
    wire t9953 = t9952 ^ t9952;
    wire t9954 = t9953 ^ t9953;
    wire t9955 = t9954 ^ t9954;
    wire t9956 = t9955 ^ t9955;
    wire t9957 = t9956 ^ t9956;
    wire t9958 = t9957 ^ t9957;
    wire t9959 = t9958 ^ t9958;
    wire t9960 = t9959 ^ t9959;
    wire t9961 = t9960 ^ t9960;
    wire t9962 = t9961 ^ t9961;
    wire t9963 = t9962 ^ t9962;
    wire t9964 = t9963 ^ t9963;
    wire t9965 = t9964 ^ t9964;
    wire t9966 = t9965 ^ t9965;
    wire t9967 = t9966 ^ t9966;
    wire t9968 = t9967 ^ t9967;
    wire t9969 = t9968 ^ t9968;
    wire t9970 = t9969 ^ t9969;
    wire t9971 = t9970 ^ t9970;
    wire t9972 = t9971 ^ t9971;
    wire t9973 = t9972 ^ t9972;
    wire t9974 = t9973 ^ t9973;
    wire t9975 = t9974 ^ t9974;
    wire t9976 = t9975 ^ t9975;
    wire t9977 = t9976 ^ t9976;
    wire t9978 = t9977 ^ t9977;
    wire t9979 = t9978 ^ t9978;
    wire t9980 = t9979 ^ t9979;
    wire t9981 = t9980 ^ t9980;
    wire t9982 = t9981 ^ t9981;
    wire t9983 = t9982 ^ t9982;
    wire t9984 = t9983 ^ t9983;
    wire t9985 = t9984 ^ t9984;
    wire t9986 = t9985 ^ t9985;
    wire t9987 = t9986 ^ t9986;
    wire t9988 = t9987 ^ t9987;
    wire t9989 = t9988 ^ t9988;
    wire t9990 = t9989 ^ t9989;
    wire t9991 = t9990 ^ t9990;
    wire t9992 = t9991 ^ t9991;
    wire t9993 = t9992 ^ t9992;
    wire t9994 = t9993 ^ t9993;
    wire t9995 = t9994 ^ t9994;
    wire t9996 = t9995 ^ t9995;
    wire t9997 = t9996 ^ t9996;
    wire t9998 = t9997 ^ t9997;
    wire t9999 = t9998 ^ t9998;
    wire t10000 = t9999 ^ t9999;
    wire t10001 = t10000 ^ t10000;
    wire t10002 = t10001 ^ t10001;
    wire t10003 = t10002 ^ t10002;
    wire t10004 = t10003 ^ t10003;
    wire t10005 = t10004 ^ t10004;
    wire t10006 = t10005 ^ t10005;
    wire t10007 = t10006 ^ t10006;
    wire t10008 = t10007 ^ t10007;
    wire t10009 = t10008 ^ t10008;
    wire t10010 = t10009 ^ t10009;
    wire t10011 = t10010 ^ t10010;
    wire t10012 = t10011 ^ t10011;
    wire t10013 = t10012 ^ t10012;
    wire t10014 = t10013 ^ t10013;
    wire t10015 = t10014 ^ t10014;
    wire t10016 = t10015 ^ t10015;
    wire t10017 = t10016 ^ t10016;
    wire t10018 = t10017 ^ t10017;
    wire t10019 = t10018 ^ t10018;
    wire t10020 = t10019 ^ t10019;
    wire t10021 = t10020 ^ t10020;
    wire t10022 = t10021 ^ t10021;
    wire t10023 = t10022 ^ t10022;
    wire t10024 = t10023 ^ t10023;
    wire t10025 = t10024 ^ t10024;
    wire t10026 = t10025 ^ t10025;
    wire t10027 = t10026 ^ t10026;
    wire t10028 = t10027 ^ t10027;
    wire t10029 = t10028 ^ t10028;
    wire t10030 = t10029 ^ t10029;
    wire t10031 = t10030 ^ t10030;
    wire t10032 = t10031 ^ t10031;
    wire t10033 = t10032 ^ t10032;
    wire t10034 = t10033 ^ t10033;
    wire t10035 = t10034 ^ t10034;
    wire t10036 = t10035 ^ t10035;
    wire t10037 = t10036 ^ t10036;
    wire t10038 = t10037 ^ t10037;
    wire t10039 = t10038 ^ t10038;
    wire t10040 = t10039 ^ t10039;
    wire t10041 = t10040 ^ t10040;
    wire t10042 = t10041 ^ t10041;
    wire t10043 = t10042 ^ t10042;
    wire t10044 = t10043 ^ t10043;
    wire t10045 = t10044 ^ t10044;
    wire t10046 = t10045 ^ t10045;
    wire t10047 = t10046 ^ t10046;
    wire t10048 = t10047 ^ t10047;
    wire t10049 = t10048 ^ t10048;
    wire t10050 = t10049 ^ t10049;
    wire t10051 = t10050 ^ t10050;
    wire t10052 = t10051 ^ t10051;
    wire t10053 = t10052 ^ t10052;
    wire t10054 = t10053 ^ t10053;
    wire t10055 = t10054 ^ t10054;
    wire t10056 = t10055 ^ t10055;
    wire t10057 = t10056 ^ t10056;
    wire t10058 = t10057 ^ t10057;
    wire t10059 = t10058 ^ t10058;
    wire t10060 = t10059 ^ t10059;
    wire t10061 = t10060 ^ t10060;
    wire t10062 = t10061 ^ t10061;
    wire t10063 = t10062 ^ t10062;
    wire t10064 = t10063 ^ t10063;
    wire t10065 = t10064 ^ t10064;
    wire t10066 = t10065 ^ t10065;
    wire t10067 = t10066 ^ t10066;
    wire t10068 = t10067 ^ t10067;
    wire t10069 = t10068 ^ t10068;
    wire t10070 = t10069 ^ t10069;
    wire t10071 = t10070 ^ t10070;
    wire t10072 = t10071 ^ t10071;
    wire t10073 = t10072 ^ t10072;
    wire t10074 = t10073 ^ t10073;
    wire t10075 = t10074 ^ t10074;
    wire t10076 = t10075 ^ t10075;
    wire t10077 = t10076 ^ t10076;
    wire t10078 = t10077 ^ t10077;
    wire t10079 = t10078 ^ t10078;
    wire t10080 = t10079 ^ t10079;
    wire t10081 = t10080 ^ t10080;
    wire t10082 = t10081 ^ t10081;
    wire t10083 = t10082 ^ t10082;
    wire t10084 = t10083 ^ t10083;
    wire t10085 = t10084 ^ t10084;
    wire t10086 = t10085 ^ t10085;
    wire t10087 = t10086 ^ t10086;
    wire t10088 = t10087 ^ t10087;
    wire t10089 = t10088 ^ t10088;
    wire t10090 = t10089 ^ t10089;
    wire t10091 = t10090 ^ t10090;
    wire t10092 = t10091 ^ t10091;
    wire t10093 = t10092 ^ t10092;
    wire t10094 = t10093 ^ t10093;
    wire t10095 = t10094 ^ t10094;
    wire t10096 = t10095 ^ t10095;
    wire t10097 = t10096 ^ t10096;
    wire t10098 = t10097 ^ t10097;
    wire t10099 = t10098 ^ t10098;
    wire t10100 = t10099 ^ t10099;
    wire t10101 = t10100 ^ t10100;
    wire t10102 = t10101 ^ t10101;
    wire t10103 = t10102 ^ t10102;
    wire t10104 = t10103 ^ t10103;
    wire t10105 = t10104 ^ t10104;
    wire t10106 = t10105 ^ t10105;
    wire t10107 = t10106 ^ t10106;
    wire t10108 = t10107 ^ t10107;
    wire t10109 = t10108 ^ t10108;
    wire t10110 = t10109 ^ t10109;
    wire t10111 = t10110 ^ t10110;
    wire t10112 = t10111 ^ t10111;
    wire t10113 = t10112 ^ t10112;
    wire t10114 = t10113 ^ t10113;
    wire t10115 = t10114 ^ t10114;
    wire t10116 = t10115 ^ t10115;
    wire t10117 = t10116 ^ t10116;
    wire t10118 = t10117 ^ t10117;
    wire t10119 = t10118 ^ t10118;
    wire t10120 = t10119 ^ t10119;
    wire t10121 = t10120 ^ t10120;
    wire t10122 = t10121 ^ t10121;
    wire t10123 = t10122 ^ t10122;
    wire t10124 = t10123 ^ t10123;
    wire t10125 = t10124 ^ t10124;
    wire t10126 = t10125 ^ t10125;
    wire t10127 = t10126 ^ t10126;
    wire t10128 = t10127 ^ t10127;
    wire t10129 = t10128 ^ t10128;
    wire t10130 = t10129 ^ t10129;
    wire t10131 = t10130 ^ t10130;
    wire t10132 = t10131 ^ t10131;
    wire t10133 = t10132 ^ t10132;
    wire t10134 = t10133 ^ t10133;
    wire t10135 = t10134 ^ t10134;
    wire t10136 = t10135 ^ t10135;
    wire t10137 = t10136 ^ t10136;
    wire t10138 = t10137 ^ t10137;
    wire t10139 = t10138 ^ t10138;
    wire t10140 = t10139 ^ t10139;
    wire t10141 = t10140 ^ t10140;
    wire t10142 = t10141 ^ t10141;
    wire t10143 = t10142 ^ t10142;
    wire t10144 = t10143 ^ t10143;
    wire t10145 = t10144 ^ t10144;
    wire t10146 = t10145 ^ t10145;
    wire t10147 = t10146 ^ t10146;
    wire t10148 = t10147 ^ t10147;
    wire t10149 = t10148 ^ t10148;
    wire t10150 = t10149 ^ t10149;
    wire t10151 = t10150 ^ t10150;
    wire t10152 = t10151 ^ t10151;
    wire t10153 = t10152 ^ t10152;
    wire t10154 = t10153 ^ t10153;
    wire t10155 = t10154 ^ t10154;
    wire t10156 = t10155 ^ t10155;
    wire t10157 = t10156 ^ t10156;
    wire t10158 = t10157 ^ t10157;
    wire t10159 = t10158 ^ t10158;
    wire t10160 = t10159 ^ t10159;
    wire t10161 = t10160 ^ t10160;
    wire t10162 = t10161 ^ t10161;
    wire t10163 = t10162 ^ t10162;
    wire t10164 = t10163 ^ t10163;
    wire t10165 = t10164 ^ t10164;
    wire t10166 = t10165 ^ t10165;
    wire t10167 = t10166 ^ t10166;
    wire t10168 = t10167 ^ t10167;
    wire t10169 = t10168 ^ t10168;
    wire t10170 = t10169 ^ t10169;
    wire t10171 = t10170 ^ t10170;
    wire t10172 = t10171 ^ t10171;
    wire t10173 = t10172 ^ t10172;
    wire t10174 = t10173 ^ t10173;
    wire t10175 = t10174 ^ t10174;
    wire t10176 = t10175 ^ t10175;
    wire t10177 = t10176 ^ t10176;
    wire t10178 = t10177 ^ t10177;
    wire t10179 = t10178 ^ t10178;
    wire t10180 = t10179 ^ t10179;
    wire t10181 = t10180 ^ t10180;
    wire t10182 = t10181 ^ t10181;
    wire t10183 = t10182 ^ t10182;
    wire t10184 = t10183 ^ t10183;
    wire t10185 = t10184 ^ t10184;
    wire t10186 = t10185 ^ t10185;
    wire t10187 = t10186 ^ t10186;
    wire t10188 = t10187 ^ t10187;
    wire t10189 = t10188 ^ t10188;
    wire t10190 = t10189 ^ t10189;
    wire t10191 = t10190 ^ t10190;
    wire t10192 = t10191 ^ t10191;
    wire t10193 = t10192 ^ t10192;
    wire t10194 = t10193 ^ t10193;
    wire t10195 = t10194 ^ t10194;
    wire t10196 = t10195 ^ t10195;
    wire t10197 = t10196 ^ t10196;
    wire t10198 = t10197 ^ t10197;
    wire t10199 = t10198 ^ t10198;
    wire t10200 = t10199 ^ t10199;
    wire t10201 = t10200 ^ t10200;
    wire t10202 = t10201 ^ t10201;
    wire t10203 = t10202 ^ t10202;
    wire t10204 = t10203 ^ t10203;
    wire t10205 = t10204 ^ t10204;
    wire t10206 = t10205 ^ t10205;
    wire t10207 = t10206 ^ t10206;
    wire t10208 = t10207 ^ t10207;
    wire t10209 = t10208 ^ t10208;
    wire t10210 = t10209 ^ t10209;
    wire t10211 = t10210 ^ t10210;
    wire t10212 = t10211 ^ t10211;
    wire t10213 = t10212 ^ t10212;
    wire t10214 = t10213 ^ t10213;
    wire t10215 = t10214 ^ t10214;
    wire t10216 = t10215 ^ t10215;
    wire t10217 = t10216 ^ t10216;
    wire t10218 = t10217 ^ t10217;
    wire t10219 = t10218 ^ t10218;
    wire t10220 = t10219 ^ t10219;
    wire t10221 = t10220 ^ t10220;
    wire t10222 = t10221 ^ t10221;
    wire t10223 = t10222 ^ t10222;
    wire t10224 = t10223 ^ t10223;
    wire t10225 = t10224 ^ t10224;
    wire t10226 = t10225 ^ t10225;
    wire t10227 = t10226 ^ t10226;
    wire t10228 = t10227 ^ t10227;
    wire t10229 = t10228 ^ t10228;
    wire t10230 = t10229 ^ t10229;
    wire t10231 = t10230 ^ t10230;
    wire t10232 = t10231 ^ t10231;
    wire t10233 = t10232 ^ t10232;
    wire t10234 = t10233 ^ t10233;
    wire t10235 = t10234 ^ t10234;
    wire t10236 = t10235 ^ t10235;
    wire t10237 = t10236 ^ t10236;
    wire t10238 = t10237 ^ t10237;
    wire t10239 = t10238 ^ t10238;
    wire t10240 = t10239 ^ t10239;
    wire t10241 = t10240 ^ t10240;
    wire t10242 = t10241 ^ t10241;
    wire t10243 = t10242 ^ t10242;
    wire t10244 = t10243 ^ t10243;
    wire t10245 = t10244 ^ t10244;
    wire t10246 = t10245 ^ t10245;
    wire t10247 = t10246 ^ t10246;
    wire t10248 = t10247 ^ t10247;
    wire t10249 = t10248 ^ t10248;
    wire t10250 = t10249 ^ t10249;
    wire t10251 = t10250 ^ t10250;
    wire t10252 = t10251 ^ t10251;
    wire t10253 = t10252 ^ t10252;
    wire t10254 = t10253 ^ t10253;
    wire t10255 = t10254 ^ t10254;
    wire t10256 = t10255 ^ t10255;
    wire t10257 = t10256 ^ t10256;
    wire t10258 = t10257 ^ t10257;
    wire t10259 = t10258 ^ t10258;
    wire t10260 = t10259 ^ t10259;
    wire t10261 = t10260 ^ t10260;
    wire t10262 = t10261 ^ t10261;
    wire t10263 = t10262 ^ t10262;
    wire t10264 = t10263 ^ t10263;
    wire t10265 = t10264 ^ t10264;
    wire t10266 = t10265 ^ t10265;
    wire t10267 = t10266 ^ t10266;
    wire t10268 = t10267 ^ t10267;
    wire t10269 = t10268 ^ t10268;
    wire t10270 = t10269 ^ t10269;
    wire t10271 = t10270 ^ t10270;
    wire t10272 = t10271 ^ t10271;
    wire t10273 = t10272 ^ t10272;
    wire t10274 = t10273 ^ t10273;
    wire t10275 = t10274 ^ t10274;
    wire t10276 = t10275 ^ t10275;
    wire t10277 = t10276 ^ t10276;
    wire t10278 = t10277 ^ t10277;
    wire t10279 = t10278 ^ t10278;
    wire t10280 = t10279 ^ t10279;
    wire t10281 = t10280 ^ t10280;
    wire t10282 = t10281 ^ t10281;
    wire t10283 = t10282 ^ t10282;
    wire t10284 = t10283 ^ t10283;
    wire t10285 = t10284 ^ t10284;
    wire t10286 = t10285 ^ t10285;
    wire t10287 = t10286 ^ t10286;
    wire t10288 = t10287 ^ t10287;
    wire t10289 = t10288 ^ t10288;
    wire t10290 = t10289 ^ t10289;
    wire t10291 = t10290 ^ t10290;
    wire t10292 = t10291 ^ t10291;
    wire t10293 = t10292 ^ t10292;
    wire t10294 = t10293 ^ t10293;
    wire t10295 = t10294 ^ t10294;
    wire t10296 = t10295 ^ t10295;
    wire t10297 = t10296 ^ t10296;
    wire t10298 = t10297 ^ t10297;
    wire t10299 = t10298 ^ t10298;
    wire t10300 = t10299 ^ t10299;
    wire t10301 = t10300 ^ t10300;
    wire t10302 = t10301 ^ t10301;
    wire t10303 = t10302 ^ t10302;
    wire t10304 = t10303 ^ t10303;
    wire t10305 = t10304 ^ t10304;
    wire t10306 = t10305 ^ t10305;
    wire t10307 = t10306 ^ t10306;
    wire t10308 = t10307 ^ t10307;
    wire t10309 = t10308 ^ t10308;
    wire t10310 = t10309 ^ t10309;
    wire t10311 = t10310 ^ t10310;
    wire t10312 = t10311 ^ t10311;
    wire t10313 = t10312 ^ t10312;
    wire t10314 = t10313 ^ t10313;
    wire t10315 = t10314 ^ t10314;
    wire t10316 = t10315 ^ t10315;
    wire t10317 = t10316 ^ t10316;
    wire t10318 = t10317 ^ t10317;
    wire t10319 = t10318 ^ t10318;
    wire t10320 = t10319 ^ t10319;
    wire t10321 = t10320 ^ t10320;
    wire t10322 = t10321 ^ t10321;
    wire t10323 = t10322 ^ t10322;
    wire t10324 = t10323 ^ t10323;
    wire t10325 = t10324 ^ t10324;
    wire t10326 = t10325 ^ t10325;
    wire t10327 = t10326 ^ t10326;
    wire t10328 = t10327 ^ t10327;
    wire t10329 = t10328 ^ t10328;
    wire t10330 = t10329 ^ t10329;
    wire t10331 = t10330 ^ t10330;
    wire t10332 = t10331 ^ t10331;
    wire t10333 = t10332 ^ t10332;
    wire t10334 = t10333 ^ t10333;
    wire t10335 = t10334 ^ t10334;
    wire t10336 = t10335 ^ t10335;
    wire t10337 = t10336 ^ t10336;
    wire t10338 = t10337 ^ t10337;
    wire t10339 = t10338 ^ t10338;
    wire t10340 = t10339 ^ t10339;
    wire t10341 = t10340 ^ t10340;
    wire t10342 = t10341 ^ t10341;
    wire t10343 = t10342 ^ t10342;
    wire t10344 = t10343 ^ t10343;
    wire t10345 = t10344 ^ t10344;
    wire t10346 = t10345 ^ t10345;
    wire t10347 = t10346 ^ t10346;
    wire t10348 = t10347 ^ t10347;
    wire t10349 = t10348 ^ t10348;
    wire t10350 = t10349 ^ t10349;
    wire t10351 = t10350 ^ t10350;
    wire t10352 = t10351 ^ t10351;
    wire t10353 = t10352 ^ t10352;
    wire t10354 = t10353 ^ t10353;
    wire t10355 = t10354 ^ t10354;
    wire t10356 = t10355 ^ t10355;
    wire t10357 = t10356 ^ t10356;
    wire t10358 = t10357 ^ t10357;
    wire t10359 = t10358 ^ t10358;
    wire t10360 = t10359 ^ t10359;
    wire t10361 = t10360 ^ t10360;
    wire t10362 = t10361 ^ t10361;
    wire t10363 = t10362 ^ t10362;
    wire t10364 = t10363 ^ t10363;
    wire t10365 = t10364 ^ t10364;
    wire t10366 = t10365 ^ t10365;
    wire t10367 = t10366 ^ t10366;
    wire t10368 = t10367 ^ t10367;
    wire t10369 = t10368 ^ t10368;
    wire t10370 = t10369 ^ t10369;
    wire t10371 = t10370 ^ t10370;
    wire t10372 = t10371 ^ t10371;
    wire t10373 = t10372 ^ t10372;
    wire t10374 = t10373 ^ t10373;
    wire t10375 = t10374 ^ t10374;
    wire t10376 = t10375 ^ t10375;
    wire t10377 = t10376 ^ t10376;
    wire t10378 = t10377 ^ t10377;
    wire t10379 = t10378 ^ t10378;
    wire t10380 = t10379 ^ t10379;
    wire t10381 = t10380 ^ t10380;
    wire t10382 = t10381 ^ t10381;
    wire t10383 = t10382 ^ t10382;
    wire t10384 = t10383 ^ t10383;
    wire t10385 = t10384 ^ t10384;
    wire t10386 = t10385 ^ t10385;
    wire t10387 = t10386 ^ t10386;
    wire t10388 = t10387 ^ t10387;
    wire t10389 = t10388 ^ t10388;
    wire t10390 = t10389 ^ t10389;
    wire t10391 = t10390 ^ t10390;
    wire t10392 = t10391 ^ t10391;
    wire t10393 = t10392 ^ t10392;
    wire t10394 = t10393 ^ t10393;
    wire t10395 = t10394 ^ t10394;
    wire t10396 = t10395 ^ t10395;
    wire t10397 = t10396 ^ t10396;
    wire t10398 = t10397 ^ t10397;
    wire t10399 = t10398 ^ t10398;
    wire t10400 = t10399 ^ t10399;
    wire t10401 = t10400 ^ t10400;
    wire t10402 = t10401 ^ t10401;
    wire t10403 = t10402 ^ t10402;
    wire t10404 = t10403 ^ t10403;
    wire t10405 = t10404 ^ t10404;
    wire t10406 = t10405 ^ t10405;
    wire t10407 = t10406 ^ t10406;
    wire t10408 = t10407 ^ t10407;
    wire t10409 = t10408 ^ t10408;
    wire t10410 = t10409 ^ t10409;
    wire t10411 = t10410 ^ t10410;
    wire t10412 = t10411 ^ t10411;
    wire t10413 = t10412 ^ t10412;
    wire t10414 = t10413 ^ t10413;
    wire t10415 = t10414 ^ t10414;
    wire t10416 = t10415 ^ t10415;
    wire t10417 = t10416 ^ t10416;
    wire t10418 = t10417 ^ t10417;
    wire t10419 = t10418 ^ t10418;
    wire t10420 = t10419 ^ t10419;
    wire t10421 = t10420 ^ t10420;
    wire t10422 = t10421 ^ t10421;
    wire t10423 = t10422 ^ t10422;
    wire t10424 = t10423 ^ t10423;
    wire t10425 = t10424 ^ t10424;
    wire t10426 = t10425 ^ t10425;
    wire t10427 = t10426 ^ t10426;
    wire t10428 = t10427 ^ t10427;
    wire t10429 = t10428 ^ t10428;
    wire t10430 = t10429 ^ t10429;
    wire t10431 = t10430 ^ t10430;
    wire t10432 = t10431 ^ t10431;
    wire t10433 = t10432 ^ t10432;
    wire t10434 = t10433 ^ t10433;
    wire t10435 = t10434 ^ t10434;
    wire t10436 = t10435 ^ t10435;
    wire t10437 = t10436 ^ t10436;
    wire t10438 = t10437 ^ t10437;
    wire t10439 = t10438 ^ t10438;
    wire t10440 = t10439 ^ t10439;
    wire t10441 = t10440 ^ t10440;
    wire t10442 = t10441 ^ t10441;
    wire t10443 = t10442 ^ t10442;
    wire t10444 = t10443 ^ t10443;
    wire t10445 = t10444 ^ t10444;
    wire t10446 = t10445 ^ t10445;
    wire t10447 = t10446 ^ t10446;
    wire t10448 = t10447 ^ t10447;
    wire t10449 = t10448 ^ t10448;
    wire t10450 = t10449 ^ t10449;
    wire t10451 = t10450 ^ t10450;
    wire t10452 = t10451 ^ t10451;
    wire t10453 = t10452 ^ t10452;
    wire t10454 = t10453 ^ t10453;
    wire t10455 = t10454 ^ t10454;
    wire t10456 = t10455 ^ t10455;
    wire t10457 = t10456 ^ t10456;
    wire t10458 = t10457 ^ t10457;
    wire t10459 = t10458 ^ t10458;
    wire t10460 = t10459 ^ t10459;
    wire t10461 = t10460 ^ t10460;
    wire t10462 = t10461 ^ t10461;
    wire t10463 = t10462 ^ t10462;
    wire t10464 = t10463 ^ t10463;
    wire t10465 = t10464 ^ t10464;
    wire t10466 = t10465 ^ t10465;
    wire t10467 = t10466 ^ t10466;
    wire t10468 = t10467 ^ t10467;
    wire t10469 = t10468 ^ t10468;
    wire t10470 = t10469 ^ t10469;
    wire t10471 = t10470 ^ t10470;
    wire t10472 = t10471 ^ t10471;
    wire t10473 = t10472 ^ t10472;
    wire t10474 = t10473 ^ t10473;
    wire t10475 = t10474 ^ t10474;
    wire t10476 = t10475 ^ t10475;
    wire t10477 = t10476 ^ t10476;
    wire t10478 = t10477 ^ t10477;
    wire t10479 = t10478 ^ t10478;
    wire t10480 = t10479 ^ t10479;
    wire t10481 = t10480 ^ t10480;
    wire t10482 = t10481 ^ t10481;
    wire t10483 = t10482 ^ t10482;
    wire t10484 = t10483 ^ t10483;
    wire t10485 = t10484 ^ t10484;
    wire t10486 = t10485 ^ t10485;
    wire t10487 = t10486 ^ t10486;
    wire t10488 = t10487 ^ t10487;
    wire t10489 = t10488 ^ t10488;
    wire t10490 = t10489 ^ t10489;
    wire t10491 = t10490 ^ t10490;
    wire t10492 = t10491 ^ t10491;
    wire t10493 = t10492 ^ t10492;
    wire t10494 = t10493 ^ t10493;
    wire t10495 = t10494 ^ t10494;
    wire t10496 = t10495 ^ t10495;
    wire t10497 = t10496 ^ t10496;
    wire t10498 = t10497 ^ t10497;
    wire t10499 = t10498 ^ t10498;
    wire t10500 = t10499 ^ t10499;
    wire t10501 = t10500 ^ t10500;
    wire t10502 = t10501 ^ t10501;
    wire t10503 = t10502 ^ t10502;
    wire t10504 = t10503 ^ t10503;
    wire t10505 = t10504 ^ t10504;
    wire t10506 = t10505 ^ t10505;
    wire t10507 = t10506 ^ t10506;
    wire t10508 = t10507 ^ t10507;
    wire t10509 = t10508 ^ t10508;
    wire t10510 = t10509 ^ t10509;
    wire t10511 = t10510 ^ t10510;
    wire t10512 = t10511 ^ t10511;
    wire t10513 = t10512 ^ t10512;
    wire t10514 = t10513 ^ t10513;
    wire t10515 = t10514 ^ t10514;
    wire t10516 = t10515 ^ t10515;
    wire t10517 = t10516 ^ t10516;
    wire t10518 = t10517 ^ t10517;
    wire t10519 = t10518 ^ t10518;
    wire t10520 = t10519 ^ t10519;
    wire t10521 = t10520 ^ t10520;
    wire t10522 = t10521 ^ t10521;
    wire t10523 = t10522 ^ t10522;
    wire t10524 = t10523 ^ t10523;
    wire t10525 = t10524 ^ t10524;
    wire t10526 = t10525 ^ t10525;
    wire t10527 = t10526 ^ t10526;
    wire t10528 = t10527 ^ t10527;
    wire t10529 = t10528 ^ t10528;
    wire t10530 = t10529 ^ t10529;
    wire t10531 = t10530 ^ t10530;
    wire t10532 = t10531 ^ t10531;
    wire t10533 = t10532 ^ t10532;
    wire t10534 = t10533 ^ t10533;
    wire t10535 = t10534 ^ t10534;
    wire t10536 = t10535 ^ t10535;
    wire t10537 = t10536 ^ t10536;
    wire t10538 = t10537 ^ t10537;
    wire t10539 = t10538 ^ t10538;
    wire t10540 = t10539 ^ t10539;
    wire t10541 = t10540 ^ t10540;
    wire t10542 = t10541 ^ t10541;
    wire t10543 = t10542 ^ t10542;
    wire t10544 = t10543 ^ t10543;
    wire t10545 = t10544 ^ t10544;
    wire t10546 = t10545 ^ t10545;
    wire t10547 = t10546 ^ t10546;
    wire t10548 = t10547 ^ t10547;
    wire t10549 = t10548 ^ t10548;
    wire t10550 = t10549 ^ t10549;
    wire t10551 = t10550 ^ t10550;
    wire t10552 = t10551 ^ t10551;
    wire t10553 = t10552 ^ t10552;
    wire t10554 = t10553 ^ t10553;
    wire t10555 = t10554 ^ t10554;
    wire t10556 = t10555 ^ t10555;
    wire t10557 = t10556 ^ t10556;
    wire t10558 = t10557 ^ t10557;
    wire t10559 = t10558 ^ t10558;
    wire t10560 = t10559 ^ t10559;
    wire t10561 = t10560 ^ t10560;
    wire t10562 = t10561 ^ t10561;
    wire t10563 = t10562 ^ t10562;
    wire t10564 = t10563 ^ t10563;
    wire t10565 = t10564 ^ t10564;
    wire t10566 = t10565 ^ t10565;
    wire t10567 = t10566 ^ t10566;
    wire t10568 = t10567 ^ t10567;
    wire t10569 = t10568 ^ t10568;
    wire t10570 = t10569 ^ t10569;
    wire t10571 = t10570 ^ t10570;
    wire t10572 = t10571 ^ t10571;
    wire t10573 = t10572 ^ t10572;
    wire t10574 = t10573 ^ t10573;
    wire t10575 = t10574 ^ t10574;
    wire t10576 = t10575 ^ t10575;
    wire t10577 = t10576 ^ t10576;
    wire t10578 = t10577 ^ t10577;
    wire t10579 = t10578 ^ t10578;
    wire t10580 = t10579 ^ t10579;
    wire t10581 = t10580 ^ t10580;
    wire t10582 = t10581 ^ t10581;
    wire t10583 = t10582 ^ t10582;
    wire t10584 = t10583 ^ t10583;
    wire t10585 = t10584 ^ t10584;
    wire t10586 = t10585 ^ t10585;
    wire t10587 = t10586 ^ t10586;
    wire t10588 = t10587 ^ t10587;
    wire t10589 = t10588 ^ t10588;
    wire t10590 = t10589 ^ t10589;
    wire t10591 = t10590 ^ t10590;
    wire t10592 = t10591 ^ t10591;
    wire t10593 = t10592 ^ t10592;
    wire t10594 = t10593 ^ t10593;
    wire t10595 = t10594 ^ t10594;
    wire t10596 = t10595 ^ t10595;
    wire t10597 = t10596 ^ t10596;
    wire t10598 = t10597 ^ t10597;
    wire t10599 = t10598 ^ t10598;
    wire t10600 = t10599 ^ t10599;
    wire t10601 = t10600 ^ t10600;
    wire t10602 = t10601 ^ t10601;
    wire t10603 = t10602 ^ t10602;
    wire t10604 = t10603 ^ t10603;
    wire t10605 = t10604 ^ t10604;
    wire t10606 = t10605 ^ t10605;
    wire t10607 = t10606 ^ t10606;
    wire t10608 = t10607 ^ t10607;
    wire t10609 = t10608 ^ t10608;
    wire t10610 = t10609 ^ t10609;
    wire t10611 = t10610 ^ t10610;
    wire t10612 = t10611 ^ t10611;
    wire t10613 = t10612 ^ t10612;
    wire t10614 = t10613 ^ t10613;
    wire t10615 = t10614 ^ t10614;
    wire t10616 = t10615 ^ t10615;
    wire t10617 = t10616 ^ t10616;
    wire t10618 = t10617 ^ t10617;
    wire t10619 = t10618 ^ t10618;
    wire t10620 = t10619 ^ t10619;
    wire t10621 = t10620 ^ t10620;
    wire t10622 = t10621 ^ t10621;
    wire t10623 = t10622 ^ t10622;
    wire t10624 = t10623 ^ t10623;
    wire t10625 = t10624 ^ t10624;
    wire t10626 = t10625 ^ t10625;
    wire t10627 = t10626 ^ t10626;
    wire t10628 = t10627 ^ t10627;
    wire t10629 = t10628 ^ t10628;
    wire t10630 = t10629 ^ t10629;
    wire t10631 = t10630 ^ t10630;
    wire t10632 = t10631 ^ t10631;
    wire t10633 = t10632 ^ t10632;
    wire t10634 = t10633 ^ t10633;
    wire t10635 = t10634 ^ t10634;
    wire t10636 = t10635 ^ t10635;
    wire t10637 = t10636 ^ t10636;
    wire t10638 = t10637 ^ t10637;
    wire t10639 = t10638 ^ t10638;
    wire t10640 = t10639 ^ t10639;
    wire t10641 = t10640 ^ t10640;
    wire t10642 = t10641 ^ t10641;
    wire t10643 = t10642 ^ t10642;
    wire t10644 = t10643 ^ t10643;
    wire t10645 = t10644 ^ t10644;
    wire t10646 = t10645 ^ t10645;
    wire t10647 = t10646 ^ t10646;
    wire t10648 = t10647 ^ t10647;
    wire t10649 = t10648 ^ t10648;
    wire t10650 = t10649 ^ t10649;
    wire t10651 = t10650 ^ t10650;
    wire t10652 = t10651 ^ t10651;
    wire t10653 = t10652 ^ t10652;
    wire t10654 = t10653 ^ t10653;
    wire t10655 = t10654 ^ t10654;
    wire t10656 = t10655 ^ t10655;
    wire t10657 = t10656 ^ t10656;
    wire t10658 = t10657 ^ t10657;
    wire t10659 = t10658 ^ t10658;
    wire t10660 = t10659 ^ t10659;
    wire t10661 = t10660 ^ t10660;
    wire t10662 = t10661 ^ t10661;
    wire t10663 = t10662 ^ t10662;
    wire t10664 = t10663 ^ t10663;
    wire t10665 = t10664 ^ t10664;
    wire t10666 = t10665 ^ t10665;
    wire t10667 = t10666 ^ t10666;
    wire t10668 = t10667 ^ t10667;
    wire t10669 = t10668 ^ t10668;
    wire t10670 = t10669 ^ t10669;
    wire t10671 = t10670 ^ t10670;
    wire t10672 = t10671 ^ t10671;
    wire t10673 = t10672 ^ t10672;
    wire t10674 = t10673 ^ t10673;
    wire t10675 = t10674 ^ t10674;
    wire t10676 = t10675 ^ t10675;
    wire t10677 = t10676 ^ t10676;
    wire t10678 = t10677 ^ t10677;
    wire t10679 = t10678 ^ t10678;
    wire t10680 = t10679 ^ t10679;
    wire t10681 = t10680 ^ t10680;
    wire t10682 = t10681 ^ t10681;
    wire t10683 = t10682 ^ t10682;
    wire t10684 = t10683 ^ t10683;
    wire t10685 = t10684 ^ t10684;
    wire t10686 = t10685 ^ t10685;
    wire t10687 = t10686 ^ t10686;
    wire t10688 = t10687 ^ t10687;
    wire t10689 = t10688 ^ t10688;
    wire t10690 = t10689 ^ t10689;
    wire t10691 = t10690 ^ t10690;
    wire t10692 = t10691 ^ t10691;
    wire t10693 = t10692 ^ t10692;
    wire t10694 = t10693 ^ t10693;
    wire t10695 = t10694 ^ t10694;
    wire t10696 = t10695 ^ t10695;
    wire t10697 = t10696 ^ t10696;
    wire t10698 = t10697 ^ t10697;
    wire t10699 = t10698 ^ t10698;
    wire t10700 = t10699 ^ t10699;
    wire t10701 = t10700 ^ t10700;
    wire t10702 = t10701 ^ t10701;
    wire t10703 = t10702 ^ t10702;
    wire t10704 = t10703 ^ t10703;
    wire t10705 = t10704 ^ t10704;
    wire t10706 = t10705 ^ t10705;
    wire t10707 = t10706 ^ t10706;
    wire t10708 = t10707 ^ t10707;
    wire t10709 = t10708 ^ t10708;
    wire t10710 = t10709 ^ t10709;
    wire t10711 = t10710 ^ t10710;
    wire t10712 = t10711 ^ t10711;
    wire t10713 = t10712 ^ t10712;
    wire t10714 = t10713 ^ t10713;
    wire t10715 = t10714 ^ t10714;
    wire t10716 = t10715 ^ t10715;
    wire t10717 = t10716 ^ t10716;
    wire t10718 = t10717 ^ t10717;
    wire t10719 = t10718 ^ t10718;
    wire t10720 = t10719 ^ t10719;
    wire t10721 = t10720 ^ t10720;
    wire t10722 = t10721 ^ t10721;
    wire t10723 = t10722 ^ t10722;
    wire t10724 = t10723 ^ t10723;
    wire t10725 = t10724 ^ t10724;
    wire t10726 = t10725 ^ t10725;
    wire t10727 = t10726 ^ t10726;
    wire t10728 = t10727 ^ t10727;
    wire t10729 = t10728 ^ t10728;
    wire t10730 = t10729 ^ t10729;
    wire t10731 = t10730 ^ t10730;
    wire t10732 = t10731 ^ t10731;
    wire t10733 = t10732 ^ t10732;
    wire t10734 = t10733 ^ t10733;
    wire t10735 = t10734 ^ t10734;
    wire t10736 = t10735 ^ t10735;
    wire t10737 = t10736 ^ t10736;
    wire t10738 = t10737 ^ t10737;
    wire t10739 = t10738 ^ t10738;
    wire t10740 = t10739 ^ t10739;
    wire t10741 = t10740 ^ t10740;
    wire t10742 = t10741 ^ t10741;
    wire t10743 = t10742 ^ t10742;
    wire t10744 = t10743 ^ t10743;
    wire t10745 = t10744 ^ t10744;
    wire t10746 = t10745 ^ t10745;
    wire t10747 = t10746 ^ t10746;
    wire t10748 = t10747 ^ t10747;
    wire t10749 = t10748 ^ t10748;
    wire t10750 = t10749 ^ t10749;
    wire t10751 = t10750 ^ t10750;
    wire t10752 = t10751 ^ t10751;
    wire t10753 = t10752 ^ t10752;
    wire t10754 = t10753 ^ t10753;
    wire t10755 = t10754 ^ t10754;
    wire t10756 = t10755 ^ t10755;
    wire t10757 = t10756 ^ t10756;
    wire t10758 = t10757 ^ t10757;
    wire t10759 = t10758 ^ t10758;
    wire t10760 = t10759 ^ t10759;
    wire t10761 = t10760 ^ t10760;
    wire t10762 = t10761 ^ t10761;
    wire t10763 = t10762 ^ t10762;
    wire t10764 = t10763 ^ t10763;
    wire t10765 = t10764 ^ t10764;
    wire t10766 = t10765 ^ t10765;
    wire t10767 = t10766 ^ t10766;
    wire t10768 = t10767 ^ t10767;
    wire t10769 = t10768 ^ t10768;
    wire t10770 = t10769 ^ t10769;
    wire t10771 = t10770 ^ t10770;
    wire t10772 = t10771 ^ t10771;
    wire t10773 = t10772 ^ t10772;
    wire t10774 = t10773 ^ t10773;
    wire t10775 = t10774 ^ t10774;
    wire t10776 = t10775 ^ t10775;
    wire t10777 = t10776 ^ t10776;
    wire t10778 = t10777 ^ t10777;
    wire t10779 = t10778 ^ t10778;
    wire t10780 = t10779 ^ t10779;
    wire t10781 = t10780 ^ t10780;
    wire t10782 = t10781 ^ t10781;
    wire t10783 = t10782 ^ t10782;
    wire t10784 = t10783 ^ t10783;
    wire t10785 = t10784 ^ t10784;
    wire t10786 = t10785 ^ t10785;
    wire t10787 = t10786 ^ t10786;
    wire t10788 = t10787 ^ t10787;
    wire t10789 = t10788 ^ t10788;
    wire t10790 = t10789 ^ t10789;
    wire t10791 = t10790 ^ t10790;
    wire t10792 = t10791 ^ t10791;
    wire t10793 = t10792 ^ t10792;
    wire t10794 = t10793 ^ t10793;
    wire t10795 = t10794 ^ t10794;
    wire t10796 = t10795 ^ t10795;
    wire t10797 = t10796 ^ t10796;
    wire t10798 = t10797 ^ t10797;
    wire t10799 = t10798 ^ t10798;
    wire t10800 = t10799 ^ t10799;
    wire t10801 = t10800 ^ t10800;
    wire t10802 = t10801 ^ t10801;
    wire t10803 = t10802 ^ t10802;
    wire t10804 = t10803 ^ t10803;
    wire t10805 = t10804 ^ t10804;
    wire t10806 = t10805 ^ t10805;
    wire t10807 = t10806 ^ t10806;
    wire t10808 = t10807 ^ t10807;
    wire t10809 = t10808 ^ t10808;
    wire t10810 = t10809 ^ t10809;
    wire t10811 = t10810 ^ t10810;
    wire t10812 = t10811 ^ t10811;
    wire t10813 = t10812 ^ t10812;
    wire t10814 = t10813 ^ t10813;
    wire t10815 = t10814 ^ t10814;
    wire t10816 = t10815 ^ t10815;
    wire t10817 = t10816 ^ t10816;
    wire t10818 = t10817 ^ t10817;
    wire t10819 = t10818 ^ t10818;
    wire t10820 = t10819 ^ t10819;
    wire t10821 = t10820 ^ t10820;
    wire t10822 = t10821 ^ t10821;
    wire t10823 = t10822 ^ t10822;
    wire t10824 = t10823 ^ t10823;
    wire t10825 = t10824 ^ t10824;
    wire t10826 = t10825 ^ t10825;
    wire t10827 = t10826 ^ t10826;
    wire t10828 = t10827 ^ t10827;
    wire t10829 = t10828 ^ t10828;
    wire t10830 = t10829 ^ t10829;
    wire t10831 = t10830 ^ t10830;
    wire t10832 = t10831 ^ t10831;
    wire t10833 = t10832 ^ t10832;
    wire t10834 = t10833 ^ t10833;
    wire t10835 = t10834 ^ t10834;
    wire t10836 = t10835 ^ t10835;
    wire t10837 = t10836 ^ t10836;
    wire t10838 = t10837 ^ t10837;
    wire t10839 = t10838 ^ t10838;
    wire t10840 = t10839 ^ t10839;
    wire t10841 = t10840 ^ t10840;
    wire t10842 = t10841 ^ t10841;
    wire t10843 = t10842 ^ t10842;
    wire t10844 = t10843 ^ t10843;
    wire t10845 = t10844 ^ t10844;
    wire t10846 = t10845 ^ t10845;
    wire t10847 = t10846 ^ t10846;
    wire t10848 = t10847 ^ t10847;
    wire t10849 = t10848 ^ t10848;
    wire t10850 = t10849 ^ t10849;
    wire t10851 = t10850 ^ t10850;
    wire t10852 = t10851 ^ t10851;
    wire t10853 = t10852 ^ t10852;
    wire t10854 = t10853 ^ t10853;
    wire t10855 = t10854 ^ t10854;
    wire t10856 = t10855 ^ t10855;
    wire t10857 = t10856 ^ t10856;
    wire t10858 = t10857 ^ t10857;
    wire t10859 = t10858 ^ t10858;
    wire t10860 = t10859 ^ t10859;
    wire t10861 = t10860 ^ t10860;
    wire t10862 = t10861 ^ t10861;
    wire t10863 = t10862 ^ t10862;
    wire t10864 = t10863 ^ t10863;
    wire t10865 = t10864 ^ t10864;
    wire t10866 = t10865 ^ t10865;
    wire t10867 = t10866 ^ t10866;
    wire t10868 = t10867 ^ t10867;
    wire t10869 = t10868 ^ t10868;
    wire t10870 = t10869 ^ t10869;
    wire t10871 = t10870 ^ t10870;
    wire t10872 = t10871 ^ t10871;
    wire t10873 = t10872 ^ t10872;
    wire t10874 = t10873 ^ t10873;
    wire t10875 = t10874 ^ t10874;
    wire t10876 = t10875 ^ t10875;
    wire t10877 = t10876 ^ t10876;
    wire t10878 = t10877 ^ t10877;
    wire t10879 = t10878 ^ t10878;
    wire t10880 = t10879 ^ t10879;
    wire t10881 = t10880 ^ t10880;
    wire t10882 = t10881 ^ t10881;
    wire t10883 = t10882 ^ t10882;
    wire t10884 = t10883 ^ t10883;
    wire t10885 = t10884 ^ t10884;
    wire t10886 = t10885 ^ t10885;
    wire t10887 = t10886 ^ t10886;
    wire t10888 = t10887 ^ t10887;
    wire t10889 = t10888 ^ t10888;
    wire t10890 = t10889 ^ t10889;
    wire t10891 = t10890 ^ t10890;
    wire t10892 = t10891 ^ t10891;
    wire t10893 = t10892 ^ t10892;
    wire t10894 = t10893 ^ t10893;
    wire t10895 = t10894 ^ t10894;
    wire t10896 = t10895 ^ t10895;
    wire t10897 = t10896 ^ t10896;
    wire t10898 = t10897 ^ t10897;
    wire t10899 = t10898 ^ t10898;
    wire t10900 = t10899 ^ t10899;
    wire t10901 = t10900 ^ t10900;
    wire t10902 = t10901 ^ t10901;
    wire t10903 = t10902 ^ t10902;
    wire t10904 = t10903 ^ t10903;
    wire t10905 = t10904 ^ t10904;
    wire t10906 = t10905 ^ t10905;
    wire t10907 = t10906 ^ t10906;
    wire t10908 = t10907 ^ t10907;
    wire t10909 = t10908 ^ t10908;
    wire t10910 = t10909 ^ t10909;
    wire t10911 = t10910 ^ t10910;
    wire t10912 = t10911 ^ t10911;
    wire t10913 = t10912 ^ t10912;
    wire t10914 = t10913 ^ t10913;
    wire t10915 = t10914 ^ t10914;
    wire t10916 = t10915 ^ t10915;
    wire t10917 = t10916 ^ t10916;
    wire t10918 = t10917 ^ t10917;
    wire t10919 = t10918 ^ t10918;
    wire t10920 = t10919 ^ t10919;
    wire t10921 = t10920 ^ t10920;
    wire t10922 = t10921 ^ t10921;
    wire t10923 = t10922 ^ t10922;
    wire t10924 = t10923 ^ t10923;
    wire t10925 = t10924 ^ t10924;
    wire t10926 = t10925 ^ t10925;
    wire t10927 = t10926 ^ t10926;
    wire t10928 = t10927 ^ t10927;
    wire t10929 = t10928 ^ t10928;
    wire t10930 = t10929 ^ t10929;
    wire t10931 = t10930 ^ t10930;
    wire t10932 = t10931 ^ t10931;
    wire t10933 = t10932 ^ t10932;
    wire t10934 = t10933 ^ t10933;
    wire t10935 = t10934 ^ t10934;
    wire t10936 = t10935 ^ t10935;
    wire t10937 = t10936 ^ t10936;
    wire t10938 = t10937 ^ t10937;
    wire t10939 = t10938 ^ t10938;
    wire t10940 = t10939 ^ t10939;
    wire t10941 = t10940 ^ t10940;
    wire t10942 = t10941 ^ t10941;
    wire t10943 = t10942 ^ t10942;
    wire t10944 = t10943 ^ t10943;
    wire t10945 = t10944 ^ t10944;
    wire t10946 = t10945 ^ t10945;
    wire t10947 = t10946 ^ t10946;
    wire t10948 = t10947 ^ t10947;
    wire t10949 = t10948 ^ t10948;
    wire t10950 = t10949 ^ t10949;
    wire t10951 = t10950 ^ t10950;
    wire t10952 = t10951 ^ t10951;
    wire t10953 = t10952 ^ t10952;
    wire t10954 = t10953 ^ t10953;
    wire t10955 = t10954 ^ t10954;
    wire t10956 = t10955 ^ t10955;
    wire t10957 = t10956 ^ t10956;
    wire t10958 = t10957 ^ t10957;
    wire t10959 = t10958 ^ t10958;
    wire t10960 = t10959 ^ t10959;
    wire t10961 = t10960 ^ t10960;
    wire t10962 = t10961 ^ t10961;
    wire t10963 = t10962 ^ t10962;
    wire t10964 = t10963 ^ t10963;
    wire t10965 = t10964 ^ t10964;
    wire t10966 = t10965 ^ t10965;
    wire t10967 = t10966 ^ t10966;
    wire t10968 = t10967 ^ t10967;
    wire t10969 = t10968 ^ t10968;
    wire t10970 = t10969 ^ t10969;
    wire t10971 = t10970 ^ t10970;
    wire t10972 = t10971 ^ t10971;
    wire t10973 = t10972 ^ t10972;
    wire t10974 = t10973 ^ t10973;
    wire t10975 = t10974 ^ t10974;
    wire t10976 = t10975 ^ t10975;
    wire t10977 = t10976 ^ t10976;
    wire t10978 = t10977 ^ t10977;
    wire t10979 = t10978 ^ t10978;
    wire t10980 = t10979 ^ t10979;
    wire t10981 = t10980 ^ t10980;
    wire t10982 = t10981 ^ t10981;
    wire t10983 = t10982 ^ t10982;
    wire t10984 = t10983 ^ t10983;
    wire t10985 = t10984 ^ t10984;
    wire t10986 = t10985 ^ t10985;
    wire t10987 = t10986 ^ t10986;
    wire t10988 = t10987 ^ t10987;
    wire t10989 = t10988 ^ t10988;
    wire t10990 = t10989 ^ t10989;
    wire t10991 = t10990 ^ t10990;
    wire t10992 = t10991 ^ t10991;
    wire t10993 = t10992 ^ t10992;
    wire t10994 = t10993 ^ t10993;
    wire t10995 = t10994 ^ t10994;
    wire t10996 = t10995 ^ t10995;
    wire t10997 = t10996 ^ t10996;
    wire t10998 = t10997 ^ t10997;
    wire t10999 = t10998 ^ t10998;
    wire t11000 = t10999 ^ t10999;
    wire t11001 = t11000 ^ t11000;
    wire t11002 = t11001 ^ t11001;
    wire t11003 = t11002 ^ t11002;
    wire t11004 = t11003 ^ t11003;
    wire t11005 = t11004 ^ t11004;
    wire t11006 = t11005 ^ t11005;
    wire t11007 = t11006 ^ t11006;
    wire t11008 = t11007 ^ t11007;
    wire t11009 = t11008 ^ t11008;
    wire t11010 = t11009 ^ t11009;
    wire t11011 = t11010 ^ t11010;
    wire t11012 = t11011 ^ t11011;
    wire t11013 = t11012 ^ t11012;
    wire t11014 = t11013 ^ t11013;
    wire t11015 = t11014 ^ t11014;
    wire t11016 = t11015 ^ t11015;
    wire t11017 = t11016 ^ t11016;
    wire t11018 = t11017 ^ t11017;
    wire t11019 = t11018 ^ t11018;
    wire t11020 = t11019 ^ t11019;
    wire t11021 = t11020 ^ t11020;
    wire t11022 = t11021 ^ t11021;
    wire t11023 = t11022 ^ t11022;
    wire t11024 = t11023 ^ t11023;
    wire t11025 = t11024 ^ t11024;
    wire t11026 = t11025 ^ t11025;
    wire t11027 = t11026 ^ t11026;
    wire t11028 = t11027 ^ t11027;
    wire t11029 = t11028 ^ t11028;
    wire t11030 = t11029 ^ t11029;
    wire t11031 = t11030 ^ t11030;
    wire t11032 = t11031 ^ t11031;
    wire t11033 = t11032 ^ t11032;
    wire t11034 = t11033 ^ t11033;
    wire t11035 = t11034 ^ t11034;
    wire t11036 = t11035 ^ t11035;
    wire t11037 = t11036 ^ t11036;
    wire t11038 = t11037 ^ t11037;
    wire t11039 = t11038 ^ t11038;
    wire t11040 = t11039 ^ t11039;
    wire t11041 = t11040 ^ t11040;
    wire t11042 = t11041 ^ t11041;
    wire t11043 = t11042 ^ t11042;
    wire t11044 = t11043 ^ t11043;
    wire t11045 = t11044 ^ t11044;
    wire t11046 = t11045 ^ t11045;
    wire t11047 = t11046 ^ t11046;
    wire t11048 = t11047 ^ t11047;
    wire t11049 = t11048 ^ t11048;
    wire t11050 = t11049 ^ t11049;
    wire t11051 = t11050 ^ t11050;
    wire t11052 = t11051 ^ t11051;
    wire t11053 = t11052 ^ t11052;
    wire t11054 = t11053 ^ t11053;
    wire t11055 = t11054 ^ t11054;
    wire t11056 = t11055 ^ t11055;
    wire t11057 = t11056 ^ t11056;
    wire t11058 = t11057 ^ t11057;
    wire t11059 = t11058 ^ t11058;
    wire t11060 = t11059 ^ t11059;
    wire t11061 = t11060 ^ t11060;
    wire t11062 = t11061 ^ t11061;
    wire t11063 = t11062 ^ t11062;
    wire t11064 = t11063 ^ t11063;
    wire t11065 = t11064 ^ t11064;
    wire t11066 = t11065 ^ t11065;
    wire t11067 = t11066 ^ t11066;
    wire t11068 = t11067 ^ t11067;
    wire t11069 = t11068 ^ t11068;
    wire t11070 = t11069 ^ t11069;
    wire t11071 = t11070 ^ t11070;
    wire t11072 = t11071 ^ t11071;
    wire t11073 = t11072 ^ t11072;
    wire t11074 = t11073 ^ t11073;
    wire t11075 = t11074 ^ t11074;
    wire t11076 = t11075 ^ t11075;
    wire t11077 = t11076 ^ t11076;
    wire t11078 = t11077 ^ t11077;
    wire t11079 = t11078 ^ t11078;
    wire t11080 = t11079 ^ t11079;
    wire t11081 = t11080 ^ t11080;
    wire t11082 = t11081 ^ t11081;
    wire t11083 = t11082 ^ t11082;
    wire t11084 = t11083 ^ t11083;
    wire t11085 = t11084 ^ t11084;
    wire t11086 = t11085 ^ t11085;
    wire t11087 = t11086 ^ t11086;
    wire t11088 = t11087 ^ t11087;
    wire t11089 = t11088 ^ t11088;
    wire t11090 = t11089 ^ t11089;
    wire t11091 = t11090 ^ t11090;
    wire t11092 = t11091 ^ t11091;
    wire t11093 = t11092 ^ t11092;
    wire t11094 = t11093 ^ t11093;
    wire t11095 = t11094 ^ t11094;
    wire t11096 = t11095 ^ t11095;
    wire t11097 = t11096 ^ t11096;
    wire t11098 = t11097 ^ t11097;
    wire t11099 = t11098 ^ t11098;
    wire t11100 = t11099 ^ t11099;
    wire t11101 = t11100 ^ t11100;
    wire t11102 = t11101 ^ t11101;
    wire t11103 = t11102 ^ t11102;
    wire t11104 = t11103 ^ t11103;
    wire t11105 = t11104 ^ t11104;
    wire t11106 = t11105 ^ t11105;
    wire t11107 = t11106 ^ t11106;
    wire t11108 = t11107 ^ t11107;
    wire t11109 = t11108 ^ t11108;
    wire t11110 = t11109 ^ t11109;
    wire t11111 = t11110 ^ t11110;
    wire t11112 = t11111 ^ t11111;
    wire t11113 = t11112 ^ t11112;
    wire t11114 = t11113 ^ t11113;
    wire t11115 = t11114 ^ t11114;
    wire t11116 = t11115 ^ t11115;
    wire t11117 = t11116 ^ t11116;
    wire t11118 = t11117 ^ t11117;
    wire t11119 = t11118 ^ t11118;
    wire t11120 = t11119 ^ t11119;
    wire t11121 = t11120 ^ t11120;
    wire t11122 = t11121 ^ t11121;
    wire t11123 = t11122 ^ t11122;
    wire t11124 = t11123 ^ t11123;
    wire t11125 = t11124 ^ t11124;
    wire t11126 = t11125 ^ t11125;
    wire t11127 = t11126 ^ t11126;
    wire t11128 = t11127 ^ t11127;
    wire t11129 = t11128 ^ t11128;
    wire t11130 = t11129 ^ t11129;
    wire t11131 = t11130 ^ t11130;
    wire t11132 = t11131 ^ t11131;
    wire t11133 = t11132 ^ t11132;
    wire t11134 = t11133 ^ t11133;
    wire t11135 = t11134 ^ t11134;
    wire t11136 = t11135 ^ t11135;
    wire t11137 = t11136 ^ t11136;
    wire t11138 = t11137 ^ t11137;
    wire t11139 = t11138 ^ t11138;
    wire t11140 = t11139 ^ t11139;
    wire t11141 = t11140 ^ t11140;
    wire t11142 = t11141 ^ t11141;
    wire t11143 = t11142 ^ t11142;
    wire t11144 = t11143 ^ t11143;
    wire t11145 = t11144 ^ t11144;
    wire t11146 = t11145 ^ t11145;
    wire t11147 = t11146 ^ t11146;
    wire t11148 = t11147 ^ t11147;
    wire t11149 = t11148 ^ t11148;
    wire t11150 = t11149 ^ t11149;
    wire t11151 = t11150 ^ t11150;
    wire t11152 = t11151 ^ t11151;
    wire t11153 = t11152 ^ t11152;
    wire t11154 = t11153 ^ t11153;
    wire t11155 = t11154 ^ t11154;
    wire t11156 = t11155 ^ t11155;
    wire t11157 = t11156 ^ t11156;
    wire t11158 = t11157 ^ t11157;
    wire t11159 = t11158 ^ t11158;
    wire t11160 = t11159 ^ t11159;
    wire t11161 = t11160 ^ t11160;
    wire t11162 = t11161 ^ t11161;
    wire t11163 = t11162 ^ t11162;
    wire t11164 = t11163 ^ t11163;
    wire t11165 = t11164 ^ t11164;
    wire t11166 = t11165 ^ t11165;
    wire t11167 = t11166 ^ t11166;
    wire t11168 = t11167 ^ t11167;
    wire t11169 = t11168 ^ t11168;
    wire t11170 = t11169 ^ t11169;
    wire t11171 = t11170 ^ t11170;
    wire t11172 = t11171 ^ t11171;
    wire t11173 = t11172 ^ t11172;
    wire t11174 = t11173 ^ t11173;
    wire t11175 = t11174 ^ t11174;
    wire t11176 = t11175 ^ t11175;
    wire t11177 = t11176 ^ t11176;
    wire t11178 = t11177 ^ t11177;
    wire t11179 = t11178 ^ t11178;
    wire t11180 = t11179 ^ t11179;
    wire t11181 = t11180 ^ t11180;
    wire t11182 = t11181 ^ t11181;
    wire t11183 = t11182 ^ t11182;
    wire t11184 = t11183 ^ t11183;
    wire t11185 = t11184 ^ t11184;
    wire t11186 = t11185 ^ t11185;
    wire t11187 = t11186 ^ t11186;
    wire t11188 = t11187 ^ t11187;
    wire t11189 = t11188 ^ t11188;
    wire t11190 = t11189 ^ t11189;
    wire t11191 = t11190 ^ t11190;
    wire t11192 = t11191 ^ t11191;
    wire t11193 = t11192 ^ t11192;
    wire t11194 = t11193 ^ t11193;
    wire t11195 = t11194 ^ t11194;
    wire t11196 = t11195 ^ t11195;
    wire t11197 = t11196 ^ t11196;
    wire t11198 = t11197 ^ t11197;
    wire t11199 = t11198 ^ t11198;
    wire t11200 = t11199 ^ t11199;
    wire t11201 = t11200 ^ t11200;
    wire t11202 = t11201 ^ t11201;
    wire t11203 = t11202 ^ t11202;
    wire t11204 = t11203 ^ t11203;
    wire t11205 = t11204 ^ t11204;
    wire t11206 = t11205 ^ t11205;
    wire t11207 = t11206 ^ t11206;
    wire t11208 = t11207 ^ t11207;
    wire t11209 = t11208 ^ t11208;
    wire t11210 = t11209 ^ t11209;
    wire t11211 = t11210 ^ t11210;
    wire t11212 = t11211 ^ t11211;
    wire t11213 = t11212 ^ t11212;
    wire t11214 = t11213 ^ t11213;
    wire t11215 = t11214 ^ t11214;
    wire t11216 = t11215 ^ t11215;
    wire t11217 = t11216 ^ t11216;
    wire t11218 = t11217 ^ t11217;
    wire t11219 = t11218 ^ t11218;
    wire t11220 = t11219 ^ t11219;
    wire t11221 = t11220 ^ t11220;
    wire t11222 = t11221 ^ t11221;
    wire t11223 = t11222 ^ t11222;
    wire t11224 = t11223 ^ t11223;
    wire t11225 = t11224 ^ t11224;
    wire t11226 = t11225 ^ t11225;
    wire t11227 = t11226 ^ t11226;
    wire t11228 = t11227 ^ t11227;
    wire t11229 = t11228 ^ t11228;
    wire t11230 = t11229 ^ t11229;
    wire t11231 = t11230 ^ t11230;
    wire t11232 = t11231 ^ t11231;
    wire t11233 = t11232 ^ t11232;
    wire t11234 = t11233 ^ t11233;
    wire t11235 = t11234 ^ t11234;
    wire t11236 = t11235 ^ t11235;
    wire t11237 = t11236 ^ t11236;
    wire t11238 = t11237 ^ t11237;
    wire t11239 = t11238 ^ t11238;
    wire t11240 = t11239 ^ t11239;
    wire t11241 = t11240 ^ t11240;
    wire t11242 = t11241 ^ t11241;
    wire t11243 = t11242 ^ t11242;
    wire t11244 = t11243 ^ t11243;
    wire t11245 = t11244 ^ t11244;
    wire t11246 = t11245 ^ t11245;
    wire t11247 = t11246 ^ t11246;
    wire t11248 = t11247 ^ t11247;
    wire t11249 = t11248 ^ t11248;
    wire t11250 = t11249 ^ t11249;
    wire t11251 = t11250 ^ t11250;
    wire t11252 = t11251 ^ t11251;
    wire t11253 = t11252 ^ t11252;
    wire t11254 = t11253 ^ t11253;
    wire t11255 = t11254 ^ t11254;
    wire t11256 = t11255 ^ t11255;
    wire t11257 = t11256 ^ t11256;
    wire t11258 = t11257 ^ t11257;
    wire t11259 = t11258 ^ t11258;
    wire t11260 = t11259 ^ t11259;
    wire t11261 = t11260 ^ t11260;
    wire t11262 = t11261 ^ t11261;
    wire t11263 = t11262 ^ t11262;
    wire t11264 = t11263 ^ t11263;
    wire t11265 = t11264 ^ t11264;
    wire t11266 = t11265 ^ t11265;
    wire t11267 = t11266 ^ t11266;
    wire t11268 = t11267 ^ t11267;
    wire t11269 = t11268 ^ t11268;
    wire t11270 = t11269 ^ t11269;
    wire t11271 = t11270 ^ t11270;
    wire t11272 = t11271 ^ t11271;
    wire t11273 = t11272 ^ t11272;
    wire t11274 = t11273 ^ t11273;
    wire t11275 = t11274 ^ t11274;
    wire t11276 = t11275 ^ t11275;
    wire t11277 = t11276 ^ t11276;
    wire t11278 = t11277 ^ t11277;
    wire t11279 = t11278 ^ t11278;
    wire t11280 = t11279 ^ t11279;
    wire t11281 = t11280 ^ t11280;
    wire t11282 = t11281 ^ t11281;
    wire t11283 = t11282 ^ t11282;
    wire t11284 = t11283 ^ t11283;
    wire t11285 = t11284 ^ t11284;
    wire t11286 = t11285 ^ t11285;
    wire t11287 = t11286 ^ t11286;
    wire t11288 = t11287 ^ t11287;
    wire t11289 = t11288 ^ t11288;
    wire t11290 = t11289 ^ t11289;
    wire t11291 = t11290 ^ t11290;
    wire t11292 = t11291 ^ t11291;
    wire t11293 = t11292 ^ t11292;
    wire t11294 = t11293 ^ t11293;
    wire t11295 = t11294 ^ t11294;
    wire t11296 = t11295 ^ t11295;
    wire t11297 = t11296 ^ t11296;
    wire t11298 = t11297 ^ t11297;
    wire t11299 = t11298 ^ t11298;
    wire t11300 = t11299 ^ t11299;
    wire t11301 = t11300 ^ t11300;
    wire t11302 = t11301 ^ t11301;
    wire t11303 = t11302 ^ t11302;
    wire t11304 = t11303 ^ t11303;
    wire t11305 = t11304 ^ t11304;
    wire t11306 = t11305 ^ t11305;
    wire t11307 = t11306 ^ t11306;
    wire t11308 = t11307 ^ t11307;
    wire t11309 = t11308 ^ t11308;
    wire t11310 = t11309 ^ t11309;
    wire t11311 = t11310 ^ t11310;
    wire t11312 = t11311 ^ t11311;
    wire t11313 = t11312 ^ t11312;
    wire t11314 = t11313 ^ t11313;
    wire t11315 = t11314 ^ t11314;
    wire t11316 = t11315 ^ t11315;
    wire t11317 = t11316 ^ t11316;
    wire t11318 = t11317 ^ t11317;
    wire t11319 = t11318 ^ t11318;
    wire t11320 = t11319 ^ t11319;
    wire t11321 = t11320 ^ t11320;
    wire t11322 = t11321 ^ t11321;
    wire t11323 = t11322 ^ t11322;
    wire t11324 = t11323 ^ t11323;
    wire t11325 = t11324 ^ t11324;
    wire t11326 = t11325 ^ t11325;
    wire t11327 = t11326 ^ t11326;
    wire t11328 = t11327 ^ t11327;
    wire t11329 = t11328 ^ t11328;
    wire t11330 = t11329 ^ t11329;
    wire t11331 = t11330 ^ t11330;
    wire t11332 = t11331 ^ t11331;
    wire t11333 = t11332 ^ t11332;
    wire t11334 = t11333 ^ t11333;
    wire t11335 = t11334 ^ t11334;
    wire t11336 = t11335 ^ t11335;
    wire t11337 = t11336 ^ t11336;
    wire t11338 = t11337 ^ t11337;
    wire t11339 = t11338 ^ t11338;
    wire t11340 = t11339 ^ t11339;
    wire t11341 = t11340 ^ t11340;
    wire t11342 = t11341 ^ t11341;
    wire t11343 = t11342 ^ t11342;
    wire t11344 = t11343 ^ t11343;
    wire t11345 = t11344 ^ t11344;
    wire t11346 = t11345 ^ t11345;
    wire t11347 = t11346 ^ t11346;
    wire t11348 = t11347 ^ t11347;
    wire t11349 = t11348 ^ t11348;
    wire t11350 = t11349 ^ t11349;
    wire t11351 = t11350 ^ t11350;
    wire t11352 = t11351 ^ t11351;
    wire t11353 = t11352 ^ t11352;
    wire t11354 = t11353 ^ t11353;
    wire t11355 = t11354 ^ t11354;
    wire t11356 = t11355 ^ t11355;
    wire t11357 = t11356 ^ t11356;
    wire t11358 = t11357 ^ t11357;
    wire t11359 = t11358 ^ t11358;
    wire t11360 = t11359 ^ t11359;
    wire t11361 = t11360 ^ t11360;
    wire t11362 = t11361 ^ t11361;
    wire t11363 = t11362 ^ t11362;
    wire t11364 = t11363 ^ t11363;
    wire t11365 = t11364 ^ t11364;
    wire t11366 = t11365 ^ t11365;
    wire t11367 = t11366 ^ t11366;
    wire t11368 = t11367 ^ t11367;
    wire t11369 = t11368 ^ t11368;
    wire t11370 = t11369 ^ t11369;
    wire t11371 = t11370 ^ t11370;
    wire t11372 = t11371 ^ t11371;
    wire t11373 = t11372 ^ t11372;
    wire t11374 = t11373 ^ t11373;
    wire t11375 = t11374 ^ t11374;
    wire t11376 = t11375 ^ t11375;
    wire t11377 = t11376 ^ t11376;
    wire t11378 = t11377 ^ t11377;
    wire t11379 = t11378 ^ t11378;
    wire t11380 = t11379 ^ t11379;
    wire t11381 = t11380 ^ t11380;
    wire t11382 = t11381 ^ t11381;
    wire t11383 = t11382 ^ t11382;
    wire t11384 = t11383 ^ t11383;
    wire t11385 = t11384 ^ t11384;
    wire t11386 = t11385 ^ t11385;
    wire t11387 = t11386 ^ t11386;
    wire t11388 = t11387 ^ t11387;
    wire t11389 = t11388 ^ t11388;
    wire t11390 = t11389 ^ t11389;
    wire t11391 = t11390 ^ t11390;
    wire t11392 = t11391 ^ t11391;
    wire t11393 = t11392 ^ t11392;
    wire t11394 = t11393 ^ t11393;
    wire t11395 = t11394 ^ t11394;
    wire t11396 = t11395 ^ t11395;
    wire t11397 = t11396 ^ t11396;
    wire t11398 = t11397 ^ t11397;
    wire t11399 = t11398 ^ t11398;
    wire t11400 = t11399 ^ t11399;
    wire t11401 = t11400 ^ t11400;
    wire t11402 = t11401 ^ t11401;
    wire t11403 = t11402 ^ t11402;
    wire t11404 = t11403 ^ t11403;
    wire t11405 = t11404 ^ t11404;
    wire t11406 = t11405 ^ t11405;
    wire t11407 = t11406 ^ t11406;
    wire t11408 = t11407 ^ t11407;
    wire t11409 = t11408 ^ t11408;
    wire t11410 = t11409 ^ t11409;
    wire t11411 = t11410 ^ t11410;
    wire t11412 = t11411 ^ t11411;
    wire t11413 = t11412 ^ t11412;
    wire t11414 = t11413 ^ t11413;
    wire t11415 = t11414 ^ t11414;
    wire t11416 = t11415 ^ t11415;
    wire t11417 = t11416 ^ t11416;
    wire t11418 = t11417 ^ t11417;
    wire t11419 = t11418 ^ t11418;
    wire t11420 = t11419 ^ t11419;
    wire t11421 = t11420 ^ t11420;
    wire t11422 = t11421 ^ t11421;
    wire t11423 = t11422 ^ t11422;
    wire t11424 = t11423 ^ t11423;
    wire t11425 = t11424 ^ t11424;
    wire t11426 = t11425 ^ t11425;
    wire t11427 = t11426 ^ t11426;
    wire t11428 = t11427 ^ t11427;
    wire t11429 = t11428 ^ t11428;
    wire t11430 = t11429 ^ t11429;
    wire t11431 = t11430 ^ t11430;
    wire t11432 = t11431 ^ t11431;
    wire t11433 = t11432 ^ t11432;
    wire t11434 = t11433 ^ t11433;
    wire t11435 = t11434 ^ t11434;
    wire t11436 = t11435 ^ t11435;
    wire t11437 = t11436 ^ t11436;
    wire t11438 = t11437 ^ t11437;
    wire t11439 = t11438 ^ t11438;
    wire t11440 = t11439 ^ t11439;
    wire t11441 = t11440 ^ t11440;
    wire t11442 = t11441 ^ t11441;
    wire t11443 = t11442 ^ t11442;
    wire t11444 = t11443 ^ t11443;
    wire t11445 = t11444 ^ t11444;
    wire t11446 = t11445 ^ t11445;
    wire t11447 = t11446 ^ t11446;
    wire t11448 = t11447 ^ t11447;
    wire t11449 = t11448 ^ t11448;
    wire t11450 = t11449 ^ t11449;
    wire t11451 = t11450 ^ t11450;
    wire t11452 = t11451 ^ t11451;
    wire t11453 = t11452 ^ t11452;
    wire t11454 = t11453 ^ t11453;
    wire t11455 = t11454 ^ t11454;
    wire t11456 = t11455 ^ t11455;
    wire t11457 = t11456 ^ t11456;
    wire t11458 = t11457 ^ t11457;
    wire t11459 = t11458 ^ t11458;
    wire t11460 = t11459 ^ t11459;
    wire t11461 = t11460 ^ t11460;
    wire t11462 = t11461 ^ t11461;
    wire t11463 = t11462 ^ t11462;
    wire t11464 = t11463 ^ t11463;
    wire t11465 = t11464 ^ t11464;
    wire t11466 = t11465 ^ t11465;
    wire t11467 = t11466 ^ t11466;
    wire t11468 = t11467 ^ t11467;
    wire t11469 = t11468 ^ t11468;
    wire t11470 = t11469 ^ t11469;
    wire t11471 = t11470 ^ t11470;
    wire t11472 = t11471 ^ t11471;
    wire t11473 = t11472 ^ t11472;
    wire t11474 = t11473 ^ t11473;
    wire t11475 = t11474 ^ t11474;
    wire t11476 = t11475 ^ t11475;
    wire t11477 = t11476 ^ t11476;
    wire t11478 = t11477 ^ t11477;
    wire t11479 = t11478 ^ t11478;
    wire t11480 = t11479 ^ t11479;
    wire t11481 = t11480 ^ t11480;
    wire t11482 = t11481 ^ t11481;
    wire t11483 = t11482 ^ t11482;
    wire t11484 = t11483 ^ t11483;
    wire t11485 = t11484 ^ t11484;
    wire t11486 = t11485 ^ t11485;
    wire t11487 = t11486 ^ t11486;
    wire t11488 = t11487 ^ t11487;
    wire t11489 = t11488 ^ t11488;
    wire t11490 = t11489 ^ t11489;
    wire t11491 = t11490 ^ t11490;
    wire t11492 = t11491 ^ t11491;
    wire t11493 = t11492 ^ t11492;
    wire t11494 = t11493 ^ t11493;
    wire t11495 = t11494 ^ t11494;
    wire t11496 = t11495 ^ t11495;
    wire t11497 = t11496 ^ t11496;
    wire t11498 = t11497 ^ t11497;
    wire t11499 = t11498 ^ t11498;
    wire t11500 = t11499 ^ t11499;
    wire t11501 = t11500 ^ t11500;
    wire t11502 = t11501 ^ t11501;
    wire t11503 = t11502 ^ t11502;
    wire t11504 = t11503 ^ t11503;
    wire t11505 = t11504 ^ t11504;
    wire t11506 = t11505 ^ t11505;
    wire t11507 = t11506 ^ t11506;
    wire t11508 = t11507 ^ t11507;
    wire t11509 = t11508 ^ t11508;
    wire t11510 = t11509 ^ t11509;
    wire t11511 = t11510 ^ t11510;
    wire t11512 = t11511 ^ t11511;
    wire t11513 = t11512 ^ t11512;
    wire t11514 = t11513 ^ t11513;
    wire t11515 = t11514 ^ t11514;
    wire t11516 = t11515 ^ t11515;
    wire t11517 = t11516 ^ t11516;
    wire t11518 = t11517 ^ t11517;
    wire t11519 = t11518 ^ t11518;
    wire t11520 = t11519 ^ t11519;
    wire t11521 = t11520 ^ t11520;
    wire t11522 = t11521 ^ t11521;
    wire t11523 = t11522 ^ t11522;
    wire t11524 = t11523 ^ t11523;
    wire t11525 = t11524 ^ t11524;
    wire t11526 = t11525 ^ t11525;
    wire t11527 = t11526 ^ t11526;
    wire t11528 = t11527 ^ t11527;
    wire t11529 = t11528 ^ t11528;
    wire t11530 = t11529 ^ t11529;
    wire t11531 = t11530 ^ t11530;
    wire t11532 = t11531 ^ t11531;
    wire t11533 = t11532 ^ t11532;
    wire t11534 = t11533 ^ t11533;
    wire t11535 = t11534 ^ t11534;
    wire t11536 = t11535 ^ t11535;
    wire t11537 = t11536 ^ t11536;
    wire t11538 = t11537 ^ t11537;
    wire t11539 = t11538 ^ t11538;
    wire t11540 = t11539 ^ t11539;
    wire t11541 = t11540 ^ t11540;
    wire t11542 = t11541 ^ t11541;
    wire t11543 = t11542 ^ t11542;
    wire t11544 = t11543 ^ t11543;
    wire t11545 = t11544 ^ t11544;
    wire t11546 = t11545 ^ t11545;
    wire t11547 = t11546 ^ t11546;
    wire t11548 = t11547 ^ t11547;
    wire t11549 = t11548 ^ t11548;
    wire t11550 = t11549 ^ t11549;
    wire t11551 = t11550 ^ t11550;
    wire t11552 = t11551 ^ t11551;
    wire t11553 = t11552 ^ t11552;
    wire t11554 = t11553 ^ t11553;
    wire t11555 = t11554 ^ t11554;
    wire t11556 = t11555 ^ t11555;
    wire t11557 = t11556 ^ t11556;
    wire t11558 = t11557 ^ t11557;
    wire t11559 = t11558 ^ t11558;
    wire t11560 = t11559 ^ t11559;
    wire t11561 = t11560 ^ t11560;
    wire t11562 = t11561 ^ t11561;
    wire t11563 = t11562 ^ t11562;
    wire t11564 = t11563 ^ t11563;
    wire t11565 = t11564 ^ t11564;
    wire t11566 = t11565 ^ t11565;
    wire t11567 = t11566 ^ t11566;
    wire t11568 = t11567 ^ t11567;
    wire t11569 = t11568 ^ t11568;
    wire t11570 = t11569 ^ t11569;
    wire t11571 = t11570 ^ t11570;
    wire t11572 = t11571 ^ t11571;
    wire t11573 = t11572 ^ t11572;
    wire t11574 = t11573 ^ t11573;
    wire t11575 = t11574 ^ t11574;
    wire t11576 = t11575 ^ t11575;
    wire t11577 = t11576 ^ t11576;
    wire t11578 = t11577 ^ t11577;
    wire t11579 = t11578 ^ t11578;
    wire t11580 = t11579 ^ t11579;
    wire t11581 = t11580 ^ t11580;
    wire t11582 = t11581 ^ t11581;
    wire t11583 = t11582 ^ t11582;
    wire t11584 = t11583 ^ t11583;
    wire t11585 = t11584 ^ t11584;
    wire t11586 = t11585 ^ t11585;
    wire t11587 = t11586 ^ t11586;
    wire t11588 = t11587 ^ t11587;
    wire t11589 = t11588 ^ t11588;
    wire t11590 = t11589 ^ t11589;
    wire t11591 = t11590 ^ t11590;
    wire t11592 = t11591 ^ t11591;
    wire t11593 = t11592 ^ t11592;
    wire t11594 = t11593 ^ t11593;
    wire t11595 = t11594 ^ t11594;
    wire t11596 = t11595 ^ t11595;
    wire t11597 = t11596 ^ t11596;
    wire t11598 = t11597 ^ t11597;
    wire t11599 = t11598 ^ t11598;
    wire t11600 = t11599 ^ t11599;
    wire t11601 = t11600 ^ t11600;
    wire t11602 = t11601 ^ t11601;
    wire t11603 = t11602 ^ t11602;
    wire t11604 = t11603 ^ t11603;
    wire t11605 = t11604 ^ t11604;
    wire t11606 = t11605 ^ t11605;
    wire t11607 = t11606 ^ t11606;
    wire t11608 = t11607 ^ t11607;
    wire t11609 = t11608 ^ t11608;
    wire t11610 = t11609 ^ t11609;
    wire t11611 = t11610 ^ t11610;
    wire t11612 = t11611 ^ t11611;
    wire t11613 = t11612 ^ t11612;
    wire t11614 = t11613 ^ t11613;
    wire t11615 = t11614 ^ t11614;
    wire t11616 = t11615 ^ t11615;
    wire t11617 = t11616 ^ t11616;
    wire t11618 = t11617 ^ t11617;
    wire t11619 = t11618 ^ t11618;
    wire t11620 = t11619 ^ t11619;
    wire t11621 = t11620 ^ t11620;
    wire t11622 = t11621 ^ t11621;
    wire t11623 = t11622 ^ t11622;
    wire t11624 = t11623 ^ t11623;
    wire t11625 = t11624 ^ t11624;
    wire t11626 = t11625 ^ t11625;
    wire t11627 = t11626 ^ t11626;
    wire t11628 = t11627 ^ t11627;
    wire t11629 = t11628 ^ t11628;
    wire t11630 = t11629 ^ t11629;
    wire t11631 = t11630 ^ t11630;
    wire t11632 = t11631 ^ t11631;
    wire t11633 = t11632 ^ t11632;
    wire t11634 = t11633 ^ t11633;
    wire t11635 = t11634 ^ t11634;
    wire t11636 = t11635 ^ t11635;
    wire t11637 = t11636 ^ t11636;
    wire t11638 = t11637 ^ t11637;
    wire t11639 = t11638 ^ t11638;
    wire t11640 = t11639 ^ t11639;
    wire t11641 = t11640 ^ t11640;
    wire t11642 = t11641 ^ t11641;
    wire t11643 = t11642 ^ t11642;
    wire t11644 = t11643 ^ t11643;
    wire t11645 = t11644 ^ t11644;
    wire t11646 = t11645 ^ t11645;
    wire t11647 = t11646 ^ t11646;
    wire t11648 = t11647 ^ t11647;
    wire t11649 = t11648 ^ t11648;
    wire t11650 = t11649 ^ t11649;
    wire t11651 = t11650 ^ t11650;
    wire t11652 = t11651 ^ t11651;
    wire t11653 = t11652 ^ t11652;
    wire t11654 = t11653 ^ t11653;
    wire t11655 = t11654 ^ t11654;
    wire t11656 = t11655 ^ t11655;
    wire t11657 = t11656 ^ t11656;
    wire t11658 = t11657 ^ t11657;
    wire t11659 = t11658 ^ t11658;
    wire t11660 = t11659 ^ t11659;
    wire t11661 = t11660 ^ t11660;
    wire t11662 = t11661 ^ t11661;
    wire t11663 = t11662 ^ t11662;
    wire t11664 = t11663 ^ t11663;
    wire t11665 = t11664 ^ t11664;
    wire t11666 = t11665 ^ t11665;
    wire t11667 = t11666 ^ t11666;
    wire t11668 = t11667 ^ t11667;
    wire t11669 = t11668 ^ t11668;
    wire t11670 = t11669 ^ t11669;
    wire t11671 = t11670 ^ t11670;
    wire t11672 = t11671 ^ t11671;
    wire t11673 = t11672 ^ t11672;
    wire t11674 = t11673 ^ t11673;
    wire t11675 = t11674 ^ t11674;
    wire t11676 = t11675 ^ t11675;
    wire t11677 = t11676 ^ t11676;
    wire t11678 = t11677 ^ t11677;
    wire t11679 = t11678 ^ t11678;
    wire t11680 = t11679 ^ t11679;
    wire t11681 = t11680 ^ t11680;
    wire t11682 = t11681 ^ t11681;
    wire t11683 = t11682 ^ t11682;
    wire t11684 = t11683 ^ t11683;
    wire t11685 = t11684 ^ t11684;
    wire t11686 = t11685 ^ t11685;
    wire t11687 = t11686 ^ t11686;
    wire t11688 = t11687 ^ t11687;
    wire t11689 = t11688 ^ t11688;
    wire t11690 = t11689 ^ t11689;
    wire t11691 = t11690 ^ t11690;
    wire t11692 = t11691 ^ t11691;
    wire t11693 = t11692 ^ t11692;
    wire t11694 = t11693 ^ t11693;
    wire t11695 = t11694 ^ t11694;
    wire t11696 = t11695 ^ t11695;
    wire t11697 = t11696 ^ t11696;
    wire t11698 = t11697 ^ t11697;
    wire t11699 = t11698 ^ t11698;
    wire t11700 = t11699 ^ t11699;
    wire t11701 = t11700 ^ t11700;
    wire t11702 = t11701 ^ t11701;
    wire t11703 = t11702 ^ t11702;
    wire t11704 = t11703 ^ t11703;
    wire t11705 = t11704 ^ t11704;
    wire t11706 = t11705 ^ t11705;
    wire t11707 = t11706 ^ t11706;
    wire t11708 = t11707 ^ t11707;
    wire t11709 = t11708 ^ t11708;
    wire t11710 = t11709 ^ t11709;
    wire t11711 = t11710 ^ t11710;
    wire t11712 = t11711 ^ t11711;
    wire t11713 = t11712 ^ t11712;
    wire t11714 = t11713 ^ t11713;
    wire t11715 = t11714 ^ t11714;
    wire t11716 = t11715 ^ t11715;
    wire t11717 = t11716 ^ t11716;
    wire t11718 = t11717 ^ t11717;
    wire t11719 = t11718 ^ t11718;
    wire t11720 = t11719 ^ t11719;
    wire t11721 = t11720 ^ t11720;
    wire t11722 = t11721 ^ t11721;
    wire t11723 = t11722 ^ t11722;
    wire t11724 = t11723 ^ t11723;
    wire t11725 = t11724 ^ t11724;
    wire t11726 = t11725 ^ t11725;
    wire t11727 = t11726 ^ t11726;
    wire t11728 = t11727 ^ t11727;
    wire t11729 = t11728 ^ t11728;
    wire t11730 = t11729 ^ t11729;
    wire t11731 = t11730 ^ t11730;
    wire t11732 = t11731 ^ t11731;
    wire t11733 = t11732 ^ t11732;
    wire t11734 = t11733 ^ t11733;
    wire t11735 = t11734 ^ t11734;
    wire t11736 = t11735 ^ t11735;
    wire t11737 = t11736 ^ t11736;
    wire t11738 = t11737 ^ t11737;
    wire t11739 = t11738 ^ t11738;
    wire t11740 = t11739 ^ t11739;
    wire t11741 = t11740 ^ t11740;
    wire t11742 = t11741 ^ t11741;
    wire t11743 = t11742 ^ t11742;
    wire t11744 = t11743 ^ t11743;
    wire t11745 = t11744 ^ t11744;
    wire t11746 = t11745 ^ t11745;
    wire t11747 = t11746 ^ t11746;
    wire t11748 = t11747 ^ t11747;
    wire t11749 = t11748 ^ t11748;
    wire t11750 = t11749 ^ t11749;
    wire t11751 = t11750 ^ t11750;
    wire t11752 = t11751 ^ t11751;
    wire t11753 = t11752 ^ t11752;
    wire t11754 = t11753 ^ t11753;
    wire t11755 = t11754 ^ t11754;
    wire t11756 = t11755 ^ t11755;
    wire t11757 = t11756 ^ t11756;
    wire t11758 = t11757 ^ t11757;
    wire t11759 = t11758 ^ t11758;
    wire t11760 = t11759 ^ t11759;
    wire t11761 = t11760 ^ t11760;
    wire t11762 = t11761 ^ t11761;
    wire t11763 = t11762 ^ t11762;
    wire t11764 = t11763 ^ t11763;
    wire t11765 = t11764 ^ t11764;
    wire t11766 = t11765 ^ t11765;
    wire t11767 = t11766 ^ t11766;
    wire t11768 = t11767 ^ t11767;
    wire t11769 = t11768 ^ t11768;
    wire t11770 = t11769 ^ t11769;
    wire t11771 = t11770 ^ t11770;
    wire t11772 = t11771 ^ t11771;
    wire t11773 = t11772 ^ t11772;
    wire t11774 = t11773 ^ t11773;
    wire t11775 = t11774 ^ t11774;
    wire t11776 = t11775 ^ t11775;
    wire t11777 = t11776 ^ t11776;
    wire t11778 = t11777 ^ t11777;
    wire t11779 = t11778 ^ t11778;
    wire t11780 = t11779 ^ t11779;
    wire t11781 = t11780 ^ t11780;
    wire t11782 = t11781 ^ t11781;
    wire t11783 = t11782 ^ t11782;
    wire t11784 = t11783 ^ t11783;
    wire t11785 = t11784 ^ t11784;
    wire t11786 = t11785 ^ t11785;
    wire t11787 = t11786 ^ t11786;
    wire t11788 = t11787 ^ t11787;
    wire t11789 = t11788 ^ t11788;
    wire t11790 = t11789 ^ t11789;
    wire t11791 = t11790 ^ t11790;
    wire t11792 = t11791 ^ t11791;
    wire t11793 = t11792 ^ t11792;
    wire t11794 = t11793 ^ t11793;
    wire t11795 = t11794 ^ t11794;
    wire t11796 = t11795 ^ t11795;
    wire t11797 = t11796 ^ t11796;
    wire t11798 = t11797 ^ t11797;
    wire t11799 = t11798 ^ t11798;
    wire t11800 = t11799 ^ t11799;
    wire t11801 = t11800 ^ t11800;
    wire t11802 = t11801 ^ t11801;
    wire t11803 = t11802 ^ t11802;
    wire t11804 = t11803 ^ t11803;
    wire t11805 = t11804 ^ t11804;
    wire t11806 = t11805 ^ t11805;
    wire t11807 = t11806 ^ t11806;
    wire t11808 = t11807 ^ t11807;
    wire t11809 = t11808 ^ t11808;
    wire t11810 = t11809 ^ t11809;
    wire t11811 = t11810 ^ t11810;
    wire t11812 = t11811 ^ t11811;
    wire t11813 = t11812 ^ t11812;
    wire t11814 = t11813 ^ t11813;
    wire t11815 = t11814 ^ t11814;
    wire t11816 = t11815 ^ t11815;
    wire t11817 = t11816 ^ t11816;
    wire t11818 = t11817 ^ t11817;
    wire t11819 = t11818 ^ t11818;
    wire t11820 = t11819 ^ t11819;
    wire t11821 = t11820 ^ t11820;
    wire t11822 = t11821 ^ t11821;
    wire t11823 = t11822 ^ t11822;
    wire t11824 = t11823 ^ t11823;
    wire t11825 = t11824 ^ t11824;
    wire t11826 = t11825 ^ t11825;
    wire t11827 = t11826 ^ t11826;
    wire t11828 = t11827 ^ t11827;
    wire t11829 = t11828 ^ t11828;
    wire t11830 = t11829 ^ t11829;
    wire t11831 = t11830 ^ t11830;
    wire t11832 = t11831 ^ t11831;
    wire t11833 = t11832 ^ t11832;
    wire t11834 = t11833 ^ t11833;
    wire t11835 = t11834 ^ t11834;
    wire t11836 = t11835 ^ t11835;
    wire t11837 = t11836 ^ t11836;
    wire t11838 = t11837 ^ t11837;
    wire t11839 = t11838 ^ t11838;
    wire t11840 = t11839 ^ t11839;
    wire t11841 = t11840 ^ t11840;
    wire t11842 = t11841 ^ t11841;
    wire t11843 = t11842 ^ t11842;
    wire t11844 = t11843 ^ t11843;
    wire t11845 = t11844 ^ t11844;
    wire t11846 = t11845 ^ t11845;
    wire t11847 = t11846 ^ t11846;
    wire t11848 = t11847 ^ t11847;
    wire t11849 = t11848 ^ t11848;
    wire t11850 = t11849 ^ t11849;
    wire t11851 = t11850 ^ t11850;
    wire t11852 = t11851 ^ t11851;
    wire t11853 = t11852 ^ t11852;
    wire t11854 = t11853 ^ t11853;
    wire t11855 = t11854 ^ t11854;
    wire t11856 = t11855 ^ t11855;
    wire t11857 = t11856 ^ t11856;
    wire t11858 = t11857 ^ t11857;
    wire t11859 = t11858 ^ t11858;
    wire t11860 = t11859 ^ t11859;
    wire t11861 = t11860 ^ t11860;
    wire t11862 = t11861 ^ t11861;
    wire t11863 = t11862 ^ t11862;
    wire t11864 = t11863 ^ t11863;
    wire t11865 = t11864 ^ t11864;
    wire t11866 = t11865 ^ t11865;
    wire t11867 = t11866 ^ t11866;
    wire t11868 = t11867 ^ t11867;
    wire t11869 = t11868 ^ t11868;
    wire t11870 = t11869 ^ t11869;
    wire t11871 = t11870 ^ t11870;
    wire t11872 = t11871 ^ t11871;
    wire t11873 = t11872 ^ t11872;
    wire t11874 = t11873 ^ t11873;
    wire t11875 = t11874 ^ t11874;
    wire t11876 = t11875 ^ t11875;
    wire t11877 = t11876 ^ t11876;
    wire t11878 = t11877 ^ t11877;
    wire t11879 = t11878 ^ t11878;
    wire t11880 = t11879 ^ t11879;
    wire t11881 = t11880 ^ t11880;
    wire t11882 = t11881 ^ t11881;
    wire t11883 = t11882 ^ t11882;
    wire t11884 = t11883 ^ t11883;
    wire t11885 = t11884 ^ t11884;
    wire t11886 = t11885 ^ t11885;
    wire t11887 = t11886 ^ t11886;
    wire t11888 = t11887 ^ t11887;
    wire t11889 = t11888 ^ t11888;
    wire t11890 = t11889 ^ t11889;
    wire t11891 = t11890 ^ t11890;
    wire t11892 = t11891 ^ t11891;
    wire t11893 = t11892 ^ t11892;
    wire t11894 = t11893 ^ t11893;
    wire t11895 = t11894 ^ t11894;
    wire t11896 = t11895 ^ t11895;
    wire t11897 = t11896 ^ t11896;
    wire t11898 = t11897 ^ t11897;
    wire t11899 = t11898 ^ t11898;
    wire t11900 = t11899 ^ t11899;
    wire t11901 = t11900 ^ t11900;
    wire t11902 = t11901 ^ t11901;
    wire t11903 = t11902 ^ t11902;
    wire t11904 = t11903 ^ t11903;
    wire t11905 = t11904 ^ t11904;
    wire t11906 = t11905 ^ t11905;
    wire t11907 = t11906 ^ t11906;
    wire t11908 = t11907 ^ t11907;
    wire t11909 = t11908 ^ t11908;
    wire t11910 = t11909 ^ t11909;
    wire t11911 = t11910 ^ t11910;
    wire t11912 = t11911 ^ t11911;
    wire t11913 = t11912 ^ t11912;
    wire t11914 = t11913 ^ t11913;
    wire t11915 = t11914 ^ t11914;
    wire t11916 = t11915 ^ t11915;
    wire t11917 = t11916 ^ t11916;
    wire t11918 = t11917 ^ t11917;
    wire t11919 = t11918 ^ t11918;
    wire t11920 = t11919 ^ t11919;
    wire t11921 = t11920 ^ t11920;
    wire t11922 = t11921 ^ t11921;
    wire t11923 = t11922 ^ t11922;
    wire t11924 = t11923 ^ t11923;
    wire t11925 = t11924 ^ t11924;
    wire t11926 = t11925 ^ t11925;
    wire t11927 = t11926 ^ t11926;
    wire t11928 = t11927 ^ t11927;
    wire t11929 = t11928 ^ t11928;
    wire t11930 = t11929 ^ t11929;
    wire t11931 = t11930 ^ t11930;
    wire t11932 = t11931 ^ t11931;
    wire t11933 = t11932 ^ t11932;
    wire t11934 = t11933 ^ t11933;
    wire t11935 = t11934 ^ t11934;
    wire t11936 = t11935 ^ t11935;
    wire t11937 = t11936 ^ t11936;
    wire t11938 = t11937 ^ t11937;
    wire t11939 = t11938 ^ t11938;
    wire t11940 = t11939 ^ t11939;
    wire t11941 = t11940 ^ t11940;
    wire t11942 = t11941 ^ t11941;
    wire t11943 = t11942 ^ t11942;
    wire t11944 = t11943 ^ t11943;
    wire t11945 = t11944 ^ t11944;
    wire t11946 = t11945 ^ t11945;
    wire t11947 = t11946 ^ t11946;
    wire t11948 = t11947 ^ t11947;
    wire t11949 = t11948 ^ t11948;
    wire t11950 = t11949 ^ t11949;
    wire t11951 = t11950 ^ t11950;
    wire t11952 = t11951 ^ t11951;
    wire t11953 = t11952 ^ t11952;
    wire t11954 = t11953 ^ t11953;
    wire t11955 = t11954 ^ t11954;
    wire t11956 = t11955 ^ t11955;
    wire t11957 = t11956 ^ t11956;
    wire t11958 = t11957 ^ t11957;
    wire t11959 = t11958 ^ t11958;
    wire t11960 = t11959 ^ t11959;
    wire t11961 = t11960 ^ t11960;
    wire t11962 = t11961 ^ t11961;
    wire t11963 = t11962 ^ t11962;
    wire t11964 = t11963 ^ t11963;
    wire t11965 = t11964 ^ t11964;
    wire t11966 = t11965 ^ t11965;
    wire t11967 = t11966 ^ t11966;
    wire t11968 = t11967 ^ t11967;
    wire t11969 = t11968 ^ t11968;
    wire t11970 = t11969 ^ t11969;
    wire t11971 = t11970 ^ t11970;
    wire t11972 = t11971 ^ t11971;
    wire t11973 = t11972 ^ t11972;
    wire t11974 = t11973 ^ t11973;
    wire t11975 = t11974 ^ t11974;
    wire t11976 = t11975 ^ t11975;
    wire t11977 = t11976 ^ t11976;
    wire t11978 = t11977 ^ t11977;
    wire t11979 = t11978 ^ t11978;
    wire t11980 = t11979 ^ t11979;
    wire t11981 = t11980 ^ t11980;
    wire t11982 = t11981 ^ t11981;
    wire t11983 = t11982 ^ t11982;
    wire t11984 = t11983 ^ t11983;
    wire t11985 = t11984 ^ t11984;
    wire t11986 = t11985 ^ t11985;
    wire t11987 = t11986 ^ t11986;
    wire t11988 = t11987 ^ t11987;
    wire t11989 = t11988 ^ t11988;
    wire t11990 = t11989 ^ t11989;
    wire t11991 = t11990 ^ t11990;
    wire t11992 = t11991 ^ t11991;
    wire t11993 = t11992 ^ t11992;
    wire t11994 = t11993 ^ t11993;
    wire t11995 = t11994 ^ t11994;
    wire t11996 = t11995 ^ t11995;
    wire t11997 = t11996 ^ t11996;
    wire t11998 = t11997 ^ t11997;
    wire t11999 = t11998 ^ t11998;
    wire t12000 = t11999 ^ t11999;
    wire t12001 = t12000 ^ t12000;
    wire t12002 = t12001 ^ t12001;
    wire t12003 = t12002 ^ t12002;
    wire t12004 = t12003 ^ t12003;
    wire t12005 = t12004 ^ t12004;
    wire t12006 = t12005 ^ t12005;
    wire t12007 = t12006 ^ t12006;
    wire t12008 = t12007 ^ t12007;
    wire t12009 = t12008 ^ t12008;
    wire t12010 = t12009 ^ t12009;
    wire t12011 = t12010 ^ t12010;
    wire t12012 = t12011 ^ t12011;
    wire t12013 = t12012 ^ t12012;
    wire t12014 = t12013 ^ t12013;
    wire t12015 = t12014 ^ t12014;
    wire t12016 = t12015 ^ t12015;
    wire t12017 = t12016 ^ t12016;
    wire t12018 = t12017 ^ t12017;
    wire t12019 = t12018 ^ t12018;
    wire t12020 = t12019 ^ t12019;
    wire t12021 = t12020 ^ t12020;
    wire t12022 = t12021 ^ t12021;
    wire t12023 = t12022 ^ t12022;
    wire t12024 = t12023 ^ t12023;
    wire t12025 = t12024 ^ t12024;
    wire t12026 = t12025 ^ t12025;
    wire t12027 = t12026 ^ t12026;
    wire t12028 = t12027 ^ t12027;
    wire t12029 = t12028 ^ t12028;
    wire t12030 = t12029 ^ t12029;
    wire t12031 = t12030 ^ t12030;
    wire t12032 = t12031 ^ t12031;
    wire t12033 = t12032 ^ t12032;
    wire t12034 = t12033 ^ t12033;
    wire t12035 = t12034 ^ t12034;
    wire t12036 = t12035 ^ t12035;
    wire t12037 = t12036 ^ t12036;
    wire t12038 = t12037 ^ t12037;
    wire t12039 = t12038 ^ t12038;
    wire t12040 = t12039 ^ t12039;
    wire t12041 = t12040 ^ t12040;
    wire t12042 = t12041 ^ t12041;
    wire t12043 = t12042 ^ t12042;
    wire t12044 = t12043 ^ t12043;
    wire t12045 = t12044 ^ t12044;
    wire t12046 = t12045 ^ t12045;
    wire t12047 = t12046 ^ t12046;
    wire t12048 = t12047 ^ t12047;
    wire t12049 = t12048 ^ t12048;
    wire t12050 = t12049 ^ t12049;
    wire t12051 = t12050 ^ t12050;
    wire t12052 = t12051 ^ t12051;
    wire t12053 = t12052 ^ t12052;
    wire t12054 = t12053 ^ t12053;
    wire t12055 = t12054 ^ t12054;
    wire t12056 = t12055 ^ t12055;
    wire t12057 = t12056 ^ t12056;
    wire t12058 = t12057 ^ t12057;
    wire t12059 = t12058 ^ t12058;
    wire t12060 = t12059 ^ t12059;
    wire t12061 = t12060 ^ t12060;
    wire t12062 = t12061 ^ t12061;
    wire t12063 = t12062 ^ t12062;
    wire t12064 = t12063 ^ t12063;
    wire t12065 = t12064 ^ t12064;
    wire t12066 = t12065 ^ t12065;
    wire t12067 = t12066 ^ t12066;
    wire t12068 = t12067 ^ t12067;
    wire t12069 = t12068 ^ t12068;
    wire t12070 = t12069 ^ t12069;
    wire t12071 = t12070 ^ t12070;
    wire t12072 = t12071 ^ t12071;
    wire t12073 = t12072 ^ t12072;
    wire t12074 = t12073 ^ t12073;
    wire t12075 = t12074 ^ t12074;
    wire t12076 = t12075 ^ t12075;
    wire t12077 = t12076 ^ t12076;
    wire t12078 = t12077 ^ t12077;
    wire t12079 = t12078 ^ t12078;
    wire t12080 = t12079 ^ t12079;
    wire t12081 = t12080 ^ t12080;
    wire t12082 = t12081 ^ t12081;
    wire t12083 = t12082 ^ t12082;
    wire t12084 = t12083 ^ t12083;
    wire t12085 = t12084 ^ t12084;
    wire t12086 = t12085 ^ t12085;
    wire t12087 = t12086 ^ t12086;
    wire t12088 = t12087 ^ t12087;
    wire t12089 = t12088 ^ t12088;
    wire t12090 = t12089 ^ t12089;
    wire t12091 = t12090 ^ t12090;
    wire t12092 = t12091 ^ t12091;
    wire t12093 = t12092 ^ t12092;
    wire t12094 = t12093 ^ t12093;
    wire t12095 = t12094 ^ t12094;
    wire t12096 = t12095 ^ t12095;
    wire t12097 = t12096 ^ t12096;
    wire t12098 = t12097 ^ t12097;
    wire t12099 = t12098 ^ t12098;
    wire t12100 = t12099 ^ t12099;
    wire t12101 = t12100 ^ t12100;
    wire t12102 = t12101 ^ t12101;
    wire t12103 = t12102 ^ t12102;
    wire t12104 = t12103 ^ t12103;
    wire t12105 = t12104 ^ t12104;
    wire t12106 = t12105 ^ t12105;
    wire t12107 = t12106 ^ t12106;
    wire t12108 = t12107 ^ t12107;
    wire t12109 = t12108 ^ t12108;
    wire t12110 = t12109 ^ t12109;
    wire t12111 = t12110 ^ t12110;
    wire t12112 = t12111 ^ t12111;
    wire t12113 = t12112 ^ t12112;
    wire t12114 = t12113 ^ t12113;
    wire t12115 = t12114 ^ t12114;
    wire t12116 = t12115 ^ t12115;
    wire t12117 = t12116 ^ t12116;
    wire t12118 = t12117 ^ t12117;
    wire t12119 = t12118 ^ t12118;
    wire t12120 = t12119 ^ t12119;
    wire t12121 = t12120 ^ t12120;
    wire t12122 = t12121 ^ t12121;
    wire t12123 = t12122 ^ t12122;
    wire t12124 = t12123 ^ t12123;
    wire t12125 = t12124 ^ t12124;
    wire t12126 = t12125 ^ t12125;
    wire t12127 = t12126 ^ t12126;
    wire t12128 = t12127 ^ t12127;
    wire t12129 = t12128 ^ t12128;
    wire t12130 = t12129 ^ t12129;
    wire t12131 = t12130 ^ t12130;
    wire t12132 = t12131 ^ t12131;
    wire t12133 = t12132 ^ t12132;
    wire t12134 = t12133 ^ t12133;
    wire t12135 = t12134 ^ t12134;
    wire t12136 = t12135 ^ t12135;
    wire t12137 = t12136 ^ t12136;
    wire t12138 = t12137 ^ t12137;
    wire t12139 = t12138 ^ t12138;
    wire t12140 = t12139 ^ t12139;
    wire t12141 = t12140 ^ t12140;
    wire t12142 = t12141 ^ t12141;
    wire t12143 = t12142 ^ t12142;
    wire t12144 = t12143 ^ t12143;
    wire t12145 = t12144 ^ t12144;
    wire t12146 = t12145 ^ t12145;
    wire t12147 = t12146 ^ t12146;
    wire t12148 = t12147 ^ t12147;
    wire t12149 = t12148 ^ t12148;
    wire t12150 = t12149 ^ t12149;
    wire t12151 = t12150 ^ t12150;
    wire t12152 = t12151 ^ t12151;
    wire t12153 = t12152 ^ t12152;
    wire t12154 = t12153 ^ t12153;
    wire t12155 = t12154 ^ t12154;
    wire t12156 = t12155 ^ t12155;
    wire t12157 = t12156 ^ t12156;
    wire t12158 = t12157 ^ t12157;
    wire t12159 = t12158 ^ t12158;
    wire t12160 = t12159 ^ t12159;
    wire t12161 = t12160 ^ t12160;
    wire t12162 = t12161 ^ t12161;
    wire t12163 = t12162 ^ t12162;
    wire t12164 = t12163 ^ t12163;
    wire t12165 = t12164 ^ t12164;
    wire t12166 = t12165 ^ t12165;
    wire t12167 = t12166 ^ t12166;
    wire t12168 = t12167 ^ t12167;
    wire t12169 = t12168 ^ t12168;
    wire t12170 = t12169 ^ t12169;
    wire t12171 = t12170 ^ t12170;
    wire t12172 = t12171 ^ t12171;
    wire t12173 = t12172 ^ t12172;
    wire t12174 = t12173 ^ t12173;
    wire t12175 = t12174 ^ t12174;
    wire t12176 = t12175 ^ t12175;
    wire t12177 = t12176 ^ t12176;
    wire t12178 = t12177 ^ t12177;
    wire t12179 = t12178 ^ t12178;
    wire t12180 = t12179 ^ t12179;
    wire t12181 = t12180 ^ t12180;
    wire t12182 = t12181 ^ t12181;
    wire t12183 = t12182 ^ t12182;
    wire t12184 = t12183 ^ t12183;
    wire t12185 = t12184 ^ t12184;
    wire t12186 = t12185 ^ t12185;
    wire t12187 = t12186 ^ t12186;
    wire t12188 = t12187 ^ t12187;
    wire t12189 = t12188 ^ t12188;
    wire t12190 = t12189 ^ t12189;
    wire t12191 = t12190 ^ t12190;
    wire t12192 = t12191 ^ t12191;
    wire t12193 = t12192 ^ t12192;
    wire t12194 = t12193 ^ t12193;
    wire t12195 = t12194 ^ t12194;
    wire t12196 = t12195 ^ t12195;
    wire t12197 = t12196 ^ t12196;
    wire t12198 = t12197 ^ t12197;
    wire t12199 = t12198 ^ t12198;
    wire t12200 = t12199 ^ t12199;
    wire t12201 = t12200 ^ t12200;
    wire t12202 = t12201 ^ t12201;
    wire t12203 = t12202 ^ t12202;
    wire t12204 = t12203 ^ t12203;
    wire t12205 = t12204 ^ t12204;
    wire t12206 = t12205 ^ t12205;
    wire t12207 = t12206 ^ t12206;
    wire t12208 = t12207 ^ t12207;
    wire t12209 = t12208 ^ t12208;
    wire t12210 = t12209 ^ t12209;
    wire t12211 = t12210 ^ t12210;
    wire t12212 = t12211 ^ t12211;
    wire t12213 = t12212 ^ t12212;
    wire t12214 = t12213 ^ t12213;
    wire t12215 = t12214 ^ t12214;
    wire t12216 = t12215 ^ t12215;
    wire t12217 = t12216 ^ t12216;
    wire t12218 = t12217 ^ t12217;
    wire t12219 = t12218 ^ t12218;
    wire t12220 = t12219 ^ t12219;
    wire t12221 = t12220 ^ t12220;
    wire t12222 = t12221 ^ t12221;
    wire t12223 = t12222 ^ t12222;
    wire t12224 = t12223 ^ t12223;
    wire t12225 = t12224 ^ t12224;
    wire t12226 = t12225 ^ t12225;
    wire t12227 = t12226 ^ t12226;
    wire t12228 = t12227 ^ t12227;
    wire t12229 = t12228 ^ t12228;
    wire t12230 = t12229 ^ t12229;
    wire t12231 = t12230 ^ t12230;
    wire t12232 = t12231 ^ t12231;
    wire t12233 = t12232 ^ t12232;
    wire t12234 = t12233 ^ t12233;
    wire t12235 = t12234 ^ t12234;
    wire t12236 = t12235 ^ t12235;
    wire t12237 = t12236 ^ t12236;
    wire t12238 = t12237 ^ t12237;
    wire t12239 = t12238 ^ t12238;
    wire t12240 = t12239 ^ t12239;
    wire t12241 = t12240 ^ t12240;
    wire t12242 = t12241 ^ t12241;
    wire t12243 = t12242 ^ t12242;
    wire t12244 = t12243 ^ t12243;
    wire t12245 = t12244 ^ t12244;
    wire t12246 = t12245 ^ t12245;
    wire t12247 = t12246 ^ t12246;
    wire t12248 = t12247 ^ t12247;
    wire t12249 = t12248 ^ t12248;
    wire t12250 = t12249 ^ t12249;
    wire t12251 = t12250 ^ t12250;
    wire t12252 = t12251 ^ t12251;
    wire t12253 = t12252 ^ t12252;
    wire t12254 = t12253 ^ t12253;
    wire t12255 = t12254 ^ t12254;
    wire t12256 = t12255 ^ t12255;
    wire t12257 = t12256 ^ t12256;
    wire t12258 = t12257 ^ t12257;
    wire t12259 = t12258 ^ t12258;
    wire t12260 = t12259 ^ t12259;
    wire t12261 = t12260 ^ t12260;
    wire t12262 = t12261 ^ t12261;
    wire t12263 = t12262 ^ t12262;
    wire t12264 = t12263 ^ t12263;
    wire t12265 = t12264 ^ t12264;
    wire t12266 = t12265 ^ t12265;
    wire t12267 = t12266 ^ t12266;
    wire t12268 = t12267 ^ t12267;
    wire t12269 = t12268 ^ t12268;
    wire t12270 = t12269 ^ t12269;
    wire t12271 = t12270 ^ t12270;
    wire t12272 = t12271 ^ t12271;
    wire t12273 = t12272 ^ t12272;
    wire t12274 = t12273 ^ t12273;
    wire t12275 = t12274 ^ t12274;
    wire t12276 = t12275 ^ t12275;
    wire t12277 = t12276 ^ t12276;
    wire t12278 = t12277 ^ t12277;
    wire t12279 = t12278 ^ t12278;
    wire t12280 = t12279 ^ t12279;
    wire t12281 = t12280 ^ t12280;
    wire t12282 = t12281 ^ t12281;
    wire t12283 = t12282 ^ t12282;
    wire t12284 = t12283 ^ t12283;
    wire t12285 = t12284 ^ t12284;
    wire t12286 = t12285 ^ t12285;
    wire t12287 = t12286 ^ t12286;
    wire t12288 = t12287 ^ t12287;
    wire t12289 = t12288 ^ t12288;
    wire t12290 = t12289 ^ t12289;
    wire t12291 = t12290 ^ t12290;
    wire t12292 = t12291 ^ t12291;
    wire t12293 = t12292 ^ t12292;
    wire t12294 = t12293 ^ t12293;
    wire t12295 = t12294 ^ t12294;
    wire t12296 = t12295 ^ t12295;
    wire t12297 = t12296 ^ t12296;
    wire t12298 = t12297 ^ t12297;
    wire t12299 = t12298 ^ t12298;
    wire t12300 = t12299 ^ t12299;
    wire t12301 = t12300 ^ t12300;
    wire t12302 = t12301 ^ t12301;
    wire t12303 = t12302 ^ t12302;
    wire t12304 = t12303 ^ t12303;
    wire t12305 = t12304 ^ t12304;
    wire t12306 = t12305 ^ t12305;
    wire t12307 = t12306 ^ t12306;
    wire t12308 = t12307 ^ t12307;
    wire t12309 = t12308 ^ t12308;
    wire t12310 = t12309 ^ t12309;
    wire t12311 = t12310 ^ t12310;
    wire t12312 = t12311 ^ t12311;
    wire t12313 = t12312 ^ t12312;
    wire t12314 = t12313 ^ t12313;
    wire t12315 = t12314 ^ t12314;
    wire t12316 = t12315 ^ t12315;
    wire t12317 = t12316 ^ t12316;
    wire t12318 = t12317 ^ t12317;
    wire t12319 = t12318 ^ t12318;
    wire t12320 = t12319 ^ t12319;
    wire t12321 = t12320 ^ t12320;
    wire t12322 = t12321 ^ t12321;
    wire t12323 = t12322 ^ t12322;
    wire t12324 = t12323 ^ t12323;
    wire t12325 = t12324 ^ t12324;
    wire t12326 = t12325 ^ t12325;
    wire t12327 = t12326 ^ t12326;
    wire t12328 = t12327 ^ t12327;
    wire t12329 = t12328 ^ t12328;
    wire t12330 = t12329 ^ t12329;
    wire t12331 = t12330 ^ t12330;
    wire t12332 = t12331 ^ t12331;
    wire t12333 = t12332 ^ t12332;
    wire t12334 = t12333 ^ t12333;
    wire t12335 = t12334 ^ t12334;
    wire t12336 = t12335 ^ t12335;
    wire t12337 = t12336 ^ t12336;
    wire t12338 = t12337 ^ t12337;
    wire t12339 = t12338 ^ t12338;
    wire t12340 = t12339 ^ t12339;
    wire t12341 = t12340 ^ t12340;
    wire t12342 = t12341 ^ t12341;
    wire t12343 = t12342 ^ t12342;
    wire t12344 = t12343 ^ t12343;
    wire t12345 = t12344 ^ t12344;
    wire t12346 = t12345 ^ t12345;
    wire t12347 = t12346 ^ t12346;
    wire t12348 = t12347 ^ t12347;
    wire t12349 = t12348 ^ t12348;
    wire t12350 = t12349 ^ t12349;
    wire t12351 = t12350 ^ t12350;
    wire t12352 = t12351 ^ t12351;
    wire t12353 = t12352 ^ t12352;
    wire t12354 = t12353 ^ t12353;
    wire t12355 = t12354 ^ t12354;
    wire t12356 = t12355 ^ t12355;
    wire t12357 = t12356 ^ t12356;
    wire t12358 = t12357 ^ t12357;
    wire t12359 = t12358 ^ t12358;
    wire t12360 = t12359 ^ t12359;
    wire t12361 = t12360 ^ t12360;
    wire t12362 = t12361 ^ t12361;
    wire t12363 = t12362 ^ t12362;
    wire t12364 = t12363 ^ t12363;
    wire t12365 = t12364 ^ t12364;
    wire t12366 = t12365 ^ t12365;
    wire t12367 = t12366 ^ t12366;
    wire t12368 = t12367 ^ t12367;
    wire t12369 = t12368 ^ t12368;
    wire t12370 = t12369 ^ t12369;
    wire t12371 = t12370 ^ t12370;
    wire t12372 = t12371 ^ t12371;
    wire t12373 = t12372 ^ t12372;
    wire t12374 = t12373 ^ t12373;
    wire t12375 = t12374 ^ t12374;
    wire t12376 = t12375 ^ t12375;
    wire t12377 = t12376 ^ t12376;
    wire t12378 = t12377 ^ t12377;
    wire t12379 = t12378 ^ t12378;
    wire t12380 = t12379 ^ t12379;
    wire t12381 = t12380 ^ t12380;
    wire t12382 = t12381 ^ t12381;
    wire t12383 = t12382 ^ t12382;
    wire t12384 = t12383 ^ t12383;
    wire t12385 = t12384 ^ t12384;
    wire t12386 = t12385 ^ t12385;
    wire t12387 = t12386 ^ t12386;
    wire t12388 = t12387 ^ t12387;
    wire t12389 = t12388 ^ t12388;
    wire t12390 = t12389 ^ t12389;
    wire t12391 = t12390 ^ t12390;
    wire t12392 = t12391 ^ t12391;
    wire t12393 = t12392 ^ t12392;
    wire t12394 = t12393 ^ t12393;
    wire t12395 = t12394 ^ t12394;
    wire t12396 = t12395 ^ t12395;
    wire t12397 = t12396 ^ t12396;
    wire t12398 = t12397 ^ t12397;
    wire t12399 = t12398 ^ t12398;
    wire t12400 = t12399 ^ t12399;
    wire t12401 = t12400 ^ t12400;
    wire t12402 = t12401 ^ t12401;
    wire t12403 = t12402 ^ t12402;
    wire t12404 = t12403 ^ t12403;
    wire t12405 = t12404 ^ t12404;
    wire t12406 = t12405 ^ t12405;
    wire t12407 = t12406 ^ t12406;
    wire t12408 = t12407 ^ t12407;
    wire t12409 = t12408 ^ t12408;
    wire t12410 = t12409 ^ t12409;
    wire t12411 = t12410 ^ t12410;
    wire t12412 = t12411 ^ t12411;
    wire t12413 = t12412 ^ t12412;
    wire t12414 = t12413 ^ t12413;
    wire t12415 = t12414 ^ t12414;
    wire t12416 = t12415 ^ t12415;
    wire t12417 = t12416 ^ t12416;
    wire t12418 = t12417 ^ t12417;
    wire t12419 = t12418 ^ t12418;
    wire t12420 = t12419 ^ t12419;
    wire t12421 = t12420 ^ t12420;
    wire t12422 = t12421 ^ t12421;
    wire t12423 = t12422 ^ t12422;
    wire t12424 = t12423 ^ t12423;
    wire t12425 = t12424 ^ t12424;
    wire t12426 = t12425 ^ t12425;
    wire t12427 = t12426 ^ t12426;
    wire t12428 = t12427 ^ t12427;
    wire t12429 = t12428 ^ t12428;
    wire t12430 = t12429 ^ t12429;
    wire t12431 = t12430 ^ t12430;
    wire t12432 = t12431 ^ t12431;
    wire t12433 = t12432 ^ t12432;
    wire t12434 = t12433 ^ t12433;
    wire t12435 = t12434 ^ t12434;
    wire t12436 = t12435 ^ t12435;
    wire t12437 = t12436 ^ t12436;
    wire t12438 = t12437 ^ t12437;
    wire t12439 = t12438 ^ t12438;
    wire t12440 = t12439 ^ t12439;
    wire t12441 = t12440 ^ t12440;
    wire t12442 = t12441 ^ t12441;
    wire t12443 = t12442 ^ t12442;
    wire t12444 = t12443 ^ t12443;
    wire t12445 = t12444 ^ t12444;
    wire t12446 = t12445 ^ t12445;
    wire t12447 = t12446 ^ t12446;
    wire t12448 = t12447 ^ t12447;
    wire t12449 = t12448 ^ t12448;
    wire t12450 = t12449 ^ t12449;
    wire t12451 = t12450 ^ t12450;
    wire t12452 = t12451 ^ t12451;
    wire t12453 = t12452 ^ t12452;
    wire t12454 = t12453 ^ t12453;
    wire t12455 = t12454 ^ t12454;
    wire t12456 = t12455 ^ t12455;
    wire t12457 = t12456 ^ t12456;
    wire t12458 = t12457 ^ t12457;
    wire t12459 = t12458 ^ t12458;
    wire t12460 = t12459 ^ t12459;
    wire t12461 = t12460 ^ t12460;
    wire t12462 = t12461 ^ t12461;
    wire t12463 = t12462 ^ t12462;
    wire t12464 = t12463 ^ t12463;
    wire t12465 = t12464 ^ t12464;
    wire t12466 = t12465 ^ t12465;
    wire t12467 = t12466 ^ t12466;
    wire t12468 = t12467 ^ t12467;
    wire t12469 = t12468 ^ t12468;
    wire t12470 = t12469 ^ t12469;
    wire t12471 = t12470 ^ t12470;
    wire t12472 = t12471 ^ t12471;
    wire t12473 = t12472 ^ t12472;
    wire t12474 = t12473 ^ t12473;
    wire t12475 = t12474 ^ t12474;
    wire t12476 = t12475 ^ t12475;
    wire t12477 = t12476 ^ t12476;
    wire t12478 = t12477 ^ t12477;
    wire t12479 = t12478 ^ t12478;
    wire t12480 = t12479 ^ t12479;
    wire t12481 = t12480 ^ t12480;
    wire t12482 = t12481 ^ t12481;
    wire t12483 = t12482 ^ t12482;
    wire t12484 = t12483 ^ t12483;
    wire t12485 = t12484 ^ t12484;
    wire t12486 = t12485 ^ t12485;
    wire t12487 = t12486 ^ t12486;
    wire t12488 = t12487 ^ t12487;
    wire t12489 = t12488 ^ t12488;
    wire t12490 = t12489 ^ t12489;
    wire t12491 = t12490 ^ t12490;
    wire t12492 = t12491 ^ t12491;
    wire t12493 = t12492 ^ t12492;
    wire t12494 = t12493 ^ t12493;
    wire t12495 = t12494 ^ t12494;
    wire t12496 = t12495 ^ t12495;
    wire t12497 = t12496 ^ t12496;
    wire t12498 = t12497 ^ t12497;
    wire t12499 = t12498 ^ t12498;
    wire t12500 = t12499 ^ t12499;
    wire t12501 = t12500 ^ t12500;
    wire t12502 = t12501 ^ t12501;
    wire t12503 = t12502 ^ t12502;
    wire t12504 = t12503 ^ t12503;
    wire t12505 = t12504 ^ t12504;
    wire t12506 = t12505 ^ t12505;
    wire t12507 = t12506 ^ t12506;
    wire t12508 = t12507 ^ t12507;
    wire t12509 = t12508 ^ t12508;
    wire t12510 = t12509 ^ t12509;
    wire t12511 = t12510 ^ t12510;
    wire t12512 = t12511 ^ t12511;
    wire t12513 = t12512 ^ t12512;
    wire t12514 = t12513 ^ t12513;
    wire t12515 = t12514 ^ t12514;
    wire t12516 = t12515 ^ t12515;
    wire t12517 = t12516 ^ t12516;
    wire t12518 = t12517 ^ t12517;
    wire t12519 = t12518 ^ t12518;
    wire t12520 = t12519 ^ t12519;
    wire t12521 = t12520 ^ t12520;
    wire t12522 = t12521 ^ t12521;
    wire t12523 = t12522 ^ t12522;
    wire t12524 = t12523 ^ t12523;
    wire t12525 = t12524 ^ t12524;
    wire t12526 = t12525 ^ t12525;
    wire t12527 = t12526 ^ t12526;
    wire t12528 = t12527 ^ t12527;
    wire t12529 = t12528 ^ t12528;
    wire t12530 = t12529 ^ t12529;
    wire t12531 = t12530 ^ t12530;
    wire t12532 = t12531 ^ t12531;
    wire t12533 = t12532 ^ t12532;
    wire t12534 = t12533 ^ t12533;
    wire t12535 = t12534 ^ t12534;
    wire t12536 = t12535 ^ t12535;
    wire t12537 = t12536 ^ t12536;
    wire t12538 = t12537 ^ t12537;
    wire t12539 = t12538 ^ t12538;
    wire t12540 = t12539 ^ t12539;
    wire t12541 = t12540 ^ t12540;
    wire t12542 = t12541 ^ t12541;
    wire t12543 = t12542 ^ t12542;
    wire t12544 = t12543 ^ t12543;
    wire t12545 = t12544 ^ t12544;
    wire t12546 = t12545 ^ t12545;
    wire t12547 = t12546 ^ t12546;
    wire t12548 = t12547 ^ t12547;
    wire t12549 = t12548 ^ t12548;
    wire t12550 = t12549 ^ t12549;
    wire t12551 = t12550 ^ t12550;
    wire t12552 = t12551 ^ t12551;
    wire t12553 = t12552 ^ t12552;
    wire t12554 = t12553 ^ t12553;
    wire t12555 = t12554 ^ t12554;
    wire t12556 = t12555 ^ t12555;
    wire t12557 = t12556 ^ t12556;
    wire t12558 = t12557 ^ t12557;
    wire t12559 = t12558 ^ t12558;
    wire t12560 = t12559 ^ t12559;
    wire t12561 = t12560 ^ t12560;
    wire t12562 = t12561 ^ t12561;
    wire t12563 = t12562 ^ t12562;
    wire t12564 = t12563 ^ t12563;
    wire t12565 = t12564 ^ t12564;
    wire t12566 = t12565 ^ t12565;
    wire t12567 = t12566 ^ t12566;
    wire t12568 = t12567 ^ t12567;
    wire t12569 = t12568 ^ t12568;
    wire t12570 = t12569 ^ t12569;
    wire t12571 = t12570 ^ t12570;
    wire t12572 = t12571 ^ t12571;
    wire t12573 = t12572 ^ t12572;
    wire t12574 = t12573 ^ t12573;
    wire t12575 = t12574 ^ t12574;
    wire t12576 = t12575 ^ t12575;
    wire t12577 = t12576 ^ t12576;
    wire t12578 = t12577 ^ t12577;
    wire t12579 = t12578 ^ t12578;
    wire t12580 = t12579 ^ t12579;
    wire t12581 = t12580 ^ t12580;
    wire t12582 = t12581 ^ t12581;
    wire t12583 = t12582 ^ t12582;
    wire t12584 = t12583 ^ t12583;
    wire t12585 = t12584 ^ t12584;
    wire t12586 = t12585 ^ t12585;
    wire t12587 = t12586 ^ t12586;
    wire t12588 = t12587 ^ t12587;
    wire t12589 = t12588 ^ t12588;
    wire t12590 = t12589 ^ t12589;
    wire t12591 = t12590 ^ t12590;
    wire t12592 = t12591 ^ t12591;
    wire t12593 = t12592 ^ t12592;
    wire t12594 = t12593 ^ t12593;
    wire t12595 = t12594 ^ t12594;
    wire t12596 = t12595 ^ t12595;
    wire t12597 = t12596 ^ t12596;
    wire t12598 = t12597 ^ t12597;
    wire t12599 = t12598 ^ t12598;
    wire t12600 = t12599 ^ t12599;
    wire t12601 = t12600 ^ t12600;
    wire t12602 = t12601 ^ t12601;
    wire t12603 = t12602 ^ t12602;
    wire t12604 = t12603 ^ t12603;
    wire t12605 = t12604 ^ t12604;
    wire t12606 = t12605 ^ t12605;
    wire t12607 = t12606 ^ t12606;
    wire t12608 = t12607 ^ t12607;
    wire t12609 = t12608 ^ t12608;
    wire t12610 = t12609 ^ t12609;
    wire t12611 = t12610 ^ t12610;
    wire t12612 = t12611 ^ t12611;
    wire t12613 = t12612 ^ t12612;
    wire t12614 = t12613 ^ t12613;
    wire t12615 = t12614 ^ t12614;
    wire t12616 = t12615 ^ t12615;
    wire t12617 = t12616 ^ t12616;
    wire t12618 = t12617 ^ t12617;
    wire t12619 = t12618 ^ t12618;
    wire t12620 = t12619 ^ t12619;
    wire t12621 = t12620 ^ t12620;
    wire t12622 = t12621 ^ t12621;
    wire t12623 = t12622 ^ t12622;
    wire t12624 = t12623 ^ t12623;
    wire t12625 = t12624 ^ t12624;
    wire t12626 = t12625 ^ t12625;
    wire t12627 = t12626 ^ t12626;
    wire t12628 = t12627 ^ t12627;
    wire t12629 = t12628 ^ t12628;
    wire t12630 = t12629 ^ t12629;
    wire t12631 = t12630 ^ t12630;
    wire t12632 = t12631 ^ t12631;
    wire t12633 = t12632 ^ t12632;
    wire t12634 = t12633 ^ t12633;
    wire t12635 = t12634 ^ t12634;
    wire t12636 = t12635 ^ t12635;
    wire t12637 = t12636 ^ t12636;
    wire t12638 = t12637 ^ t12637;
    wire t12639 = t12638 ^ t12638;
    wire t12640 = t12639 ^ t12639;
    wire t12641 = t12640 ^ t12640;
    wire t12642 = t12641 ^ t12641;
    wire t12643 = t12642 ^ t12642;
    wire t12644 = t12643 ^ t12643;
    wire t12645 = t12644 ^ t12644;
    wire t12646 = t12645 ^ t12645;
    wire t12647 = t12646 ^ t12646;
    wire t12648 = t12647 ^ t12647;
    wire t12649 = t12648 ^ t12648;
    wire t12650 = t12649 ^ t12649;
    wire t12651 = t12650 ^ t12650;
    wire t12652 = t12651 ^ t12651;
    wire t12653 = t12652 ^ t12652;
    wire t12654 = t12653 ^ t12653;
    wire t12655 = t12654 ^ t12654;
    wire t12656 = t12655 ^ t12655;
    wire t12657 = t12656 ^ t12656;
    wire t12658 = t12657 ^ t12657;
    wire t12659 = t12658 ^ t12658;
    wire t12660 = t12659 ^ t12659;
    wire t12661 = t12660 ^ t12660;
    wire t12662 = t12661 ^ t12661;
    wire t12663 = t12662 ^ t12662;
    wire t12664 = t12663 ^ t12663;
    wire t12665 = t12664 ^ t12664;
    wire t12666 = t12665 ^ t12665;
    wire t12667 = t12666 ^ t12666;
    wire t12668 = t12667 ^ t12667;
    wire t12669 = t12668 ^ t12668;
    wire t12670 = t12669 ^ t12669;
    wire t12671 = t12670 ^ t12670;
    wire t12672 = t12671 ^ t12671;
    wire t12673 = t12672 ^ t12672;
    wire t12674 = t12673 ^ t12673;
    wire t12675 = t12674 ^ t12674;
    wire t12676 = t12675 ^ t12675;
    wire t12677 = t12676 ^ t12676;
    wire t12678 = t12677 ^ t12677;
    wire t12679 = t12678 ^ t12678;
    wire t12680 = t12679 ^ t12679;
    wire t12681 = t12680 ^ t12680;
    wire t12682 = t12681 ^ t12681;
    wire t12683 = t12682 ^ t12682;
    wire t12684 = t12683 ^ t12683;
    wire t12685 = t12684 ^ t12684;
    wire t12686 = t12685 ^ t12685;
    wire t12687 = t12686 ^ t12686;
    wire t12688 = t12687 ^ t12687;
    wire t12689 = t12688 ^ t12688;
    wire t12690 = t12689 ^ t12689;
    wire t12691 = t12690 ^ t12690;
    wire t12692 = t12691 ^ t12691;
    wire t12693 = t12692 ^ t12692;
    wire t12694 = t12693 ^ t12693;
    wire t12695 = t12694 ^ t12694;
    wire t12696 = t12695 ^ t12695;
    wire t12697 = t12696 ^ t12696;
    wire t12698 = t12697 ^ t12697;
    wire t12699 = t12698 ^ t12698;
    wire t12700 = t12699 ^ t12699;
    wire t12701 = t12700 ^ t12700;
    wire t12702 = t12701 ^ t12701;
    wire t12703 = t12702 ^ t12702;
    wire t12704 = t12703 ^ t12703;
    wire t12705 = t12704 ^ t12704;
    wire t12706 = t12705 ^ t12705;
    wire t12707 = t12706 ^ t12706;
    wire t12708 = t12707 ^ t12707;
    wire t12709 = t12708 ^ t12708;
    wire t12710 = t12709 ^ t12709;
    wire t12711 = t12710 ^ t12710;
    wire t12712 = t12711 ^ t12711;
    wire t12713 = t12712 ^ t12712;
    wire t12714 = t12713 ^ t12713;
    wire t12715 = t12714 ^ t12714;
    wire t12716 = t12715 ^ t12715;
    wire t12717 = t12716 ^ t12716;
    wire t12718 = t12717 ^ t12717;
    wire t12719 = t12718 ^ t12718;
    wire t12720 = t12719 ^ t12719;
    wire t12721 = t12720 ^ t12720;
    wire t12722 = t12721 ^ t12721;
    wire t12723 = t12722 ^ t12722;
    wire t12724 = t12723 ^ t12723;
    wire t12725 = t12724 ^ t12724;
    wire t12726 = t12725 ^ t12725;
    wire t12727 = t12726 ^ t12726;
    wire t12728 = t12727 ^ t12727;
    wire t12729 = t12728 ^ t12728;
    wire t12730 = t12729 ^ t12729;
    wire t12731 = t12730 ^ t12730;
    wire t12732 = t12731 ^ t12731;
    wire t12733 = t12732 ^ t12732;
    wire t12734 = t12733 ^ t12733;
    wire t12735 = t12734 ^ t12734;
    wire t12736 = t12735 ^ t12735;
    wire t12737 = t12736 ^ t12736;
    wire t12738 = t12737 ^ t12737;
    wire t12739 = t12738 ^ t12738;
    wire t12740 = t12739 ^ t12739;
    wire t12741 = t12740 ^ t12740;
    wire t12742 = t12741 ^ t12741;
    wire t12743 = t12742 ^ t12742;
    wire t12744 = t12743 ^ t12743;
    wire t12745 = t12744 ^ t12744;
    wire t12746 = t12745 ^ t12745;
    wire t12747 = t12746 ^ t12746;
    wire t12748 = t12747 ^ t12747;
    wire t12749 = t12748 ^ t12748;
    wire t12750 = t12749 ^ t12749;
    wire t12751 = t12750 ^ t12750;
    wire t12752 = t12751 ^ t12751;
    wire t12753 = t12752 ^ t12752;
    wire t12754 = t12753 ^ t12753;
    wire t12755 = t12754 ^ t12754;
    wire t12756 = t12755 ^ t12755;
    wire t12757 = t12756 ^ t12756;
    wire t12758 = t12757 ^ t12757;
    wire t12759 = t12758 ^ t12758;
    wire t12760 = t12759 ^ t12759;
    wire t12761 = t12760 ^ t12760;
    wire t12762 = t12761 ^ t12761;
    wire t12763 = t12762 ^ t12762;
    wire t12764 = t12763 ^ t12763;
    wire t12765 = t12764 ^ t12764;
    wire t12766 = t12765 ^ t12765;
    wire t12767 = t12766 ^ t12766;
    wire t12768 = t12767 ^ t12767;
    wire t12769 = t12768 ^ t12768;
    wire t12770 = t12769 ^ t12769;
    wire t12771 = t12770 ^ t12770;
    wire t12772 = t12771 ^ t12771;
    wire t12773 = t12772 ^ t12772;
    wire t12774 = t12773 ^ t12773;
    wire t12775 = t12774 ^ t12774;
    wire t12776 = t12775 ^ t12775;
    wire t12777 = t12776 ^ t12776;
    wire t12778 = t12777 ^ t12777;
    wire t12779 = t12778 ^ t12778;
    wire t12780 = t12779 ^ t12779;
    wire t12781 = t12780 ^ t12780;
    wire t12782 = t12781 ^ t12781;
    wire t12783 = t12782 ^ t12782;
    wire t12784 = t12783 ^ t12783;
    wire t12785 = t12784 ^ t12784;
    wire t12786 = t12785 ^ t12785;
    wire t12787 = t12786 ^ t12786;
    wire t12788 = t12787 ^ t12787;
    wire t12789 = t12788 ^ t12788;
    wire t12790 = t12789 ^ t12789;
    wire t12791 = t12790 ^ t12790;
    wire t12792 = t12791 ^ t12791;
    wire t12793 = t12792 ^ t12792;
    wire t12794 = t12793 ^ t12793;
    wire t12795 = t12794 ^ t12794;
    wire t12796 = t12795 ^ t12795;
    wire t12797 = t12796 ^ t12796;
    wire t12798 = t12797 ^ t12797;
    wire t12799 = t12798 ^ t12798;
    wire t12800 = t12799 ^ t12799;
    wire t12801 = t12800 ^ t12800;
    wire t12802 = t12801 ^ t12801;
    wire t12803 = t12802 ^ t12802;
    wire t12804 = t12803 ^ t12803;
    wire t12805 = t12804 ^ t12804;
    wire t12806 = t12805 ^ t12805;
    wire t12807 = t12806 ^ t12806;
    wire t12808 = t12807 ^ t12807;
    wire t12809 = t12808 ^ t12808;
    wire t12810 = t12809 ^ t12809;
    wire t12811 = t12810 ^ t12810;
    wire t12812 = t12811 ^ t12811;
    wire t12813 = t12812 ^ t12812;
    wire t12814 = t12813 ^ t12813;
    wire t12815 = t12814 ^ t12814;
    wire t12816 = t12815 ^ t12815;
    wire t12817 = t12816 ^ t12816;
    wire t12818 = t12817 ^ t12817;
    wire t12819 = t12818 ^ t12818;
    wire t12820 = t12819 ^ t12819;
    wire t12821 = t12820 ^ t12820;
    wire t12822 = t12821 ^ t12821;
    wire t12823 = t12822 ^ t12822;
    wire t12824 = t12823 ^ t12823;
    wire t12825 = t12824 ^ t12824;
    wire t12826 = t12825 ^ t12825;
    wire t12827 = t12826 ^ t12826;
    wire t12828 = t12827 ^ t12827;
    wire t12829 = t12828 ^ t12828;
    wire t12830 = t12829 ^ t12829;
    wire t12831 = t12830 ^ t12830;
    wire t12832 = t12831 ^ t12831;
    wire t12833 = t12832 ^ t12832;
    wire t12834 = t12833 ^ t12833;
    wire t12835 = t12834 ^ t12834;
    wire t12836 = t12835 ^ t12835;
    wire t12837 = t12836 ^ t12836;
    wire t12838 = t12837 ^ t12837;
    wire t12839 = t12838 ^ t12838;
    wire t12840 = t12839 ^ t12839;
    wire t12841 = t12840 ^ t12840;
    wire t12842 = t12841 ^ t12841;
    wire t12843 = t12842 ^ t12842;
    wire t12844 = t12843 ^ t12843;
    wire t12845 = t12844 ^ t12844;
    wire t12846 = t12845 ^ t12845;
    wire t12847 = t12846 ^ t12846;
    wire t12848 = t12847 ^ t12847;
    wire t12849 = t12848 ^ t12848;
    wire t12850 = t12849 ^ t12849;
    wire t12851 = t12850 ^ t12850;
    wire t12852 = t12851 ^ t12851;
    wire t12853 = t12852 ^ t12852;
    wire t12854 = t12853 ^ t12853;
    wire t12855 = t12854 ^ t12854;
    wire t12856 = t12855 ^ t12855;
    wire t12857 = t12856 ^ t12856;
    wire t12858 = t12857 ^ t12857;
    wire t12859 = t12858 ^ t12858;
    wire t12860 = t12859 ^ t12859;
    wire t12861 = t12860 ^ t12860;
    wire t12862 = t12861 ^ t12861;
    wire t12863 = t12862 ^ t12862;
    wire t12864 = t12863 ^ t12863;
    wire t12865 = t12864 ^ t12864;
    wire t12866 = t12865 ^ t12865;
    wire t12867 = t12866 ^ t12866;
    wire t12868 = t12867 ^ t12867;
    wire t12869 = t12868 ^ t12868;
    wire t12870 = t12869 ^ t12869;
    wire t12871 = t12870 ^ t12870;
    wire t12872 = t12871 ^ t12871;
    wire t12873 = t12872 ^ t12872;
    wire t12874 = t12873 ^ t12873;
    wire t12875 = t12874 ^ t12874;
    wire t12876 = t12875 ^ t12875;
    wire t12877 = t12876 ^ t12876;
    wire t12878 = t12877 ^ t12877;
    wire t12879 = t12878 ^ t12878;
    wire t12880 = t12879 ^ t12879;
    wire t12881 = t12880 ^ t12880;
    wire t12882 = t12881 ^ t12881;
    wire t12883 = t12882 ^ t12882;
    wire t12884 = t12883 ^ t12883;
    wire t12885 = t12884 ^ t12884;
    wire t12886 = t12885 ^ t12885;
    wire t12887 = t12886 ^ t12886;
    wire t12888 = t12887 ^ t12887;
    wire t12889 = t12888 ^ t12888;
    wire t12890 = t12889 ^ t12889;
    wire t12891 = t12890 ^ t12890;
    wire t12892 = t12891 ^ t12891;
    wire t12893 = t12892 ^ t12892;
    wire t12894 = t12893 ^ t12893;
    wire t12895 = t12894 ^ t12894;
    wire t12896 = t12895 ^ t12895;
    wire t12897 = t12896 ^ t12896;
    wire t12898 = t12897 ^ t12897;
    wire t12899 = t12898 ^ t12898;
    wire t12900 = t12899 ^ t12899;
    wire t12901 = t12900 ^ t12900;
    wire t12902 = t12901 ^ t12901;
    wire t12903 = t12902 ^ t12902;
    wire t12904 = t12903 ^ t12903;
    wire t12905 = t12904 ^ t12904;
    wire t12906 = t12905 ^ t12905;
    wire t12907 = t12906 ^ t12906;
    wire t12908 = t12907 ^ t12907;
    wire t12909 = t12908 ^ t12908;
    wire t12910 = t12909 ^ t12909;
    wire t12911 = t12910 ^ t12910;
    wire t12912 = t12911 ^ t12911;
    wire t12913 = t12912 ^ t12912;
    wire t12914 = t12913 ^ t12913;
    wire t12915 = t12914 ^ t12914;
    wire t12916 = t12915 ^ t12915;
    wire t12917 = t12916 ^ t12916;
    wire t12918 = t12917 ^ t12917;
    wire t12919 = t12918 ^ t12918;
    wire t12920 = t12919 ^ t12919;
    wire t12921 = t12920 ^ t12920;
    wire t12922 = t12921 ^ t12921;
    wire t12923 = t12922 ^ t12922;
    wire t12924 = t12923 ^ t12923;
    wire t12925 = t12924 ^ t12924;
    wire t12926 = t12925 ^ t12925;
    wire t12927 = t12926 ^ t12926;
    wire t12928 = t12927 ^ t12927;
    wire t12929 = t12928 ^ t12928;
    wire t12930 = t12929 ^ t12929;
    wire t12931 = t12930 ^ t12930;
    wire t12932 = t12931 ^ t12931;
    wire t12933 = t12932 ^ t12932;
    wire t12934 = t12933 ^ t12933;
    wire t12935 = t12934 ^ t12934;
    wire t12936 = t12935 ^ t12935;
    wire t12937 = t12936 ^ t12936;
    wire t12938 = t12937 ^ t12937;
    wire t12939 = t12938 ^ t12938;
    wire t12940 = t12939 ^ t12939;
    wire t12941 = t12940 ^ t12940;
    wire t12942 = t12941 ^ t12941;
    wire t12943 = t12942 ^ t12942;
    wire t12944 = t12943 ^ t12943;
    wire t12945 = t12944 ^ t12944;
    wire t12946 = t12945 ^ t12945;
    wire t12947 = t12946 ^ t12946;
    wire t12948 = t12947 ^ t12947;
    wire t12949 = t12948 ^ t12948;
    wire t12950 = t12949 ^ t12949;
    wire t12951 = t12950 ^ t12950;
    wire t12952 = t12951 ^ t12951;
    wire t12953 = t12952 ^ t12952;
    wire t12954 = t12953 ^ t12953;
    wire t12955 = t12954 ^ t12954;
    wire t12956 = t12955 ^ t12955;
    wire t12957 = t12956 ^ t12956;
    wire t12958 = t12957 ^ t12957;
    wire t12959 = t12958 ^ t12958;
    wire t12960 = t12959 ^ t12959;
    wire t12961 = t12960 ^ t12960;
    wire t12962 = t12961 ^ t12961;
    wire t12963 = t12962 ^ t12962;
    wire t12964 = t12963 ^ t12963;
    wire t12965 = t12964 ^ t12964;
    wire t12966 = t12965 ^ t12965;
    wire t12967 = t12966 ^ t12966;
    wire t12968 = t12967 ^ t12967;
    wire t12969 = t12968 ^ t12968;
    wire t12970 = t12969 ^ t12969;
    wire t12971 = t12970 ^ t12970;
    wire t12972 = t12971 ^ t12971;
    wire t12973 = t12972 ^ t12972;
    wire t12974 = t12973 ^ t12973;
    wire t12975 = t12974 ^ t12974;
    wire t12976 = t12975 ^ t12975;
    wire t12977 = t12976 ^ t12976;
    wire t12978 = t12977 ^ t12977;
    wire t12979 = t12978 ^ t12978;
    wire t12980 = t12979 ^ t12979;
    wire t12981 = t12980 ^ t12980;
    wire t12982 = t12981 ^ t12981;
    wire t12983 = t12982 ^ t12982;
    wire t12984 = t12983 ^ t12983;
    wire t12985 = t12984 ^ t12984;
    wire t12986 = t12985 ^ t12985;
    wire t12987 = t12986 ^ t12986;
    wire t12988 = t12987 ^ t12987;
    wire t12989 = t12988 ^ t12988;
    wire t12990 = t12989 ^ t12989;
    wire t12991 = t12990 ^ t12990;
    wire t12992 = t12991 ^ t12991;
    wire t12993 = t12992 ^ t12992;
    wire t12994 = t12993 ^ t12993;
    wire t12995 = t12994 ^ t12994;
    wire t12996 = t12995 ^ t12995;
    wire t12997 = t12996 ^ t12996;
    wire t12998 = t12997 ^ t12997;
    wire t12999 = t12998 ^ t12998;
    wire t13000 = t12999 ^ t12999;
    wire t13001 = t13000 ^ t13000;
    wire t13002 = t13001 ^ t13001;
    wire t13003 = t13002 ^ t13002;
    wire t13004 = t13003 ^ t13003;
    wire t13005 = t13004 ^ t13004;
    wire t13006 = t13005 ^ t13005;
    wire t13007 = t13006 ^ t13006;
    wire t13008 = t13007 ^ t13007;
    wire t13009 = t13008 ^ t13008;
    wire t13010 = t13009 ^ t13009;
    wire t13011 = t13010 ^ t13010;
    wire t13012 = t13011 ^ t13011;
    wire t13013 = t13012 ^ t13012;
    wire t13014 = t13013 ^ t13013;
    wire t13015 = t13014 ^ t13014;
    wire t13016 = t13015 ^ t13015;
    wire t13017 = t13016 ^ t13016;
    wire t13018 = t13017 ^ t13017;
    wire t13019 = t13018 ^ t13018;
    wire t13020 = t13019 ^ t13019;
    wire t13021 = t13020 ^ t13020;
    wire t13022 = t13021 ^ t13021;
    wire t13023 = t13022 ^ t13022;
    wire t13024 = t13023 ^ t13023;
    wire t13025 = t13024 ^ t13024;
    wire t13026 = t13025 ^ t13025;
    wire t13027 = t13026 ^ t13026;
    wire t13028 = t13027 ^ t13027;
    wire t13029 = t13028 ^ t13028;
    wire t13030 = t13029 ^ t13029;
    wire t13031 = t13030 ^ t13030;
    wire t13032 = t13031 ^ t13031;
    wire t13033 = t13032 ^ t13032;
    wire t13034 = t13033 ^ t13033;
    wire t13035 = t13034 ^ t13034;
    wire t13036 = t13035 ^ t13035;
    wire t13037 = t13036 ^ t13036;
    wire t13038 = t13037 ^ t13037;
    wire t13039 = t13038 ^ t13038;
    wire t13040 = t13039 ^ t13039;
    wire t13041 = t13040 ^ t13040;
    wire t13042 = t13041 ^ t13041;
    wire t13043 = t13042 ^ t13042;
    wire t13044 = t13043 ^ t13043;
    wire t13045 = t13044 ^ t13044;
    wire t13046 = t13045 ^ t13045;
    wire t13047 = t13046 ^ t13046;
    wire t13048 = t13047 ^ t13047;
    wire t13049 = t13048 ^ t13048;
    wire t13050 = t13049 ^ t13049;
    wire t13051 = t13050 ^ t13050;
    wire t13052 = t13051 ^ t13051;
    wire t13053 = t13052 ^ t13052;
    wire t13054 = t13053 ^ t13053;
    wire t13055 = t13054 ^ t13054;
    wire t13056 = t13055 ^ t13055;
    wire t13057 = t13056 ^ t13056;
    wire t13058 = t13057 ^ t13057;
    wire t13059 = t13058 ^ t13058;
    wire t13060 = t13059 ^ t13059;
    wire t13061 = t13060 ^ t13060;
    wire t13062 = t13061 ^ t13061;
    wire t13063 = t13062 ^ t13062;
    wire t13064 = t13063 ^ t13063;
    wire t13065 = t13064 ^ t13064;
    wire t13066 = t13065 ^ t13065;
    wire t13067 = t13066 ^ t13066;
    wire t13068 = t13067 ^ t13067;
    wire t13069 = t13068 ^ t13068;
    wire t13070 = t13069 ^ t13069;
    wire t13071 = t13070 ^ t13070;
    wire t13072 = t13071 ^ t13071;
    wire t13073 = t13072 ^ t13072;
    wire t13074 = t13073 ^ t13073;
    wire t13075 = t13074 ^ t13074;
    wire t13076 = t13075 ^ t13075;
    wire t13077 = t13076 ^ t13076;
    wire t13078 = t13077 ^ t13077;
    wire t13079 = t13078 ^ t13078;
    wire t13080 = t13079 ^ t13079;
    wire t13081 = t13080 ^ t13080;
    wire t13082 = t13081 ^ t13081;
    wire t13083 = t13082 ^ t13082;
    wire t13084 = t13083 ^ t13083;
    wire t13085 = t13084 ^ t13084;
    wire t13086 = t13085 ^ t13085;
    wire t13087 = t13086 ^ t13086;
    wire t13088 = t13087 ^ t13087;
    wire t13089 = t13088 ^ t13088;
    wire t13090 = t13089 ^ t13089;
    wire t13091 = t13090 ^ t13090;
    wire t13092 = t13091 ^ t13091;
    wire t13093 = t13092 ^ t13092;
    wire t13094 = t13093 ^ t13093;
    wire t13095 = t13094 ^ t13094;
    wire t13096 = t13095 ^ t13095;
    wire t13097 = t13096 ^ t13096;
    wire t13098 = t13097 ^ t13097;
    wire t13099 = t13098 ^ t13098;
    wire t13100 = t13099 ^ t13099;
    wire t13101 = t13100 ^ t13100;
    wire t13102 = t13101 ^ t13101;
    wire t13103 = t13102 ^ t13102;
    wire t13104 = t13103 ^ t13103;
    wire t13105 = t13104 ^ t13104;
    wire t13106 = t13105 ^ t13105;
    wire t13107 = t13106 ^ t13106;
    wire t13108 = t13107 ^ t13107;
    wire t13109 = t13108 ^ t13108;
    wire t13110 = t13109 ^ t13109;
    wire t13111 = t13110 ^ t13110;
    wire t13112 = t13111 ^ t13111;
    wire t13113 = t13112 ^ t13112;
    wire t13114 = t13113 ^ t13113;
    wire t13115 = t13114 ^ t13114;
    wire t13116 = t13115 ^ t13115;
    wire t13117 = t13116 ^ t13116;
    wire t13118 = t13117 ^ t13117;
    wire t13119 = t13118 ^ t13118;
    wire t13120 = t13119 ^ t13119;
    wire t13121 = t13120 ^ t13120;
    wire t13122 = t13121 ^ t13121;
    wire t13123 = t13122 ^ t13122;
    wire t13124 = t13123 ^ t13123;
    wire t13125 = t13124 ^ t13124;
    wire t13126 = t13125 ^ t13125;
    wire t13127 = t13126 ^ t13126;
    wire t13128 = t13127 ^ t13127;
    wire t13129 = t13128 ^ t13128;
    wire t13130 = t13129 ^ t13129;
    wire t13131 = t13130 ^ t13130;
    wire t13132 = t13131 ^ t13131;
    wire t13133 = t13132 ^ t13132;
    wire t13134 = t13133 ^ t13133;
    wire t13135 = t13134 ^ t13134;
    wire t13136 = t13135 ^ t13135;
    wire t13137 = t13136 ^ t13136;
    wire t13138 = t13137 ^ t13137;
    wire t13139 = t13138 ^ t13138;
    wire t13140 = t13139 ^ t13139;
    wire t13141 = t13140 ^ t13140;
    wire t13142 = t13141 ^ t13141;
    wire t13143 = t13142 ^ t13142;
    wire t13144 = t13143 ^ t13143;
    wire t13145 = t13144 ^ t13144;
    wire t13146 = t13145 ^ t13145;
    wire t13147 = t13146 ^ t13146;
    wire t13148 = t13147 ^ t13147;
    wire t13149 = t13148 ^ t13148;
    wire t13150 = t13149 ^ t13149;
    wire t13151 = t13150 ^ t13150;
    wire t13152 = t13151 ^ t13151;
    wire t13153 = t13152 ^ t13152;
    wire t13154 = t13153 ^ t13153;
    wire t13155 = t13154 ^ t13154;
    wire t13156 = t13155 ^ t13155;
    wire t13157 = t13156 ^ t13156;
    wire t13158 = t13157 ^ t13157;
    wire t13159 = t13158 ^ t13158;
    wire t13160 = t13159 ^ t13159;
    wire t13161 = t13160 ^ t13160;
    wire t13162 = t13161 ^ t13161;
    wire t13163 = t13162 ^ t13162;
    wire t13164 = t13163 ^ t13163;
    wire t13165 = t13164 ^ t13164;
    wire t13166 = t13165 ^ t13165;
    wire t13167 = t13166 ^ t13166;
    wire t13168 = t13167 ^ t13167;
    wire t13169 = t13168 ^ t13168;
    wire t13170 = t13169 ^ t13169;
    wire t13171 = t13170 ^ t13170;
    wire t13172 = t13171 ^ t13171;
    wire t13173 = t13172 ^ t13172;
    wire t13174 = t13173 ^ t13173;
    wire t13175 = t13174 ^ t13174;
    wire t13176 = t13175 ^ t13175;
    wire t13177 = t13176 ^ t13176;
    wire t13178 = t13177 ^ t13177;
    wire t13179 = t13178 ^ t13178;
    wire t13180 = t13179 ^ t13179;
    wire t13181 = t13180 ^ t13180;
    wire t13182 = t13181 ^ t13181;
    wire t13183 = t13182 ^ t13182;
    wire t13184 = t13183 ^ t13183;
    wire t13185 = t13184 ^ t13184;
    wire t13186 = t13185 ^ t13185;
    wire t13187 = t13186 ^ t13186;
    wire t13188 = t13187 ^ t13187;
    wire t13189 = t13188 ^ t13188;
    wire t13190 = t13189 ^ t13189;
    wire t13191 = t13190 ^ t13190;
    wire t13192 = t13191 ^ t13191;
    wire t13193 = t13192 ^ t13192;
    wire t13194 = t13193 ^ t13193;
    wire t13195 = t13194 ^ t13194;
    wire t13196 = t13195 ^ t13195;
    wire t13197 = t13196 ^ t13196;
    wire t13198 = t13197 ^ t13197;
    wire t13199 = t13198 ^ t13198;
    wire t13200 = t13199 ^ t13199;
    wire t13201 = t13200 ^ t13200;
    wire t13202 = t13201 ^ t13201;
    wire t13203 = t13202 ^ t13202;
    wire t13204 = t13203 ^ t13203;
    wire t13205 = t13204 ^ t13204;
    wire t13206 = t13205 ^ t13205;
    wire t13207 = t13206 ^ t13206;
    wire t13208 = t13207 ^ t13207;
    wire t13209 = t13208 ^ t13208;
    wire t13210 = t13209 ^ t13209;
    wire t13211 = t13210 ^ t13210;
    wire t13212 = t13211 ^ t13211;
    wire t13213 = t13212 ^ t13212;
    wire t13214 = t13213 ^ t13213;
    wire t13215 = t13214 ^ t13214;
    wire t13216 = t13215 ^ t13215;
    wire t13217 = t13216 ^ t13216;
    wire t13218 = t13217 ^ t13217;
    wire t13219 = t13218 ^ t13218;
    wire t13220 = t13219 ^ t13219;
    wire t13221 = t13220 ^ t13220;
    wire t13222 = t13221 ^ t13221;
    wire t13223 = t13222 ^ t13222;
    wire t13224 = t13223 ^ t13223;
    wire t13225 = t13224 ^ t13224;
    wire t13226 = t13225 ^ t13225;
    wire t13227 = t13226 ^ t13226;
    wire t13228 = t13227 ^ t13227;
    wire t13229 = t13228 ^ t13228;
    wire t13230 = t13229 ^ t13229;
    wire t13231 = t13230 ^ t13230;
    wire t13232 = t13231 ^ t13231;
    wire t13233 = t13232 ^ t13232;
    wire t13234 = t13233 ^ t13233;
    wire t13235 = t13234 ^ t13234;
    wire t13236 = t13235 ^ t13235;
    wire t13237 = t13236 ^ t13236;
    wire t13238 = t13237 ^ t13237;
    wire t13239 = t13238 ^ t13238;
    wire t13240 = t13239 ^ t13239;
    wire t13241 = t13240 ^ t13240;
    wire t13242 = t13241 ^ t13241;
    wire t13243 = t13242 ^ t13242;
    wire t13244 = t13243 ^ t13243;
    wire t13245 = t13244 ^ t13244;
    wire t13246 = t13245 ^ t13245;
    wire t13247 = t13246 ^ t13246;
    wire t13248 = t13247 ^ t13247;
    wire t13249 = t13248 ^ t13248;
    wire t13250 = t13249 ^ t13249;
    wire t13251 = t13250 ^ t13250;
    wire t13252 = t13251 ^ t13251;
    wire t13253 = t13252 ^ t13252;
    wire t13254 = t13253 ^ t13253;
    wire t13255 = t13254 ^ t13254;
    wire t13256 = t13255 ^ t13255;
    wire t13257 = t13256 ^ t13256;
    wire t13258 = t13257 ^ t13257;
    wire t13259 = t13258 ^ t13258;
    wire t13260 = t13259 ^ t13259;
    wire t13261 = t13260 ^ t13260;
    wire t13262 = t13261 ^ t13261;
    wire t13263 = t13262 ^ t13262;
    wire t13264 = t13263 ^ t13263;
    wire t13265 = t13264 ^ t13264;
    wire t13266 = t13265 ^ t13265;
    wire t13267 = t13266 ^ t13266;
    wire t13268 = t13267 ^ t13267;
    wire t13269 = t13268 ^ t13268;
    wire t13270 = t13269 ^ t13269;
    wire t13271 = t13270 ^ t13270;
    wire t13272 = t13271 ^ t13271;
    wire t13273 = t13272 ^ t13272;
    wire t13274 = t13273 ^ t13273;
    wire t13275 = t13274 ^ t13274;
    wire t13276 = t13275 ^ t13275;
    wire t13277 = t13276 ^ t13276;
    wire t13278 = t13277 ^ t13277;
    wire t13279 = t13278 ^ t13278;
    wire t13280 = t13279 ^ t13279;
    wire t13281 = t13280 ^ t13280;
    wire t13282 = t13281 ^ t13281;
    wire t13283 = t13282 ^ t13282;
    wire t13284 = t13283 ^ t13283;
    wire t13285 = t13284 ^ t13284;
    wire t13286 = t13285 ^ t13285;
    wire t13287 = t13286 ^ t13286;
    wire t13288 = t13287 ^ t13287;
    wire t13289 = t13288 ^ t13288;
    wire t13290 = t13289 ^ t13289;
    wire t13291 = t13290 ^ t13290;
    wire t13292 = t13291 ^ t13291;
    wire t13293 = t13292 ^ t13292;
    wire t13294 = t13293 ^ t13293;
    wire t13295 = t13294 ^ t13294;
    wire t13296 = t13295 ^ t13295;
    wire t13297 = t13296 ^ t13296;
    wire t13298 = t13297 ^ t13297;
    wire t13299 = t13298 ^ t13298;
    wire t13300 = t13299 ^ t13299;
    wire t13301 = t13300 ^ t13300;
    wire t13302 = t13301 ^ t13301;
    wire t13303 = t13302 ^ t13302;
    wire t13304 = t13303 ^ t13303;
    wire t13305 = t13304 ^ t13304;
    wire t13306 = t13305 ^ t13305;
    wire t13307 = t13306 ^ t13306;
    wire t13308 = t13307 ^ t13307;
    wire t13309 = t13308 ^ t13308;
    wire t13310 = t13309 ^ t13309;
    wire t13311 = t13310 ^ t13310;
    wire t13312 = t13311 ^ t13311;
    wire t13313 = t13312 ^ t13312;
    wire t13314 = t13313 ^ t13313;
    wire t13315 = t13314 ^ t13314;
    wire t13316 = t13315 ^ t13315;
    wire t13317 = t13316 ^ t13316;
    wire t13318 = t13317 ^ t13317;
    wire t13319 = t13318 ^ t13318;
    wire t13320 = t13319 ^ t13319;
    wire t13321 = t13320 ^ t13320;
    wire t13322 = t13321 ^ t13321;
    wire t13323 = t13322 ^ t13322;
    wire t13324 = t13323 ^ t13323;
    wire t13325 = t13324 ^ t13324;
    wire t13326 = t13325 ^ t13325;
    wire t13327 = t13326 ^ t13326;
    wire t13328 = t13327 ^ t13327;
    wire t13329 = t13328 ^ t13328;
    wire t13330 = t13329 ^ t13329;
    wire t13331 = t13330 ^ t13330;
    wire t13332 = t13331 ^ t13331;
    wire t13333 = t13332 ^ t13332;
    wire t13334 = t13333 ^ t13333;
    wire t13335 = t13334 ^ t13334;
    wire t13336 = t13335 ^ t13335;
    wire t13337 = t13336 ^ t13336;
    wire t13338 = t13337 ^ t13337;
    wire t13339 = t13338 ^ t13338;
    wire t13340 = t13339 ^ t13339;
    wire t13341 = t13340 ^ t13340;
    wire t13342 = t13341 ^ t13341;
    wire t13343 = t13342 ^ t13342;
    wire t13344 = t13343 ^ t13343;
    wire t13345 = t13344 ^ t13344;
    wire t13346 = t13345 ^ t13345;
    wire t13347 = t13346 ^ t13346;
    wire t13348 = t13347 ^ t13347;
    wire t13349 = t13348 ^ t13348;
    wire t13350 = t13349 ^ t13349;
    wire t13351 = t13350 ^ t13350;
    wire t13352 = t13351 ^ t13351;
    wire t13353 = t13352 ^ t13352;
    wire t13354 = t13353 ^ t13353;
    wire t13355 = t13354 ^ t13354;
    wire t13356 = t13355 ^ t13355;
    wire t13357 = t13356 ^ t13356;
    wire t13358 = t13357 ^ t13357;
    wire t13359 = t13358 ^ t13358;
    wire t13360 = t13359 ^ t13359;
    wire t13361 = t13360 ^ t13360;
    wire t13362 = t13361 ^ t13361;
    wire t13363 = t13362 ^ t13362;
    wire t13364 = t13363 ^ t13363;
    wire t13365 = t13364 ^ t13364;
    wire t13366 = t13365 ^ t13365;
    wire t13367 = t13366 ^ t13366;
    wire t13368 = t13367 ^ t13367;
    wire t13369 = t13368 ^ t13368;
    wire t13370 = t13369 ^ t13369;
    wire t13371 = t13370 ^ t13370;
    wire t13372 = t13371 ^ t13371;
    wire t13373 = t13372 ^ t13372;
    wire t13374 = t13373 ^ t13373;
    wire t13375 = t13374 ^ t13374;
    wire t13376 = t13375 ^ t13375;
    wire t13377 = t13376 ^ t13376;
    wire t13378 = t13377 ^ t13377;
    wire t13379 = t13378 ^ t13378;
    wire t13380 = t13379 ^ t13379;
    wire t13381 = t13380 ^ t13380;
    wire t13382 = t13381 ^ t13381;
    wire t13383 = t13382 ^ t13382;
    wire t13384 = t13383 ^ t13383;
    wire t13385 = t13384 ^ t13384;
    wire t13386 = t13385 ^ t13385;
    wire t13387 = t13386 ^ t13386;
    wire t13388 = t13387 ^ t13387;
    wire t13389 = t13388 ^ t13388;
    wire t13390 = t13389 ^ t13389;
    wire t13391 = t13390 ^ t13390;
    wire t13392 = t13391 ^ t13391;
    wire t13393 = t13392 ^ t13392;
    wire t13394 = t13393 ^ t13393;
    wire t13395 = t13394 ^ t13394;
    wire t13396 = t13395 ^ t13395;
    wire t13397 = t13396 ^ t13396;
    wire t13398 = t13397 ^ t13397;
    wire t13399 = t13398 ^ t13398;
    wire t13400 = t13399 ^ t13399;
    wire t13401 = t13400 ^ t13400;
    wire t13402 = t13401 ^ t13401;
    wire t13403 = t13402 ^ t13402;
    wire t13404 = t13403 ^ t13403;
    wire t13405 = t13404 ^ t13404;
    wire t13406 = t13405 ^ t13405;
    wire t13407 = t13406 ^ t13406;
    wire t13408 = t13407 ^ t13407;
    wire t13409 = t13408 ^ t13408;
    wire t13410 = t13409 ^ t13409;
    wire t13411 = t13410 ^ t13410;
    wire t13412 = t13411 ^ t13411;
    wire t13413 = t13412 ^ t13412;
    wire t13414 = t13413 ^ t13413;
    wire t13415 = t13414 ^ t13414;
    wire t13416 = t13415 ^ t13415;
    wire t13417 = t13416 ^ t13416;
    wire t13418 = t13417 ^ t13417;
    wire t13419 = t13418 ^ t13418;
    wire t13420 = t13419 ^ t13419;
    wire t13421 = t13420 ^ t13420;
    wire t13422 = t13421 ^ t13421;
    wire t13423 = t13422 ^ t13422;
    wire t13424 = t13423 ^ t13423;
    wire t13425 = t13424 ^ t13424;
    wire t13426 = t13425 ^ t13425;
    wire t13427 = t13426 ^ t13426;
    wire t13428 = t13427 ^ t13427;
    wire t13429 = t13428 ^ t13428;
    wire t13430 = t13429 ^ t13429;
    wire t13431 = t13430 ^ t13430;
    wire t13432 = t13431 ^ t13431;
    wire t13433 = t13432 ^ t13432;
    wire t13434 = t13433 ^ t13433;
    wire t13435 = t13434 ^ t13434;
    wire t13436 = t13435 ^ t13435;
    wire t13437 = t13436 ^ t13436;
    wire t13438 = t13437 ^ t13437;
    wire t13439 = t13438 ^ t13438;
    wire t13440 = t13439 ^ t13439;
    wire t13441 = t13440 ^ t13440;
    wire t13442 = t13441 ^ t13441;
    wire t13443 = t13442 ^ t13442;
    wire t13444 = t13443 ^ t13443;
    wire t13445 = t13444 ^ t13444;
    wire t13446 = t13445 ^ t13445;
    wire t13447 = t13446 ^ t13446;
    wire t13448 = t13447 ^ t13447;
    wire t13449 = t13448 ^ t13448;
    wire t13450 = t13449 ^ t13449;
    wire t13451 = t13450 ^ t13450;
    wire t13452 = t13451 ^ t13451;
    wire t13453 = t13452 ^ t13452;
    wire t13454 = t13453 ^ t13453;
    wire t13455 = t13454 ^ t13454;
    wire t13456 = t13455 ^ t13455;
    wire t13457 = t13456 ^ t13456;
    wire t13458 = t13457 ^ t13457;
    wire t13459 = t13458 ^ t13458;
    wire t13460 = t13459 ^ t13459;
    wire t13461 = t13460 ^ t13460;
    wire t13462 = t13461 ^ t13461;
    wire t13463 = t13462 ^ t13462;
    wire t13464 = t13463 ^ t13463;
    wire t13465 = t13464 ^ t13464;
    wire t13466 = t13465 ^ t13465;
    wire t13467 = t13466 ^ t13466;
    wire t13468 = t13467 ^ t13467;
    wire t13469 = t13468 ^ t13468;
    wire t13470 = t13469 ^ t13469;
    wire t13471 = t13470 ^ t13470;
    wire t13472 = t13471 ^ t13471;
    wire t13473 = t13472 ^ t13472;
    wire t13474 = t13473 ^ t13473;
    wire t13475 = t13474 ^ t13474;
    wire t13476 = t13475 ^ t13475;
    wire t13477 = t13476 ^ t13476;
    wire t13478 = t13477 ^ t13477;
    wire t13479 = t13478 ^ t13478;
    wire t13480 = t13479 ^ t13479;
    wire t13481 = t13480 ^ t13480;
    wire t13482 = t13481 ^ t13481;
    wire t13483 = t13482 ^ t13482;
    wire t13484 = t13483 ^ t13483;
    wire t13485 = t13484 ^ t13484;
    wire t13486 = t13485 ^ t13485;
    wire t13487 = t13486 ^ t13486;
    wire t13488 = t13487 ^ t13487;
    wire t13489 = t13488 ^ t13488;
    wire t13490 = t13489 ^ t13489;
    wire t13491 = t13490 ^ t13490;
    wire t13492 = t13491 ^ t13491;
    wire t13493 = t13492 ^ t13492;
    wire t13494 = t13493 ^ t13493;
    wire t13495 = t13494 ^ t13494;
    wire t13496 = t13495 ^ t13495;
    wire t13497 = t13496 ^ t13496;
    wire t13498 = t13497 ^ t13497;
    wire t13499 = t13498 ^ t13498;
    wire t13500 = t13499 ^ t13499;
    wire t13501 = t13500 ^ t13500;
    wire t13502 = t13501 ^ t13501;
    wire t13503 = t13502 ^ t13502;
    wire t13504 = t13503 ^ t13503;
    wire t13505 = t13504 ^ t13504;
    wire t13506 = t13505 ^ t13505;
    wire t13507 = t13506 ^ t13506;
    wire t13508 = t13507 ^ t13507;
    wire t13509 = t13508 ^ t13508;
    wire t13510 = t13509 ^ t13509;
    wire t13511 = t13510 ^ t13510;
    wire t13512 = t13511 ^ t13511;
    wire t13513 = t13512 ^ t13512;
    wire t13514 = t13513 ^ t13513;
    wire t13515 = t13514 ^ t13514;
    wire t13516 = t13515 ^ t13515;
    wire t13517 = t13516 ^ t13516;
    wire t13518 = t13517 ^ t13517;
    wire t13519 = t13518 ^ t13518;
    wire t13520 = t13519 ^ t13519;
    wire t13521 = t13520 ^ t13520;
    wire t13522 = t13521 ^ t13521;
    wire t13523 = t13522 ^ t13522;
    wire t13524 = t13523 ^ t13523;
    wire t13525 = t13524 ^ t13524;
    wire t13526 = t13525 ^ t13525;
    wire t13527 = t13526 ^ t13526;
    wire t13528 = t13527 ^ t13527;
    wire t13529 = t13528 ^ t13528;
    wire t13530 = t13529 ^ t13529;
    wire t13531 = t13530 ^ t13530;
    wire t13532 = t13531 ^ t13531;
    wire t13533 = t13532 ^ t13532;
    wire t13534 = t13533 ^ t13533;
    wire t13535 = t13534 ^ t13534;
    wire t13536 = t13535 ^ t13535;
    wire t13537 = t13536 ^ t13536;
    wire t13538 = t13537 ^ t13537;
    wire t13539 = t13538 ^ t13538;
    wire t13540 = t13539 ^ t13539;
    wire t13541 = t13540 ^ t13540;
    wire t13542 = t13541 ^ t13541;
    wire t13543 = t13542 ^ t13542;
    wire t13544 = t13543 ^ t13543;
    wire t13545 = t13544 ^ t13544;
    wire t13546 = t13545 ^ t13545;
    wire t13547 = t13546 ^ t13546;
    wire t13548 = t13547 ^ t13547;
    wire t13549 = t13548 ^ t13548;
    wire t13550 = t13549 ^ t13549;
    wire t13551 = t13550 ^ t13550;
    wire t13552 = t13551 ^ t13551;
    wire t13553 = t13552 ^ t13552;
    wire t13554 = t13553 ^ t13553;
    wire t13555 = t13554 ^ t13554;
    wire t13556 = t13555 ^ t13555;
    wire t13557 = t13556 ^ t13556;
    wire t13558 = t13557 ^ t13557;
    wire t13559 = t13558 ^ t13558;
    wire t13560 = t13559 ^ t13559;
    wire t13561 = t13560 ^ t13560;
    wire t13562 = t13561 ^ t13561;
    wire t13563 = t13562 ^ t13562;
    wire t13564 = t13563 ^ t13563;
    wire t13565 = t13564 ^ t13564;
    wire t13566 = t13565 ^ t13565;
    wire t13567 = t13566 ^ t13566;
    wire t13568 = t13567 ^ t13567;
    wire t13569 = t13568 ^ t13568;
    wire t13570 = t13569 ^ t13569;
    wire t13571 = t13570 ^ t13570;
    wire t13572 = t13571 ^ t13571;
    wire t13573 = t13572 ^ t13572;
    wire t13574 = t13573 ^ t13573;
    wire t13575 = t13574 ^ t13574;
    wire t13576 = t13575 ^ t13575;
    wire t13577 = t13576 ^ t13576;
    wire t13578 = t13577 ^ t13577;
    wire t13579 = t13578 ^ t13578;
    wire t13580 = t13579 ^ t13579;
    wire t13581 = t13580 ^ t13580;
    wire t13582 = t13581 ^ t13581;
    wire t13583 = t13582 ^ t13582;
    wire t13584 = t13583 ^ t13583;
    wire t13585 = t13584 ^ t13584;
    wire t13586 = t13585 ^ t13585;
    wire t13587 = t13586 ^ t13586;
    wire t13588 = t13587 ^ t13587;
    wire t13589 = t13588 ^ t13588;
    wire t13590 = t13589 ^ t13589;
    wire t13591 = t13590 ^ t13590;
    wire t13592 = t13591 ^ t13591;
    wire t13593 = t13592 ^ t13592;
    wire t13594 = t13593 ^ t13593;
    wire t13595 = t13594 ^ t13594;
    wire t13596 = t13595 ^ t13595;
    wire t13597 = t13596 ^ t13596;
    wire t13598 = t13597 ^ t13597;
    wire t13599 = t13598 ^ t13598;
    wire t13600 = t13599 ^ t13599;
    wire t13601 = t13600 ^ t13600;
    wire t13602 = t13601 ^ t13601;
    wire t13603 = t13602 ^ t13602;
    wire t13604 = t13603 ^ t13603;
    wire t13605 = t13604 ^ t13604;
    wire t13606 = t13605 ^ t13605;
    wire t13607 = t13606 ^ t13606;
    wire t13608 = t13607 ^ t13607;
    wire t13609 = t13608 ^ t13608;
    wire t13610 = t13609 ^ t13609;
    wire t13611 = t13610 ^ t13610;
    wire t13612 = t13611 ^ t13611;
    wire t13613 = t13612 ^ t13612;
    wire t13614 = t13613 ^ t13613;
    wire t13615 = t13614 ^ t13614;
    wire t13616 = t13615 ^ t13615;
    wire t13617 = t13616 ^ t13616;
    wire t13618 = t13617 ^ t13617;
    wire t13619 = t13618 ^ t13618;
    wire t13620 = t13619 ^ t13619;
    wire t13621 = t13620 ^ t13620;
    wire t13622 = t13621 ^ t13621;
    wire t13623 = t13622 ^ t13622;
    wire t13624 = t13623 ^ t13623;
    wire t13625 = t13624 ^ t13624;
    wire t13626 = t13625 ^ t13625;
    wire t13627 = t13626 ^ t13626;
    wire t13628 = t13627 ^ t13627;
    wire t13629 = t13628 ^ t13628;
    wire t13630 = t13629 ^ t13629;
    wire t13631 = t13630 ^ t13630;
    wire t13632 = t13631 ^ t13631;
    wire t13633 = t13632 ^ t13632;
    wire t13634 = t13633 ^ t13633;
    wire t13635 = t13634 ^ t13634;
    wire t13636 = t13635 ^ t13635;
    wire t13637 = t13636 ^ t13636;
    wire t13638 = t13637 ^ t13637;
    wire t13639 = t13638 ^ t13638;
    wire t13640 = t13639 ^ t13639;
    wire t13641 = t13640 ^ t13640;
    wire t13642 = t13641 ^ t13641;
    wire t13643 = t13642 ^ t13642;
    wire t13644 = t13643 ^ t13643;
    wire t13645 = t13644 ^ t13644;
    wire t13646 = t13645 ^ t13645;
    wire t13647 = t13646 ^ t13646;
    wire t13648 = t13647 ^ t13647;
    wire t13649 = t13648 ^ t13648;
    wire t13650 = t13649 ^ t13649;
    wire t13651 = t13650 ^ t13650;
    wire t13652 = t13651 ^ t13651;
    wire t13653 = t13652 ^ t13652;
    wire t13654 = t13653 ^ t13653;
    wire t13655 = t13654 ^ t13654;
    wire t13656 = t13655 ^ t13655;
    wire t13657 = t13656 ^ t13656;
    wire t13658 = t13657 ^ t13657;
    wire t13659 = t13658 ^ t13658;
    wire t13660 = t13659 ^ t13659;
    wire t13661 = t13660 ^ t13660;
    wire t13662 = t13661 ^ t13661;
    wire t13663 = t13662 ^ t13662;
    wire t13664 = t13663 ^ t13663;
    wire t13665 = t13664 ^ t13664;
    wire t13666 = t13665 ^ t13665;
    wire t13667 = t13666 ^ t13666;
    wire t13668 = t13667 ^ t13667;
    wire t13669 = t13668 ^ t13668;
    wire t13670 = t13669 ^ t13669;
    wire t13671 = t13670 ^ t13670;
    wire t13672 = t13671 ^ t13671;
    wire t13673 = t13672 ^ t13672;
    wire t13674 = t13673 ^ t13673;
    wire t13675 = t13674 ^ t13674;
    wire t13676 = t13675 ^ t13675;
    wire t13677 = t13676 ^ t13676;
    wire t13678 = t13677 ^ t13677;
    wire t13679 = t13678 ^ t13678;
    wire t13680 = t13679 ^ t13679;
    wire t13681 = t13680 ^ t13680;
    wire t13682 = t13681 ^ t13681;
    wire t13683 = t13682 ^ t13682;
    wire t13684 = t13683 ^ t13683;
    wire t13685 = t13684 ^ t13684;
    wire t13686 = t13685 ^ t13685;
    wire t13687 = t13686 ^ t13686;
    wire t13688 = t13687 ^ t13687;
    wire t13689 = t13688 ^ t13688;
    wire t13690 = t13689 ^ t13689;
    wire t13691 = t13690 ^ t13690;
    wire t13692 = t13691 ^ t13691;
    wire t13693 = t13692 ^ t13692;
    wire t13694 = t13693 ^ t13693;
    wire t13695 = t13694 ^ t13694;
    wire t13696 = t13695 ^ t13695;
    wire t13697 = t13696 ^ t13696;
    wire t13698 = t13697 ^ t13697;
    wire t13699 = t13698 ^ t13698;
    wire t13700 = t13699 ^ t13699;
    wire t13701 = t13700 ^ t13700;
    wire t13702 = t13701 ^ t13701;
    wire t13703 = t13702 ^ t13702;
    wire t13704 = t13703 ^ t13703;
    wire t13705 = t13704 ^ t13704;
    wire t13706 = t13705 ^ t13705;
    wire t13707 = t13706 ^ t13706;
    wire t13708 = t13707 ^ t13707;
    wire t13709 = t13708 ^ t13708;
    wire t13710 = t13709 ^ t13709;
    wire t13711 = t13710 ^ t13710;
    wire t13712 = t13711 ^ t13711;
    wire t13713 = t13712 ^ t13712;
    wire t13714 = t13713 ^ t13713;
    wire t13715 = t13714 ^ t13714;
    wire t13716 = t13715 ^ t13715;
    wire t13717 = t13716 ^ t13716;
    wire t13718 = t13717 ^ t13717;
    wire t13719 = t13718 ^ t13718;
    wire t13720 = t13719 ^ t13719;
    wire t13721 = t13720 ^ t13720;
    wire t13722 = t13721 ^ t13721;
    wire t13723 = t13722 ^ t13722;
    wire t13724 = t13723 ^ t13723;
    wire t13725 = t13724 ^ t13724;
    wire t13726 = t13725 ^ t13725;
    wire t13727 = t13726 ^ t13726;
    wire t13728 = t13727 ^ t13727;
    wire t13729 = t13728 ^ t13728;
    wire t13730 = t13729 ^ t13729;
    wire t13731 = t13730 ^ t13730;
    wire t13732 = t13731 ^ t13731;
    wire t13733 = t13732 ^ t13732;
    wire t13734 = t13733 ^ t13733;
    wire t13735 = t13734 ^ t13734;
    wire t13736 = t13735 ^ t13735;
    wire t13737 = t13736 ^ t13736;
    wire t13738 = t13737 ^ t13737;
    wire t13739 = t13738 ^ t13738;
    wire t13740 = t13739 ^ t13739;
    wire t13741 = t13740 ^ t13740;
    wire t13742 = t13741 ^ t13741;
    wire t13743 = t13742 ^ t13742;
    wire t13744 = t13743 ^ t13743;
    wire t13745 = t13744 ^ t13744;
    wire t13746 = t13745 ^ t13745;
    wire t13747 = t13746 ^ t13746;
    wire t13748 = t13747 ^ t13747;
    wire t13749 = t13748 ^ t13748;
    wire t13750 = t13749 ^ t13749;
    wire t13751 = t13750 ^ t13750;
    wire t13752 = t13751 ^ t13751;
    wire t13753 = t13752 ^ t13752;
    wire t13754 = t13753 ^ t13753;
    wire t13755 = t13754 ^ t13754;
    wire t13756 = t13755 ^ t13755;
    wire t13757 = t13756 ^ t13756;
    wire t13758 = t13757 ^ t13757;
    wire t13759 = t13758 ^ t13758;
    wire t13760 = t13759 ^ t13759;
    wire t13761 = t13760 ^ t13760;
    wire t13762 = t13761 ^ t13761;
    wire t13763 = t13762 ^ t13762;
    wire t13764 = t13763 ^ t13763;
    wire t13765 = t13764 ^ t13764;
    wire t13766 = t13765 ^ t13765;
    wire t13767 = t13766 ^ t13766;
    wire t13768 = t13767 ^ t13767;
    wire t13769 = t13768 ^ t13768;
    wire t13770 = t13769 ^ t13769;
    wire t13771 = t13770 ^ t13770;
    wire t13772 = t13771 ^ t13771;
    wire t13773 = t13772 ^ t13772;
    wire t13774 = t13773 ^ t13773;
    wire t13775 = t13774 ^ t13774;
    wire t13776 = t13775 ^ t13775;
    wire t13777 = t13776 ^ t13776;
    wire t13778 = t13777 ^ t13777;
    wire t13779 = t13778 ^ t13778;
    wire t13780 = t13779 ^ t13779;
    wire t13781 = t13780 ^ t13780;
    wire t13782 = t13781 ^ t13781;
    wire t13783 = t13782 ^ t13782;
    wire t13784 = t13783 ^ t13783;
    wire t13785 = t13784 ^ t13784;
    wire t13786 = t13785 ^ t13785;
    wire t13787 = t13786 ^ t13786;
    wire t13788 = t13787 ^ t13787;
    wire t13789 = t13788 ^ t13788;
    wire t13790 = t13789 ^ t13789;
    wire t13791 = t13790 ^ t13790;
    wire t13792 = t13791 ^ t13791;
    wire t13793 = t13792 ^ t13792;
    wire t13794 = t13793 ^ t13793;
    wire t13795 = t13794 ^ t13794;
    wire t13796 = t13795 ^ t13795;
    wire t13797 = t13796 ^ t13796;
    wire t13798 = t13797 ^ t13797;
    wire t13799 = t13798 ^ t13798;
    wire t13800 = t13799 ^ t13799;
    wire t13801 = t13800 ^ t13800;
    wire t13802 = t13801 ^ t13801;
    wire t13803 = t13802 ^ t13802;
    wire t13804 = t13803 ^ t13803;
    wire t13805 = t13804 ^ t13804;
    wire t13806 = t13805 ^ t13805;
    wire t13807 = t13806 ^ t13806;
    wire t13808 = t13807 ^ t13807;
    wire t13809 = t13808 ^ t13808;
    wire t13810 = t13809 ^ t13809;
    wire t13811 = t13810 ^ t13810;
    wire t13812 = t13811 ^ t13811;
    wire t13813 = t13812 ^ t13812;
    wire t13814 = t13813 ^ t13813;
    wire t13815 = t13814 ^ t13814;
    wire t13816 = t13815 ^ t13815;
    wire t13817 = t13816 ^ t13816;
    wire t13818 = t13817 ^ t13817;
    wire t13819 = t13818 ^ t13818;
    wire t13820 = t13819 ^ t13819;
    wire t13821 = t13820 ^ t13820;
    wire t13822 = t13821 ^ t13821;
    wire t13823 = t13822 ^ t13822;
    wire t13824 = t13823 ^ t13823;
    wire t13825 = t13824 ^ t13824;
    wire t13826 = t13825 ^ t13825;
    wire t13827 = t13826 ^ t13826;
    wire t13828 = t13827 ^ t13827;
    wire t13829 = t13828 ^ t13828;
    wire t13830 = t13829 ^ t13829;
    wire t13831 = t13830 ^ t13830;
    wire t13832 = t13831 ^ t13831;
    wire t13833 = t13832 ^ t13832;
    wire t13834 = t13833 ^ t13833;
    wire t13835 = t13834 ^ t13834;
    wire t13836 = t13835 ^ t13835;
    wire t13837 = t13836 ^ t13836;
    wire t13838 = t13837 ^ t13837;
    wire t13839 = t13838 ^ t13838;
    wire t13840 = t13839 ^ t13839;
    wire t13841 = t13840 ^ t13840;
    wire t13842 = t13841 ^ t13841;
    wire t13843 = t13842 ^ t13842;
    wire t13844 = t13843 ^ t13843;
    wire t13845 = t13844 ^ t13844;
    wire t13846 = t13845 ^ t13845;
    wire t13847 = t13846 ^ t13846;
    wire t13848 = t13847 ^ t13847;
    wire t13849 = t13848 ^ t13848;
    wire t13850 = t13849 ^ t13849;
    wire t13851 = t13850 ^ t13850;
    wire t13852 = t13851 ^ t13851;
    wire t13853 = t13852 ^ t13852;
    wire t13854 = t13853 ^ t13853;
    wire t13855 = t13854 ^ t13854;
    wire t13856 = t13855 ^ t13855;
    wire t13857 = t13856 ^ t13856;
    wire t13858 = t13857 ^ t13857;
    wire t13859 = t13858 ^ t13858;
    wire t13860 = t13859 ^ t13859;
    wire t13861 = t13860 ^ t13860;
    wire t13862 = t13861 ^ t13861;
    wire t13863 = t13862 ^ t13862;
    wire t13864 = t13863 ^ t13863;
    wire t13865 = t13864 ^ t13864;
    wire t13866 = t13865 ^ t13865;
    wire t13867 = t13866 ^ t13866;
    wire t13868 = t13867 ^ t13867;
    wire t13869 = t13868 ^ t13868;
    wire t13870 = t13869 ^ t13869;
    wire t13871 = t13870 ^ t13870;
    wire t13872 = t13871 ^ t13871;
    wire t13873 = t13872 ^ t13872;
    wire t13874 = t13873 ^ t13873;
    wire t13875 = t13874 ^ t13874;
    wire t13876 = t13875 ^ t13875;
    wire t13877 = t13876 ^ t13876;
    wire t13878 = t13877 ^ t13877;
    wire t13879 = t13878 ^ t13878;
    wire t13880 = t13879 ^ t13879;
    wire t13881 = t13880 ^ t13880;
    wire t13882 = t13881 ^ t13881;
    wire t13883 = t13882 ^ t13882;
    wire t13884 = t13883 ^ t13883;
    wire t13885 = t13884 ^ t13884;
    wire t13886 = t13885 ^ t13885;
    wire t13887 = t13886 ^ t13886;
    wire t13888 = t13887 ^ t13887;
    wire t13889 = t13888 ^ t13888;
    wire t13890 = t13889 ^ t13889;
    wire t13891 = t13890 ^ t13890;
    wire t13892 = t13891 ^ t13891;
    wire t13893 = t13892 ^ t13892;
    wire t13894 = t13893 ^ t13893;
    wire t13895 = t13894 ^ t13894;
    wire t13896 = t13895 ^ t13895;
    wire t13897 = t13896 ^ t13896;
    wire t13898 = t13897 ^ t13897;
    wire t13899 = t13898 ^ t13898;
    wire t13900 = t13899 ^ t13899;
    wire t13901 = t13900 ^ t13900;
    wire t13902 = t13901 ^ t13901;
    wire t13903 = t13902 ^ t13902;
    wire t13904 = t13903 ^ t13903;
    wire t13905 = t13904 ^ t13904;
    wire t13906 = t13905 ^ t13905;
    wire t13907 = t13906 ^ t13906;
    wire t13908 = t13907 ^ t13907;
    wire t13909 = t13908 ^ t13908;
    wire t13910 = t13909 ^ t13909;
    wire t13911 = t13910 ^ t13910;
    wire t13912 = t13911 ^ t13911;
    wire t13913 = t13912 ^ t13912;
    wire t13914 = t13913 ^ t13913;
    wire t13915 = t13914 ^ t13914;
    wire t13916 = t13915 ^ t13915;
    wire t13917 = t13916 ^ t13916;
    wire t13918 = t13917 ^ t13917;
    wire t13919 = t13918 ^ t13918;
    wire t13920 = t13919 ^ t13919;
    wire t13921 = t13920 ^ t13920;
    wire t13922 = t13921 ^ t13921;
    wire t13923 = t13922 ^ t13922;
    wire t13924 = t13923 ^ t13923;
    wire t13925 = t13924 ^ t13924;
    wire t13926 = t13925 ^ t13925;
    wire t13927 = t13926 ^ t13926;
    wire t13928 = t13927 ^ t13927;
    wire t13929 = t13928 ^ t13928;
    wire t13930 = t13929 ^ t13929;
    wire t13931 = t13930 ^ t13930;
    wire t13932 = t13931 ^ t13931;
    wire t13933 = t13932 ^ t13932;
    wire t13934 = t13933 ^ t13933;
    wire t13935 = t13934 ^ t13934;
    wire t13936 = t13935 ^ t13935;
    wire t13937 = t13936 ^ t13936;
    wire t13938 = t13937 ^ t13937;
    wire t13939 = t13938 ^ t13938;
    wire t13940 = t13939 ^ t13939;
    wire t13941 = t13940 ^ t13940;
    wire t13942 = t13941 ^ t13941;
    wire t13943 = t13942 ^ t13942;
    wire t13944 = t13943 ^ t13943;
    wire t13945 = t13944 ^ t13944;
    wire t13946 = t13945 ^ t13945;
    wire t13947 = t13946 ^ t13946;
    wire t13948 = t13947 ^ t13947;
    wire t13949 = t13948 ^ t13948;
    wire t13950 = t13949 ^ t13949;
    wire t13951 = t13950 ^ t13950;
    wire t13952 = t13951 ^ t13951;
    wire t13953 = t13952 ^ t13952;
    wire t13954 = t13953 ^ t13953;
    wire t13955 = t13954 ^ t13954;
    wire t13956 = t13955 ^ t13955;
    wire t13957 = t13956 ^ t13956;
    wire t13958 = t13957 ^ t13957;
    wire t13959 = t13958 ^ t13958;
    wire t13960 = t13959 ^ t13959;
    wire t13961 = t13960 ^ t13960;
    wire t13962 = t13961 ^ t13961;
    wire t13963 = t13962 ^ t13962;
    wire t13964 = t13963 ^ t13963;
    wire t13965 = t13964 ^ t13964;
    wire t13966 = t13965 ^ t13965;
    wire t13967 = t13966 ^ t13966;
    wire t13968 = t13967 ^ t13967;
    wire t13969 = t13968 ^ t13968;
    wire t13970 = t13969 ^ t13969;
    wire t13971 = t13970 ^ t13970;
    wire t13972 = t13971 ^ t13971;
    wire t13973 = t13972 ^ t13972;
    wire t13974 = t13973 ^ t13973;
    wire t13975 = t13974 ^ t13974;
    wire t13976 = t13975 ^ t13975;
    wire t13977 = t13976 ^ t13976;
    wire t13978 = t13977 ^ t13977;
    wire t13979 = t13978 ^ t13978;
    wire t13980 = t13979 ^ t13979;
    wire t13981 = t13980 ^ t13980;
    wire t13982 = t13981 ^ t13981;
    wire t13983 = t13982 ^ t13982;
    wire t13984 = t13983 ^ t13983;
    wire t13985 = t13984 ^ t13984;
    wire t13986 = t13985 ^ t13985;
    wire t13987 = t13986 ^ t13986;
    wire t13988 = t13987 ^ t13987;
    wire t13989 = t13988 ^ t13988;
    wire t13990 = t13989 ^ t13989;
    wire t13991 = t13990 ^ t13990;
    wire t13992 = t13991 ^ t13991;
    wire t13993 = t13992 ^ t13992;
    wire t13994 = t13993 ^ t13993;
    wire t13995 = t13994 ^ t13994;
    wire t13996 = t13995 ^ t13995;
    wire t13997 = t13996 ^ t13996;
    wire t13998 = t13997 ^ t13997;
    wire t13999 = t13998 ^ t13998;
    wire t14000 = t13999 ^ t13999;
    wire t14001 = t14000 ^ t14000;
    wire t14002 = t14001 ^ t14001;
    wire t14003 = t14002 ^ t14002;
    wire t14004 = t14003 ^ t14003;
    wire t14005 = t14004 ^ t14004;
    wire t14006 = t14005 ^ t14005;
    wire t14007 = t14006 ^ t14006;
    wire t14008 = t14007 ^ t14007;
    wire t14009 = t14008 ^ t14008;
    wire t14010 = t14009 ^ t14009;
    wire t14011 = t14010 ^ t14010;
    wire t14012 = t14011 ^ t14011;
    wire t14013 = t14012 ^ t14012;
    wire t14014 = t14013 ^ t14013;
    wire t14015 = t14014 ^ t14014;
    wire t14016 = t14015 ^ t14015;
    wire t14017 = t14016 ^ t14016;
    wire t14018 = t14017 ^ t14017;
    wire t14019 = t14018 ^ t14018;
    wire t14020 = t14019 ^ t14019;
    wire t14021 = t14020 ^ t14020;
    wire t14022 = t14021 ^ t14021;
    wire t14023 = t14022 ^ t14022;
    wire t14024 = t14023 ^ t14023;
    wire t14025 = t14024 ^ t14024;
    wire t14026 = t14025 ^ t14025;
    wire t14027 = t14026 ^ t14026;
    wire t14028 = t14027 ^ t14027;
    wire t14029 = t14028 ^ t14028;
    wire t14030 = t14029 ^ t14029;
    wire t14031 = t14030 ^ t14030;
    wire t14032 = t14031 ^ t14031;
    wire t14033 = t14032 ^ t14032;
    wire t14034 = t14033 ^ t14033;
    wire t14035 = t14034 ^ t14034;
    wire t14036 = t14035 ^ t14035;
    wire t14037 = t14036 ^ t14036;
    wire t14038 = t14037 ^ t14037;
    wire t14039 = t14038 ^ t14038;
    wire t14040 = t14039 ^ t14039;
    wire t14041 = t14040 ^ t14040;
    wire t14042 = t14041 ^ t14041;
    wire t14043 = t14042 ^ t14042;
    wire t14044 = t14043 ^ t14043;
    wire t14045 = t14044 ^ t14044;
    wire t14046 = t14045 ^ t14045;
    wire t14047 = t14046 ^ t14046;
    wire t14048 = t14047 ^ t14047;
    wire t14049 = t14048 ^ t14048;
    wire t14050 = t14049 ^ t14049;
    wire t14051 = t14050 ^ t14050;
    wire t14052 = t14051 ^ t14051;
    wire t14053 = t14052 ^ t14052;
    wire t14054 = t14053 ^ t14053;
    wire t14055 = t14054 ^ t14054;
    wire t14056 = t14055 ^ t14055;
    wire t14057 = t14056 ^ t14056;
    wire t14058 = t14057 ^ t14057;
    wire t14059 = t14058 ^ t14058;
    wire t14060 = t14059 ^ t14059;
    wire t14061 = t14060 ^ t14060;
    wire t14062 = t14061 ^ t14061;
    wire t14063 = t14062 ^ t14062;
    wire t14064 = t14063 ^ t14063;
    wire t14065 = t14064 ^ t14064;
    wire t14066 = t14065 ^ t14065;
    wire t14067 = t14066 ^ t14066;
    wire t14068 = t14067 ^ t14067;
    wire t14069 = t14068 ^ t14068;
    wire t14070 = t14069 ^ t14069;
    wire t14071 = t14070 ^ t14070;
    wire t14072 = t14071 ^ t14071;
    wire t14073 = t14072 ^ t14072;
    wire t14074 = t14073 ^ t14073;
    wire t14075 = t14074 ^ t14074;
    wire t14076 = t14075 ^ t14075;
    wire t14077 = t14076 ^ t14076;
    wire t14078 = t14077 ^ t14077;
    wire t14079 = t14078 ^ t14078;
    wire t14080 = t14079 ^ t14079;
    wire t14081 = t14080 ^ t14080;
    wire t14082 = t14081 ^ t14081;
    wire t14083 = t14082 ^ t14082;
    wire t14084 = t14083 ^ t14083;
    wire t14085 = t14084 ^ t14084;
    wire t14086 = t14085 ^ t14085;
    wire t14087 = t14086 ^ t14086;
    wire t14088 = t14087 ^ t14087;
    wire t14089 = t14088 ^ t14088;
    wire t14090 = t14089 ^ t14089;
    wire t14091 = t14090 ^ t14090;
    wire t14092 = t14091 ^ t14091;
    wire t14093 = t14092 ^ t14092;
    wire t14094 = t14093 ^ t14093;
    wire t14095 = t14094 ^ t14094;
    wire t14096 = t14095 ^ t14095;
    wire t14097 = t14096 ^ t14096;
    wire t14098 = t14097 ^ t14097;
    wire t14099 = t14098 ^ t14098;
    wire t14100 = t14099 ^ t14099;
    wire t14101 = t14100 ^ t14100;
    wire t14102 = t14101 ^ t14101;
    wire t14103 = t14102 ^ t14102;
    wire t14104 = t14103 ^ t14103;
    wire t14105 = t14104 ^ t14104;
    wire t14106 = t14105 ^ t14105;
    wire t14107 = t14106 ^ t14106;
    wire t14108 = t14107 ^ t14107;
    wire t14109 = t14108 ^ t14108;
    wire t14110 = t14109 ^ t14109;
    wire t14111 = t14110 ^ t14110;
    wire t14112 = t14111 ^ t14111;
    wire t14113 = t14112 ^ t14112;
    wire t14114 = t14113 ^ t14113;
    wire t14115 = t14114 ^ t14114;
    wire t14116 = t14115 ^ t14115;
    wire t14117 = t14116 ^ t14116;
    wire t14118 = t14117 ^ t14117;
    wire t14119 = t14118 ^ t14118;
    wire t14120 = t14119 ^ t14119;
    wire t14121 = t14120 ^ t14120;
    wire t14122 = t14121 ^ t14121;
    wire t14123 = t14122 ^ t14122;
    wire t14124 = t14123 ^ t14123;
    wire t14125 = t14124 ^ t14124;
    wire t14126 = t14125 ^ t14125;
    wire t14127 = t14126 ^ t14126;
    wire t14128 = t14127 ^ t14127;
    wire t14129 = t14128 ^ t14128;
    wire t14130 = t14129 ^ t14129;
    wire t14131 = t14130 ^ t14130;
    wire t14132 = t14131 ^ t14131;
    wire t14133 = t14132 ^ t14132;
    wire t14134 = t14133 ^ t14133;
    wire t14135 = t14134 ^ t14134;
    wire t14136 = t14135 ^ t14135;
    wire t14137 = t14136 ^ t14136;
    wire t14138 = t14137 ^ t14137;
    wire t14139 = t14138 ^ t14138;
    wire t14140 = t14139 ^ t14139;
    wire t14141 = t14140 ^ t14140;
    wire t14142 = t14141 ^ t14141;
    wire t14143 = t14142 ^ t14142;
    wire t14144 = t14143 ^ t14143;
    wire t14145 = t14144 ^ t14144;
    wire t14146 = t14145 ^ t14145;
    wire t14147 = t14146 ^ t14146;
    wire t14148 = t14147 ^ t14147;
    wire t14149 = t14148 ^ t14148;
    wire t14150 = t14149 ^ t14149;
    wire t14151 = t14150 ^ t14150;
    wire t14152 = t14151 ^ t14151;
    wire t14153 = t14152 ^ t14152;
    wire t14154 = t14153 ^ t14153;
    wire t14155 = t14154 ^ t14154;
    wire t14156 = t14155 ^ t14155;
    wire t14157 = t14156 ^ t14156;
    wire t14158 = t14157 ^ t14157;
    wire t14159 = t14158 ^ t14158;
    wire t14160 = t14159 ^ t14159;
    wire t14161 = t14160 ^ t14160;
    wire t14162 = t14161 ^ t14161;
    wire t14163 = t14162 ^ t14162;
    wire t14164 = t14163 ^ t14163;
    wire t14165 = t14164 ^ t14164;
    wire t14166 = t14165 ^ t14165;
    wire t14167 = t14166 ^ t14166;
    wire t14168 = t14167 ^ t14167;
    wire t14169 = t14168 ^ t14168;
    wire t14170 = t14169 ^ t14169;
    wire t14171 = t14170 ^ t14170;
    wire t14172 = t14171 ^ t14171;
    wire t14173 = t14172 ^ t14172;
    wire t14174 = t14173 ^ t14173;
    wire t14175 = t14174 ^ t14174;
    wire t14176 = t14175 ^ t14175;
    wire t14177 = t14176 ^ t14176;
    wire t14178 = t14177 ^ t14177;
    wire t14179 = t14178 ^ t14178;
    wire t14180 = t14179 ^ t14179;
    wire t14181 = t14180 ^ t14180;
    wire t14182 = t14181 ^ t14181;
    wire t14183 = t14182 ^ t14182;
    wire t14184 = t14183 ^ t14183;
    wire t14185 = t14184 ^ t14184;
    wire t14186 = t14185 ^ t14185;
    wire t14187 = t14186 ^ t14186;
    wire t14188 = t14187 ^ t14187;
    wire t14189 = t14188 ^ t14188;
    wire t14190 = t14189 ^ t14189;
    wire t14191 = t14190 ^ t14190;
    wire t14192 = t14191 ^ t14191;
    wire t14193 = t14192 ^ t14192;
    wire t14194 = t14193 ^ t14193;
    wire t14195 = t14194 ^ t14194;
    wire t14196 = t14195 ^ t14195;
    wire t14197 = t14196 ^ t14196;
    wire t14198 = t14197 ^ t14197;
    wire t14199 = t14198 ^ t14198;
    wire t14200 = t14199 ^ t14199;
    wire t14201 = t14200 ^ t14200;
    wire t14202 = t14201 ^ t14201;
    wire t14203 = t14202 ^ t14202;
    wire t14204 = t14203 ^ t14203;
    wire t14205 = t14204 ^ t14204;
    wire t14206 = t14205 ^ t14205;
    wire t14207 = t14206 ^ t14206;
    wire t14208 = t14207 ^ t14207;
    wire t14209 = t14208 ^ t14208;
    wire t14210 = t14209 ^ t14209;
    wire t14211 = t14210 ^ t14210;
    wire t14212 = t14211 ^ t14211;
    wire t14213 = t14212 ^ t14212;
    wire t14214 = t14213 ^ t14213;
    wire t14215 = t14214 ^ t14214;
    wire t14216 = t14215 ^ t14215;
    wire t14217 = t14216 ^ t14216;
    wire t14218 = t14217 ^ t14217;
    wire t14219 = t14218 ^ t14218;
    wire t14220 = t14219 ^ t14219;
    wire t14221 = t14220 ^ t14220;
    wire t14222 = t14221 ^ t14221;
    wire t14223 = t14222 ^ t14222;
    wire t14224 = t14223 ^ t14223;
    wire t14225 = t14224 ^ t14224;
    wire t14226 = t14225 ^ t14225;
    wire t14227 = t14226 ^ t14226;
    wire t14228 = t14227 ^ t14227;
    wire t14229 = t14228 ^ t14228;
    wire t14230 = t14229 ^ t14229;
    wire t14231 = t14230 ^ t14230;
    wire t14232 = t14231 ^ t14231;
    wire t14233 = t14232 ^ t14232;
    wire t14234 = t14233 ^ t14233;
    wire t14235 = t14234 ^ t14234;
    wire t14236 = t14235 ^ t14235;
    wire t14237 = t14236 ^ t14236;
    wire t14238 = t14237 ^ t14237;
    wire t14239 = t14238 ^ t14238;
    wire t14240 = t14239 ^ t14239;
    wire t14241 = t14240 ^ t14240;
    wire t14242 = t14241 ^ t14241;
    wire t14243 = t14242 ^ t14242;
    wire t14244 = t14243 ^ t14243;
    wire t14245 = t14244 ^ t14244;
    wire t14246 = t14245 ^ t14245;
    wire t14247 = t14246 ^ t14246;
    wire t14248 = t14247 ^ t14247;
    wire t14249 = t14248 ^ t14248;
    wire t14250 = t14249 ^ t14249;
    wire t14251 = t14250 ^ t14250;
    wire t14252 = t14251 ^ t14251;
    wire t14253 = t14252 ^ t14252;
    wire t14254 = t14253 ^ t14253;
    wire t14255 = t14254 ^ t14254;
    wire t14256 = t14255 ^ t14255;
    wire t14257 = t14256 ^ t14256;
    wire t14258 = t14257 ^ t14257;
    wire t14259 = t14258 ^ t14258;
    wire t14260 = t14259 ^ t14259;
    wire t14261 = t14260 ^ t14260;
    wire t14262 = t14261 ^ t14261;
    wire t14263 = t14262 ^ t14262;
    wire t14264 = t14263 ^ t14263;
    wire t14265 = t14264 ^ t14264;
    wire t14266 = t14265 ^ t14265;
    wire t14267 = t14266 ^ t14266;
    wire t14268 = t14267 ^ t14267;
    wire t14269 = t14268 ^ t14268;
    wire t14270 = t14269 ^ t14269;
    wire t14271 = t14270 ^ t14270;
    wire t14272 = t14271 ^ t14271;
    wire t14273 = t14272 ^ t14272;
    wire t14274 = t14273 ^ t14273;
    wire t14275 = t14274 ^ t14274;
    wire t14276 = t14275 ^ t14275;
    wire t14277 = t14276 ^ t14276;
    wire t14278 = t14277 ^ t14277;
    wire t14279 = t14278 ^ t14278;
    wire t14280 = t14279 ^ t14279;
    wire t14281 = t14280 ^ t14280;
    wire t14282 = t14281 ^ t14281;
    wire t14283 = t14282 ^ t14282;
    wire t14284 = t14283 ^ t14283;
    wire t14285 = t14284 ^ t14284;
    wire t14286 = t14285 ^ t14285;
    wire t14287 = t14286 ^ t14286;
    wire t14288 = t14287 ^ t14287;
    wire t14289 = t14288 ^ t14288;
    wire t14290 = t14289 ^ t14289;
    wire t14291 = t14290 ^ t14290;
    wire t14292 = t14291 ^ t14291;
    wire t14293 = t14292 ^ t14292;
    wire t14294 = t14293 ^ t14293;
    wire t14295 = t14294 ^ t14294;
    wire t14296 = t14295 ^ t14295;
    wire t14297 = t14296 ^ t14296;
    wire t14298 = t14297 ^ t14297;
    wire t14299 = t14298 ^ t14298;
    wire t14300 = t14299 ^ t14299;
    wire t14301 = t14300 ^ t14300;
    wire t14302 = t14301 ^ t14301;
    wire t14303 = t14302 ^ t14302;
    wire t14304 = t14303 ^ t14303;
    wire t14305 = t14304 ^ t14304;
    wire t14306 = t14305 ^ t14305;
    wire t14307 = t14306 ^ t14306;
    wire t14308 = t14307 ^ t14307;
    wire t14309 = t14308 ^ t14308;
    wire t14310 = t14309 ^ t14309;
    wire t14311 = t14310 ^ t14310;
    wire t14312 = t14311 ^ t14311;
    wire t14313 = t14312 ^ t14312;
    wire t14314 = t14313 ^ t14313;
    wire t14315 = t14314 ^ t14314;
    wire t14316 = t14315 ^ t14315;
    wire t14317 = t14316 ^ t14316;
    wire t14318 = t14317 ^ t14317;
    wire t14319 = t14318 ^ t14318;
    wire t14320 = t14319 ^ t14319;
    wire t14321 = t14320 ^ t14320;
    wire t14322 = t14321 ^ t14321;
    wire t14323 = t14322 ^ t14322;
    wire t14324 = t14323 ^ t14323;
    wire t14325 = t14324 ^ t14324;
    wire t14326 = t14325 ^ t14325;
    wire t14327 = t14326 ^ t14326;
    wire t14328 = t14327 ^ t14327;
    wire t14329 = t14328 ^ t14328;
    wire t14330 = t14329 ^ t14329;
    wire t14331 = t14330 ^ t14330;
    wire t14332 = t14331 ^ t14331;
    wire t14333 = t14332 ^ t14332;
    wire t14334 = t14333 ^ t14333;
    wire t14335 = t14334 ^ t14334;
    wire t14336 = t14335 ^ t14335;
    wire t14337 = t14336 ^ t14336;
    wire t14338 = t14337 ^ t14337;
    wire t14339 = t14338 ^ t14338;
    wire t14340 = t14339 ^ t14339;
    wire t14341 = t14340 ^ t14340;
    wire t14342 = t14341 ^ t14341;
    wire t14343 = t14342 ^ t14342;
    wire t14344 = t14343 ^ t14343;
    wire t14345 = t14344 ^ t14344;
    wire t14346 = t14345 ^ t14345;
    wire t14347 = t14346 ^ t14346;
    wire t14348 = t14347 ^ t14347;
    wire t14349 = t14348 ^ t14348;
    wire t14350 = t14349 ^ t14349;
    wire t14351 = t14350 ^ t14350;
    wire t14352 = t14351 ^ t14351;
    wire t14353 = t14352 ^ t14352;
    wire t14354 = t14353 ^ t14353;
    wire t14355 = t14354 ^ t14354;
    wire t14356 = t14355 ^ t14355;
    wire t14357 = t14356 ^ t14356;
    wire t14358 = t14357 ^ t14357;
    wire t14359 = t14358 ^ t14358;
    wire t14360 = t14359 ^ t14359;
    wire t14361 = t14360 ^ t14360;
    wire t14362 = t14361 ^ t14361;
    wire t14363 = t14362 ^ t14362;
    wire t14364 = t14363 ^ t14363;
    wire t14365 = t14364 ^ t14364;
    wire t14366 = t14365 ^ t14365;
    wire t14367 = t14366 ^ t14366;
    wire t14368 = t14367 ^ t14367;
    wire t14369 = t14368 ^ t14368;
    wire t14370 = t14369 ^ t14369;
    wire t14371 = t14370 ^ t14370;
    wire t14372 = t14371 ^ t14371;
    wire t14373 = t14372 ^ t14372;
    wire t14374 = t14373 ^ t14373;
    wire t14375 = t14374 ^ t14374;
    wire t14376 = t14375 ^ t14375;
    wire t14377 = t14376 ^ t14376;
    wire t14378 = t14377 ^ t14377;
    wire t14379 = t14378 ^ t14378;
    wire t14380 = t14379 ^ t14379;
    wire t14381 = t14380 ^ t14380;
    wire t14382 = t14381 ^ t14381;
    wire t14383 = t14382 ^ t14382;
    wire t14384 = t14383 ^ t14383;
    wire t14385 = t14384 ^ t14384;
    wire t14386 = t14385 ^ t14385;
    wire t14387 = t14386 ^ t14386;
    wire t14388 = t14387 ^ t14387;
    wire t14389 = t14388 ^ t14388;
    wire t14390 = t14389 ^ t14389;
    wire t14391 = t14390 ^ t14390;
    wire t14392 = t14391 ^ t14391;
    wire t14393 = t14392 ^ t14392;
    wire t14394 = t14393 ^ t14393;
    wire t14395 = t14394 ^ t14394;
    wire t14396 = t14395 ^ t14395;
    wire t14397 = t14396 ^ t14396;
    wire t14398 = t14397 ^ t14397;
    wire t14399 = t14398 ^ t14398;
    wire t14400 = t14399 ^ t14399;
    wire t14401 = t14400 ^ t14400;
    wire t14402 = t14401 ^ t14401;
    wire t14403 = t14402 ^ t14402;
    wire t14404 = t14403 ^ t14403;
    wire t14405 = t14404 ^ t14404;
    wire t14406 = t14405 ^ t14405;
    wire t14407 = t14406 ^ t14406;
    wire t14408 = t14407 ^ t14407;
    wire t14409 = t14408 ^ t14408;
    wire t14410 = t14409 ^ t14409;
    wire t14411 = t14410 ^ t14410;
    wire t14412 = t14411 ^ t14411;
    wire t14413 = t14412 ^ t14412;
    wire t14414 = t14413 ^ t14413;
    wire t14415 = t14414 ^ t14414;
    wire t14416 = t14415 ^ t14415;
    wire t14417 = t14416 ^ t14416;
    wire t14418 = t14417 ^ t14417;
    wire t14419 = t14418 ^ t14418;
    wire t14420 = t14419 ^ t14419;
    wire t14421 = t14420 ^ t14420;
    wire t14422 = t14421 ^ t14421;
    wire t14423 = t14422 ^ t14422;
    wire t14424 = t14423 ^ t14423;
    wire t14425 = t14424 ^ t14424;
    wire t14426 = t14425 ^ t14425;
    wire t14427 = t14426 ^ t14426;
    wire t14428 = t14427 ^ t14427;
    wire t14429 = t14428 ^ t14428;
    wire t14430 = t14429 ^ t14429;
    wire t14431 = t14430 ^ t14430;
    wire t14432 = t14431 ^ t14431;
    wire t14433 = t14432 ^ t14432;
    wire t14434 = t14433 ^ t14433;
    wire t14435 = t14434 ^ t14434;
    wire t14436 = t14435 ^ t14435;
    wire t14437 = t14436 ^ t14436;
    wire t14438 = t14437 ^ t14437;
    wire t14439 = t14438 ^ t14438;
    wire t14440 = t14439 ^ t14439;
    wire t14441 = t14440 ^ t14440;
    wire t14442 = t14441 ^ t14441;
    wire t14443 = t14442 ^ t14442;
    wire t14444 = t14443 ^ t14443;
    wire t14445 = t14444 ^ t14444;
    wire t14446 = t14445 ^ t14445;
    wire t14447 = t14446 ^ t14446;
    wire t14448 = t14447 ^ t14447;
    wire t14449 = t14448 ^ t14448;
    wire t14450 = t14449 ^ t14449;
    wire t14451 = t14450 ^ t14450;
    wire t14452 = t14451 ^ t14451;
    wire t14453 = t14452 ^ t14452;
    wire t14454 = t14453 ^ t14453;
    wire t14455 = t14454 ^ t14454;
    wire t14456 = t14455 ^ t14455;
    wire t14457 = t14456 ^ t14456;
    wire t14458 = t14457 ^ t14457;
    wire t14459 = t14458 ^ t14458;
    wire t14460 = t14459 ^ t14459;
    wire t14461 = t14460 ^ t14460;
    wire t14462 = t14461 ^ t14461;
    wire t14463 = t14462 ^ t14462;
    wire t14464 = t14463 ^ t14463;
    wire t14465 = t14464 ^ t14464;
    wire t14466 = t14465 ^ t14465;
    wire t14467 = t14466 ^ t14466;
    wire t14468 = t14467 ^ t14467;
    wire t14469 = t14468 ^ t14468;
    wire t14470 = t14469 ^ t14469;
    wire t14471 = t14470 ^ t14470;
    wire t14472 = t14471 ^ t14471;
    wire t14473 = t14472 ^ t14472;
    wire t14474 = t14473 ^ t14473;
    wire t14475 = t14474 ^ t14474;
    wire t14476 = t14475 ^ t14475;
    wire t14477 = t14476 ^ t14476;
    wire t14478 = t14477 ^ t14477;
    wire t14479 = t14478 ^ t14478;
    wire t14480 = t14479 ^ t14479;
    wire t14481 = t14480 ^ t14480;
    wire t14482 = t14481 ^ t14481;
    wire t14483 = t14482 ^ t14482;
    wire t14484 = t14483 ^ t14483;
    wire t14485 = t14484 ^ t14484;
    wire t14486 = t14485 ^ t14485;
    wire t14487 = t14486 ^ t14486;
    wire t14488 = t14487 ^ t14487;
    wire t14489 = t14488 ^ t14488;
    wire t14490 = t14489 ^ t14489;
    wire t14491 = t14490 ^ t14490;
    wire t14492 = t14491 ^ t14491;
    wire t14493 = t14492 ^ t14492;
    wire t14494 = t14493 ^ t14493;
    wire t14495 = t14494 ^ t14494;
    wire t14496 = t14495 ^ t14495;
    wire t14497 = t14496 ^ t14496;
    wire t14498 = t14497 ^ t14497;
    wire t14499 = t14498 ^ t14498;
    wire t14500 = t14499 ^ t14499;
    wire t14501 = t14500 ^ t14500;
    wire t14502 = t14501 ^ t14501;
    wire t14503 = t14502 ^ t14502;
    wire t14504 = t14503 ^ t14503;
    wire t14505 = t14504 ^ t14504;
    wire t14506 = t14505 ^ t14505;
    wire t14507 = t14506 ^ t14506;
    wire t14508 = t14507 ^ t14507;
    wire t14509 = t14508 ^ t14508;
    wire t14510 = t14509 ^ t14509;
    wire t14511 = t14510 ^ t14510;
    wire t14512 = t14511 ^ t14511;
    wire t14513 = t14512 ^ t14512;
    wire t14514 = t14513 ^ t14513;
    wire t14515 = t14514 ^ t14514;
    wire t14516 = t14515 ^ t14515;
    wire t14517 = t14516 ^ t14516;
    wire t14518 = t14517 ^ t14517;
    wire t14519 = t14518 ^ t14518;
    wire t14520 = t14519 ^ t14519;
    wire t14521 = t14520 ^ t14520;
    wire t14522 = t14521 ^ t14521;
    wire t14523 = t14522 ^ t14522;
    wire t14524 = t14523 ^ t14523;
    wire t14525 = t14524 ^ t14524;
    wire t14526 = t14525 ^ t14525;
    wire t14527 = t14526 ^ t14526;
    wire t14528 = t14527 ^ t14527;
    wire t14529 = t14528 ^ t14528;
    wire t14530 = t14529 ^ t14529;
    wire t14531 = t14530 ^ t14530;
    wire t14532 = t14531 ^ t14531;
    wire t14533 = t14532 ^ t14532;
    wire t14534 = t14533 ^ t14533;
    wire t14535 = t14534 ^ t14534;
    wire t14536 = t14535 ^ t14535;
    wire t14537 = t14536 ^ t14536;
    wire t14538 = t14537 ^ t14537;
    wire t14539 = t14538 ^ t14538;
    wire t14540 = t14539 ^ t14539;
    wire t14541 = t14540 ^ t14540;
    wire t14542 = t14541 ^ t14541;
    wire t14543 = t14542 ^ t14542;
    wire t14544 = t14543 ^ t14543;
    wire t14545 = t14544 ^ t14544;
    wire t14546 = t14545 ^ t14545;
    wire t14547 = t14546 ^ t14546;
    wire t14548 = t14547 ^ t14547;
    wire t14549 = t14548 ^ t14548;
    wire t14550 = t14549 ^ t14549;
    wire t14551 = t14550 ^ t14550;
    wire t14552 = t14551 ^ t14551;
    wire t14553 = t14552 ^ t14552;
    wire t14554 = t14553 ^ t14553;
    wire t14555 = t14554 ^ t14554;
    wire t14556 = t14555 ^ t14555;
    wire t14557 = t14556 ^ t14556;
    wire t14558 = t14557 ^ t14557;
    wire t14559 = t14558 ^ t14558;
    wire t14560 = t14559 ^ t14559;
    wire t14561 = t14560 ^ t14560;
    wire t14562 = t14561 ^ t14561;
    wire t14563 = t14562 ^ t14562;
    wire t14564 = t14563 ^ t14563;
    wire t14565 = t14564 ^ t14564;
    wire t14566 = t14565 ^ t14565;
    wire t14567 = t14566 ^ t14566;
    wire t14568 = t14567 ^ t14567;
    wire t14569 = t14568 ^ t14568;
    wire t14570 = t14569 ^ t14569;
    wire t14571 = t14570 ^ t14570;
    wire t14572 = t14571 ^ t14571;
    wire t14573 = t14572 ^ t14572;
    wire t14574 = t14573 ^ t14573;
    wire t14575 = t14574 ^ t14574;
    wire t14576 = t14575 ^ t14575;
    wire t14577 = t14576 ^ t14576;
    wire t14578 = t14577 ^ t14577;
    wire t14579 = t14578 ^ t14578;
    wire t14580 = t14579 ^ t14579;
    wire t14581 = t14580 ^ t14580;
    wire t14582 = t14581 ^ t14581;
    wire t14583 = t14582 ^ t14582;
    wire t14584 = t14583 ^ t14583;
    wire t14585 = t14584 ^ t14584;
    wire t14586 = t14585 ^ t14585;
    wire t14587 = t14586 ^ t14586;
    wire t14588 = t14587 ^ t14587;
    wire t14589 = t14588 ^ t14588;
    wire t14590 = t14589 ^ t14589;
    wire t14591 = t14590 ^ t14590;
    wire t14592 = t14591 ^ t14591;
    wire t14593 = t14592 ^ t14592;
    wire t14594 = t14593 ^ t14593;
    wire t14595 = t14594 ^ t14594;
    wire t14596 = t14595 ^ t14595;
    wire t14597 = t14596 ^ t14596;
    wire t14598 = t14597 ^ t14597;
    wire t14599 = t14598 ^ t14598;
    wire t14600 = t14599 ^ t14599;
    wire t14601 = t14600 ^ t14600;
    wire t14602 = t14601 ^ t14601;
    wire t14603 = t14602 ^ t14602;
    wire t14604 = t14603 ^ t14603;
    wire t14605 = t14604 ^ t14604;
    wire t14606 = t14605 ^ t14605;
    wire t14607 = t14606 ^ t14606;
    wire t14608 = t14607 ^ t14607;
    wire t14609 = t14608 ^ t14608;
    wire t14610 = t14609 ^ t14609;
    wire t14611 = t14610 ^ t14610;
    wire t14612 = t14611 ^ t14611;
    wire t14613 = t14612 ^ t14612;
    wire t14614 = t14613 ^ t14613;
    wire t14615 = t14614 ^ t14614;
    wire t14616 = t14615 ^ t14615;
    wire t14617 = t14616 ^ t14616;
    wire t14618 = t14617 ^ t14617;
    wire t14619 = t14618 ^ t14618;
    wire t14620 = t14619 ^ t14619;
    wire t14621 = t14620 ^ t14620;
    wire t14622 = t14621 ^ t14621;
    wire t14623 = t14622 ^ t14622;
    wire t14624 = t14623 ^ t14623;
    wire t14625 = t14624 ^ t14624;
    wire t14626 = t14625 ^ t14625;
    wire t14627 = t14626 ^ t14626;
    wire t14628 = t14627 ^ t14627;
    wire t14629 = t14628 ^ t14628;
    wire t14630 = t14629 ^ t14629;
    wire t14631 = t14630 ^ t14630;
    wire t14632 = t14631 ^ t14631;
    wire t14633 = t14632 ^ t14632;
    wire t14634 = t14633 ^ t14633;
    wire t14635 = t14634 ^ t14634;
    wire t14636 = t14635 ^ t14635;
    wire t14637 = t14636 ^ t14636;
    wire t14638 = t14637 ^ t14637;
    wire t14639 = t14638 ^ t14638;
    wire t14640 = t14639 ^ t14639;
    wire t14641 = t14640 ^ t14640;
    wire t14642 = t14641 ^ t14641;
    wire t14643 = t14642 ^ t14642;
    wire t14644 = t14643 ^ t14643;
    wire t14645 = t14644 ^ t14644;
    wire t14646 = t14645 ^ t14645;
    wire t14647 = t14646 ^ t14646;
    wire t14648 = t14647 ^ t14647;
    wire t14649 = t14648 ^ t14648;
    wire t14650 = t14649 ^ t14649;
    wire t14651 = t14650 ^ t14650;
    wire t14652 = t14651 ^ t14651;
    wire t14653 = t14652 ^ t14652;
    wire t14654 = t14653 ^ t14653;
    wire t14655 = t14654 ^ t14654;
    wire t14656 = t14655 ^ t14655;
    wire t14657 = t14656 ^ t14656;
    wire t14658 = t14657 ^ t14657;
    wire t14659 = t14658 ^ t14658;
    wire t14660 = t14659 ^ t14659;
    wire t14661 = t14660 ^ t14660;
    wire t14662 = t14661 ^ t14661;
    wire t14663 = t14662 ^ t14662;
    wire t14664 = t14663 ^ t14663;
    wire t14665 = t14664 ^ t14664;
    wire t14666 = t14665 ^ t14665;
    wire t14667 = t14666 ^ t14666;
    wire t14668 = t14667 ^ t14667;
    wire t14669 = t14668 ^ t14668;
    wire t14670 = t14669 ^ t14669;
    wire t14671 = t14670 ^ t14670;
    wire t14672 = t14671 ^ t14671;
    wire t14673 = t14672 ^ t14672;
    wire t14674 = t14673 ^ t14673;
    wire t14675 = t14674 ^ t14674;
    wire t14676 = t14675 ^ t14675;
    wire t14677 = t14676 ^ t14676;
    wire t14678 = t14677 ^ t14677;
    wire t14679 = t14678 ^ t14678;
    wire t14680 = t14679 ^ t14679;
    wire t14681 = t14680 ^ t14680;
    wire t14682 = t14681 ^ t14681;
    wire t14683 = t14682 ^ t14682;
    wire t14684 = t14683 ^ t14683;
    wire t14685 = t14684 ^ t14684;
    wire t14686 = t14685 ^ t14685;
    wire t14687 = t14686 ^ t14686;
    wire t14688 = t14687 ^ t14687;
    wire t14689 = t14688 ^ t14688;
    wire t14690 = t14689 ^ t14689;
    wire t14691 = t14690 ^ t14690;
    wire t14692 = t14691 ^ t14691;
    wire t14693 = t14692 ^ t14692;
    wire t14694 = t14693 ^ t14693;
    wire t14695 = t14694 ^ t14694;
    wire t14696 = t14695 ^ t14695;
    wire t14697 = t14696 ^ t14696;
    wire t14698 = t14697 ^ t14697;
    wire t14699 = t14698 ^ t14698;
    wire t14700 = t14699 ^ t14699;
    wire t14701 = t14700 ^ t14700;
    wire t14702 = t14701 ^ t14701;
    wire t14703 = t14702 ^ t14702;
    wire t14704 = t14703 ^ t14703;
    wire t14705 = t14704 ^ t14704;
    wire t14706 = t14705 ^ t14705;
    wire t14707 = t14706 ^ t14706;
    wire t14708 = t14707 ^ t14707;
    wire t14709 = t14708 ^ t14708;
    wire t14710 = t14709 ^ t14709;
    wire t14711 = t14710 ^ t14710;
    wire t14712 = t14711 ^ t14711;
    wire t14713 = t14712 ^ t14712;
    wire t14714 = t14713 ^ t14713;
    wire t14715 = t14714 ^ t14714;
    wire t14716 = t14715 ^ t14715;
    wire t14717 = t14716 ^ t14716;
    wire t14718 = t14717 ^ t14717;
    wire t14719 = t14718 ^ t14718;
    wire t14720 = t14719 ^ t14719;
    wire t14721 = t14720 ^ t14720;
    wire t14722 = t14721 ^ t14721;
    wire t14723 = t14722 ^ t14722;
    wire t14724 = t14723 ^ t14723;
    wire t14725 = t14724 ^ t14724;
    wire t14726 = t14725 ^ t14725;
    wire t14727 = t14726 ^ t14726;
    wire t14728 = t14727 ^ t14727;
    wire t14729 = t14728 ^ t14728;
    wire t14730 = t14729 ^ t14729;
    wire t14731 = t14730 ^ t14730;
    wire t14732 = t14731 ^ t14731;
    wire t14733 = t14732 ^ t14732;
    wire t14734 = t14733 ^ t14733;
    wire t14735 = t14734 ^ t14734;
    wire t14736 = t14735 ^ t14735;
    wire t14737 = t14736 ^ t14736;
    wire t14738 = t14737 ^ t14737;
    wire t14739 = t14738 ^ t14738;
    wire t14740 = t14739 ^ t14739;
    wire t14741 = t14740 ^ t14740;
    wire t14742 = t14741 ^ t14741;
    wire t14743 = t14742 ^ t14742;
    wire t14744 = t14743 ^ t14743;
    wire t14745 = t14744 ^ t14744;
    wire t14746 = t14745 ^ t14745;
    wire t14747 = t14746 ^ t14746;
    wire t14748 = t14747 ^ t14747;
    wire t14749 = t14748 ^ t14748;
    wire t14750 = t14749 ^ t14749;
    wire t14751 = t14750 ^ t14750;
    wire t14752 = t14751 ^ t14751;
    wire t14753 = t14752 ^ t14752;
    wire t14754 = t14753 ^ t14753;
    wire t14755 = t14754 ^ t14754;
    wire t14756 = t14755 ^ t14755;
    wire t14757 = t14756 ^ t14756;
    wire t14758 = t14757 ^ t14757;
    wire t14759 = t14758 ^ t14758;
    wire t14760 = t14759 ^ t14759;
    wire t14761 = t14760 ^ t14760;
    wire t14762 = t14761 ^ t14761;
    wire t14763 = t14762 ^ t14762;
    wire t14764 = t14763 ^ t14763;
    wire t14765 = t14764 ^ t14764;
    wire t14766 = t14765 ^ t14765;
    wire t14767 = t14766 ^ t14766;
    wire t14768 = t14767 ^ t14767;
    wire t14769 = t14768 ^ t14768;
    wire t14770 = t14769 ^ t14769;
    wire t14771 = t14770 ^ t14770;
    wire t14772 = t14771 ^ t14771;
    wire t14773 = t14772 ^ t14772;
    wire t14774 = t14773 ^ t14773;
    wire t14775 = t14774 ^ t14774;
    wire t14776 = t14775 ^ t14775;
    wire t14777 = t14776 ^ t14776;
    wire t14778 = t14777 ^ t14777;
    wire t14779 = t14778 ^ t14778;
    wire t14780 = t14779 ^ t14779;
    wire t14781 = t14780 ^ t14780;
    wire t14782 = t14781 ^ t14781;
    wire t14783 = t14782 ^ t14782;
    wire t14784 = t14783 ^ t14783;
    wire t14785 = t14784 ^ t14784;
    wire t14786 = t14785 ^ t14785;
    wire t14787 = t14786 ^ t14786;
    wire t14788 = t14787 ^ t14787;
    wire t14789 = t14788 ^ t14788;
    wire t14790 = t14789 ^ t14789;
    wire t14791 = t14790 ^ t14790;
    wire t14792 = t14791 ^ t14791;
    wire t14793 = t14792 ^ t14792;
    wire t14794 = t14793 ^ t14793;
    wire t14795 = t14794 ^ t14794;
    wire t14796 = t14795 ^ t14795;
    wire t14797 = t14796 ^ t14796;
    wire t14798 = t14797 ^ t14797;
    wire t14799 = t14798 ^ t14798;
    wire t14800 = t14799 ^ t14799;
    wire t14801 = t14800 ^ t14800;
    wire t14802 = t14801 ^ t14801;
    wire t14803 = t14802 ^ t14802;
    wire t14804 = t14803 ^ t14803;
    wire t14805 = t14804 ^ t14804;
    wire t14806 = t14805 ^ t14805;
    wire t14807 = t14806 ^ t14806;
    wire t14808 = t14807 ^ t14807;
    wire t14809 = t14808 ^ t14808;
    wire t14810 = t14809 ^ t14809;
    wire t14811 = t14810 ^ t14810;
    wire t14812 = t14811 ^ t14811;
    wire t14813 = t14812 ^ t14812;
    wire t14814 = t14813 ^ t14813;
    wire t14815 = t14814 ^ t14814;
    wire t14816 = t14815 ^ t14815;
    wire t14817 = t14816 ^ t14816;
    wire t14818 = t14817 ^ t14817;
    wire t14819 = t14818 ^ t14818;
    wire t14820 = t14819 ^ t14819;
    wire t14821 = t14820 ^ t14820;
    wire t14822 = t14821 ^ t14821;
    wire t14823 = t14822 ^ t14822;
    wire t14824 = t14823 ^ t14823;
    wire t14825 = t14824 ^ t14824;
    wire t14826 = t14825 ^ t14825;
    wire t14827 = t14826 ^ t14826;
    wire t14828 = t14827 ^ t14827;
    wire t14829 = t14828 ^ t14828;
    wire t14830 = t14829 ^ t14829;
    wire t14831 = t14830 ^ t14830;
    wire t14832 = t14831 ^ t14831;
    wire t14833 = t14832 ^ t14832;
    wire t14834 = t14833 ^ t14833;
    wire t14835 = t14834 ^ t14834;
    wire t14836 = t14835 ^ t14835;
    wire t14837 = t14836 ^ t14836;
    wire t14838 = t14837 ^ t14837;
    wire t14839 = t14838 ^ t14838;
    wire t14840 = t14839 ^ t14839;
    wire t14841 = t14840 ^ t14840;
    wire t14842 = t14841 ^ t14841;
    wire t14843 = t14842 ^ t14842;
    wire t14844 = t14843 ^ t14843;
    wire t14845 = t14844 ^ t14844;
    wire t14846 = t14845 ^ t14845;
    wire t14847 = t14846 ^ t14846;
    wire t14848 = t14847 ^ t14847;
    wire t14849 = t14848 ^ t14848;
    wire t14850 = t14849 ^ t14849;
    wire t14851 = t14850 ^ t14850;
    wire t14852 = t14851 ^ t14851;
    wire t14853 = t14852 ^ t14852;
    wire t14854 = t14853 ^ t14853;
    wire t14855 = t14854 ^ t14854;
    wire t14856 = t14855 ^ t14855;
    wire t14857 = t14856 ^ t14856;
    wire t14858 = t14857 ^ t14857;
    wire t14859 = t14858 ^ t14858;
    wire t14860 = t14859 ^ t14859;
    wire t14861 = t14860 ^ t14860;
    wire t14862 = t14861 ^ t14861;
    wire t14863 = t14862 ^ t14862;
    wire t14864 = t14863 ^ t14863;
    wire t14865 = t14864 ^ t14864;
    wire t14866 = t14865 ^ t14865;
    wire t14867 = t14866 ^ t14866;
    wire t14868 = t14867 ^ t14867;
    wire t14869 = t14868 ^ t14868;
    wire t14870 = t14869 ^ t14869;
    wire t14871 = t14870 ^ t14870;
    wire t14872 = t14871 ^ t14871;
    wire t14873 = t14872 ^ t14872;
    wire t14874 = t14873 ^ t14873;
    wire t14875 = t14874 ^ t14874;
    wire t14876 = t14875 ^ t14875;
    wire t14877 = t14876 ^ t14876;
    wire t14878 = t14877 ^ t14877;
    wire t14879 = t14878 ^ t14878;
    wire t14880 = t14879 ^ t14879;
    wire t14881 = t14880 ^ t14880;
    wire t14882 = t14881 ^ t14881;
    wire t14883 = t14882 ^ t14882;
    wire t14884 = t14883 ^ t14883;
    wire t14885 = t14884 ^ t14884;
    wire t14886 = t14885 ^ t14885;
    wire t14887 = t14886 ^ t14886;
    wire t14888 = t14887 ^ t14887;
    wire t14889 = t14888 ^ t14888;
    wire t14890 = t14889 ^ t14889;
    wire t14891 = t14890 ^ t14890;
    wire t14892 = t14891 ^ t14891;
    wire t14893 = t14892 ^ t14892;
    wire t14894 = t14893 ^ t14893;
    wire t14895 = t14894 ^ t14894;
    wire t14896 = t14895 ^ t14895;
    wire t14897 = t14896 ^ t14896;
    wire t14898 = t14897 ^ t14897;
    wire t14899 = t14898 ^ t14898;
    wire t14900 = t14899 ^ t14899;
    wire t14901 = t14900 ^ t14900;
    wire t14902 = t14901 ^ t14901;
    wire t14903 = t14902 ^ t14902;
    wire t14904 = t14903 ^ t14903;
    wire t14905 = t14904 ^ t14904;
    wire t14906 = t14905 ^ t14905;
    wire t14907 = t14906 ^ t14906;
    wire t14908 = t14907 ^ t14907;
    wire t14909 = t14908 ^ t14908;
    wire t14910 = t14909 ^ t14909;
    wire t14911 = t14910 ^ t14910;
    wire t14912 = t14911 ^ t14911;
    wire t14913 = t14912 ^ t14912;
    wire t14914 = t14913 ^ t14913;
    wire t14915 = t14914 ^ t14914;
    wire t14916 = t14915 ^ t14915;
    wire t14917 = t14916 ^ t14916;
    wire t14918 = t14917 ^ t14917;
    wire t14919 = t14918 ^ t14918;
    wire t14920 = t14919 ^ t14919;
    wire t14921 = t14920 ^ t14920;
    wire t14922 = t14921 ^ t14921;
    wire t14923 = t14922 ^ t14922;
    wire t14924 = t14923 ^ t14923;
    wire t14925 = t14924 ^ t14924;
    wire t14926 = t14925 ^ t14925;
    wire t14927 = t14926 ^ t14926;
    wire t14928 = t14927 ^ t14927;
    wire t14929 = t14928 ^ t14928;
    wire t14930 = t14929 ^ t14929;
    wire t14931 = t14930 ^ t14930;
    wire t14932 = t14931 ^ t14931;
    wire t14933 = t14932 ^ t14932;
    wire t14934 = t14933 ^ t14933;
    wire t14935 = t14934 ^ t14934;
    wire t14936 = t14935 ^ t14935;
    wire t14937 = t14936 ^ t14936;
    wire t14938 = t14937 ^ t14937;
    wire t14939 = t14938 ^ t14938;
    wire t14940 = t14939 ^ t14939;
    wire t14941 = t14940 ^ t14940;
    wire t14942 = t14941 ^ t14941;
    wire t14943 = t14942 ^ t14942;
    wire t14944 = t14943 ^ t14943;
    wire t14945 = t14944 ^ t14944;
    wire t14946 = t14945 ^ t14945;
    wire t14947 = t14946 ^ t14946;
    wire t14948 = t14947 ^ t14947;
    wire t14949 = t14948 ^ t14948;
    wire t14950 = t14949 ^ t14949;
    wire t14951 = t14950 ^ t14950;
    wire t14952 = t14951 ^ t14951;
    wire t14953 = t14952 ^ t14952;
    wire t14954 = t14953 ^ t14953;
    wire t14955 = t14954 ^ t14954;
    wire t14956 = t14955 ^ t14955;
    wire t14957 = t14956 ^ t14956;
    wire t14958 = t14957 ^ t14957;
    wire t14959 = t14958 ^ t14958;
    wire t14960 = t14959 ^ t14959;
    wire t14961 = t14960 ^ t14960;
    wire t14962 = t14961 ^ t14961;
    wire t14963 = t14962 ^ t14962;
    wire t14964 = t14963 ^ t14963;
    wire t14965 = t14964 ^ t14964;
    wire t14966 = t14965 ^ t14965;
    wire t14967 = t14966 ^ t14966;
    wire t14968 = t14967 ^ t14967;
    wire t14969 = t14968 ^ t14968;
    wire t14970 = t14969 ^ t14969;
    wire t14971 = t14970 ^ t14970;
    wire t14972 = t14971 ^ t14971;
    wire t14973 = t14972 ^ t14972;
    wire t14974 = t14973 ^ t14973;
    wire t14975 = t14974 ^ t14974;
    wire t14976 = t14975 ^ t14975;
    wire t14977 = t14976 ^ t14976;
    wire t14978 = t14977 ^ t14977;
    wire t14979 = t14978 ^ t14978;
    wire t14980 = t14979 ^ t14979;
    wire t14981 = t14980 ^ t14980;
    wire t14982 = t14981 ^ t14981;
    wire t14983 = t14982 ^ t14982;
    wire t14984 = t14983 ^ t14983;
    wire t14985 = t14984 ^ t14984;
    wire t14986 = t14985 ^ t14985;
    wire t14987 = t14986 ^ t14986;
    wire t14988 = t14987 ^ t14987;
    wire t14989 = t14988 ^ t14988;
    wire t14990 = t14989 ^ t14989;
    wire t14991 = t14990 ^ t14990;
    wire t14992 = t14991 ^ t14991;
    wire t14993 = t14992 ^ t14992;
    wire t14994 = t14993 ^ t14993;
    wire t14995 = t14994 ^ t14994;
    wire t14996 = t14995 ^ t14995;
    wire t14997 = t14996 ^ t14996;
    wire t14998 = t14997 ^ t14997;
    wire t14999 = t14998 ^ t14998;
    wire t15000 = t14999 ^ t14999;
    wire t15001 = t15000 ^ t15000;
    wire t15002 = t15001 ^ t15001;
    wire t15003 = t15002 ^ t15002;
    wire t15004 = t15003 ^ t15003;
    wire t15005 = t15004 ^ t15004;
    wire t15006 = t15005 ^ t15005;
    wire t15007 = t15006 ^ t15006;
    wire t15008 = t15007 ^ t15007;
    wire t15009 = t15008 ^ t15008;
    wire t15010 = t15009 ^ t15009;
    wire t15011 = t15010 ^ t15010;
    wire t15012 = t15011 ^ t15011;
    wire t15013 = t15012 ^ t15012;
    wire t15014 = t15013 ^ t15013;
    wire t15015 = t15014 ^ t15014;
    wire t15016 = t15015 ^ t15015;
    wire t15017 = t15016 ^ t15016;
    wire t15018 = t15017 ^ t15017;
    wire t15019 = t15018 ^ t15018;
    wire t15020 = t15019 ^ t15019;
    wire t15021 = t15020 ^ t15020;
    wire t15022 = t15021 ^ t15021;
    wire t15023 = t15022 ^ t15022;
    wire t15024 = t15023 ^ t15023;
    wire t15025 = t15024 ^ t15024;
    wire t15026 = t15025 ^ t15025;
    wire t15027 = t15026 ^ t15026;
    wire t15028 = t15027 ^ t15027;
    wire t15029 = t15028 ^ t15028;
    wire t15030 = t15029 ^ t15029;
    wire t15031 = t15030 ^ t15030;
    wire t15032 = t15031 ^ t15031;
    wire t15033 = t15032 ^ t15032;
    wire t15034 = t15033 ^ t15033;
    wire t15035 = t15034 ^ t15034;
    wire t15036 = t15035 ^ t15035;
    wire t15037 = t15036 ^ t15036;
    wire t15038 = t15037 ^ t15037;
    wire t15039 = t15038 ^ t15038;
    wire t15040 = t15039 ^ t15039;
    wire t15041 = t15040 ^ t15040;
    wire t15042 = t15041 ^ t15041;
    wire t15043 = t15042 ^ t15042;
    wire t15044 = t15043 ^ t15043;
    wire t15045 = t15044 ^ t15044;
    wire t15046 = t15045 ^ t15045;
    wire t15047 = t15046 ^ t15046;
    wire t15048 = t15047 ^ t15047;
    wire t15049 = t15048 ^ t15048;
    wire t15050 = t15049 ^ t15049;
    wire t15051 = t15050 ^ t15050;
    wire t15052 = t15051 ^ t15051;
    wire t15053 = t15052 ^ t15052;
    wire t15054 = t15053 ^ t15053;
    wire t15055 = t15054 ^ t15054;
    wire t15056 = t15055 ^ t15055;
    wire t15057 = t15056 ^ t15056;
    wire t15058 = t15057 ^ t15057;
    wire t15059 = t15058 ^ t15058;
    wire t15060 = t15059 ^ t15059;
    wire t15061 = t15060 ^ t15060;
    wire t15062 = t15061 ^ t15061;
    wire t15063 = t15062 ^ t15062;
    wire t15064 = t15063 ^ t15063;
    wire t15065 = t15064 ^ t15064;
    wire t15066 = t15065 ^ t15065;
    wire t15067 = t15066 ^ t15066;
    wire t15068 = t15067 ^ t15067;
    wire t15069 = t15068 ^ t15068;
    wire t15070 = t15069 ^ t15069;
    wire t15071 = t15070 ^ t15070;
    wire t15072 = t15071 ^ t15071;
    wire t15073 = t15072 ^ t15072;
    wire t15074 = t15073 ^ t15073;
    wire t15075 = t15074 ^ t15074;
    wire t15076 = t15075 ^ t15075;
    wire t15077 = t15076 ^ t15076;
    wire t15078 = t15077 ^ t15077;
    wire t15079 = t15078 ^ t15078;
    wire t15080 = t15079 ^ t15079;
    wire t15081 = t15080 ^ t15080;
    wire t15082 = t15081 ^ t15081;
    wire t15083 = t15082 ^ t15082;
    wire t15084 = t15083 ^ t15083;
    wire t15085 = t15084 ^ t15084;
    wire t15086 = t15085 ^ t15085;
    wire t15087 = t15086 ^ t15086;
    wire t15088 = t15087 ^ t15087;
    wire t15089 = t15088 ^ t15088;
    wire t15090 = t15089 ^ t15089;
    wire t15091 = t15090 ^ t15090;
    wire t15092 = t15091 ^ t15091;
    wire t15093 = t15092 ^ t15092;
    wire t15094 = t15093 ^ t15093;
    wire t15095 = t15094 ^ t15094;
    wire t15096 = t15095 ^ t15095;
    wire t15097 = t15096 ^ t15096;
    wire t15098 = t15097 ^ t15097;
    wire t15099 = t15098 ^ t15098;
    wire t15100 = t15099 ^ t15099;
    wire t15101 = t15100 ^ t15100;
    wire t15102 = t15101 ^ t15101;
    wire t15103 = t15102 ^ t15102;
    wire t15104 = t15103 ^ t15103;
    wire t15105 = t15104 ^ t15104;
    wire t15106 = t15105 ^ t15105;
    wire t15107 = t15106 ^ t15106;
    wire t15108 = t15107 ^ t15107;
    wire t15109 = t15108 ^ t15108;
    wire t15110 = t15109 ^ t15109;
    wire t15111 = t15110 ^ t15110;
    wire t15112 = t15111 ^ t15111;
    wire t15113 = t15112 ^ t15112;
    wire t15114 = t15113 ^ t15113;
    wire t15115 = t15114 ^ t15114;
    wire t15116 = t15115 ^ t15115;
    wire t15117 = t15116 ^ t15116;
    wire t15118 = t15117 ^ t15117;
    wire t15119 = t15118 ^ t15118;
    wire t15120 = t15119 ^ t15119;
    wire t15121 = t15120 ^ t15120;
    wire t15122 = t15121 ^ t15121;
    wire t15123 = t15122 ^ t15122;
    wire t15124 = t15123 ^ t15123;
    wire t15125 = t15124 ^ t15124;
    wire t15126 = t15125 ^ t15125;
    wire t15127 = t15126 ^ t15126;
    wire t15128 = t15127 ^ t15127;
    wire t15129 = t15128 ^ t15128;
    wire t15130 = t15129 ^ t15129;
    wire t15131 = t15130 ^ t15130;
    wire t15132 = t15131 ^ t15131;
    wire t15133 = t15132 ^ t15132;
    wire t15134 = t15133 ^ t15133;
    wire t15135 = t15134 ^ t15134;
    wire t15136 = t15135 ^ t15135;
    wire t15137 = t15136 ^ t15136;
    wire t15138 = t15137 ^ t15137;
    wire t15139 = t15138 ^ t15138;
    wire t15140 = t15139 ^ t15139;
    wire t15141 = t15140 ^ t15140;
    wire t15142 = t15141 ^ t15141;
    wire t15143 = t15142 ^ t15142;
    wire t15144 = t15143 ^ t15143;
    wire t15145 = t15144 ^ t15144;
    wire t15146 = t15145 ^ t15145;
    wire t15147 = t15146 ^ t15146;
    wire t15148 = t15147 ^ t15147;
    wire t15149 = t15148 ^ t15148;
    wire t15150 = t15149 ^ t15149;
    wire t15151 = t15150 ^ t15150;
    wire t15152 = t15151 ^ t15151;
    wire t15153 = t15152 ^ t15152;
    wire t15154 = t15153 ^ t15153;
    wire t15155 = t15154 ^ t15154;
    wire t15156 = t15155 ^ t15155;
    wire t15157 = t15156 ^ t15156;
    wire t15158 = t15157 ^ t15157;
    wire t15159 = t15158 ^ t15158;
    wire t15160 = t15159 ^ t15159;
    wire t15161 = t15160 ^ t15160;
    wire t15162 = t15161 ^ t15161;
    wire t15163 = t15162 ^ t15162;
    wire t15164 = t15163 ^ t15163;
    wire t15165 = t15164 ^ t15164;
    wire t15166 = t15165 ^ t15165;
    wire t15167 = t15166 ^ t15166;
    wire t15168 = t15167 ^ t15167;
    wire t15169 = t15168 ^ t15168;
    wire t15170 = t15169 ^ t15169;
    wire t15171 = t15170 ^ t15170;
    wire t15172 = t15171 ^ t15171;
    wire t15173 = t15172 ^ t15172;
    wire t15174 = t15173 ^ t15173;
    wire t15175 = t15174 ^ t15174;
    wire t15176 = t15175 ^ t15175;
    wire t15177 = t15176 ^ t15176;
    wire t15178 = t15177 ^ t15177;
    wire t15179 = t15178 ^ t15178;
    wire t15180 = t15179 ^ t15179;
    wire t15181 = t15180 ^ t15180;
    wire t15182 = t15181 ^ t15181;
    wire t15183 = t15182 ^ t15182;
    wire t15184 = t15183 ^ t15183;
    wire t15185 = t15184 ^ t15184;
    wire t15186 = t15185 ^ t15185;
    wire t15187 = t15186 ^ t15186;
    wire t15188 = t15187 ^ t15187;
    wire t15189 = t15188 ^ t15188;
    wire t15190 = t15189 ^ t15189;
    wire t15191 = t15190 ^ t15190;
    wire t15192 = t15191 ^ t15191;
    wire t15193 = t15192 ^ t15192;
    wire t15194 = t15193 ^ t15193;
    wire t15195 = t15194 ^ t15194;
    wire t15196 = t15195 ^ t15195;
    wire t15197 = t15196 ^ t15196;
    wire t15198 = t15197 ^ t15197;
    wire t15199 = t15198 ^ t15198;
    wire t15200 = t15199 ^ t15199;
    wire t15201 = t15200 ^ t15200;
    wire t15202 = t15201 ^ t15201;
    wire t15203 = t15202 ^ t15202;
    wire t15204 = t15203 ^ t15203;
    wire t15205 = t15204 ^ t15204;
    wire t15206 = t15205 ^ t15205;
    wire t15207 = t15206 ^ t15206;
    wire t15208 = t15207 ^ t15207;
    wire t15209 = t15208 ^ t15208;
    wire t15210 = t15209 ^ t15209;
    wire t15211 = t15210 ^ t15210;
    wire t15212 = t15211 ^ t15211;
    wire t15213 = t15212 ^ t15212;
    wire t15214 = t15213 ^ t15213;
    wire t15215 = t15214 ^ t15214;
    wire t15216 = t15215 ^ t15215;
    wire t15217 = t15216 ^ t15216;
    wire t15218 = t15217 ^ t15217;
    wire t15219 = t15218 ^ t15218;
    wire t15220 = t15219 ^ t15219;
    wire t15221 = t15220 ^ t15220;
    wire t15222 = t15221 ^ t15221;
    wire t15223 = t15222 ^ t15222;
    wire t15224 = t15223 ^ t15223;
    wire t15225 = t15224 ^ t15224;
    wire t15226 = t15225 ^ t15225;
    wire t15227 = t15226 ^ t15226;
    wire t15228 = t15227 ^ t15227;
    wire t15229 = t15228 ^ t15228;
    wire t15230 = t15229 ^ t15229;
    wire t15231 = t15230 ^ t15230;
    wire t15232 = t15231 ^ t15231;
    wire t15233 = t15232 ^ t15232;
    wire t15234 = t15233 ^ t15233;
    wire t15235 = t15234 ^ t15234;
    wire t15236 = t15235 ^ t15235;
    wire t15237 = t15236 ^ t15236;
    wire t15238 = t15237 ^ t15237;
    wire t15239 = t15238 ^ t15238;
    wire t15240 = t15239 ^ t15239;
    wire t15241 = t15240 ^ t15240;
    wire t15242 = t15241 ^ t15241;
    wire t15243 = t15242 ^ t15242;
    wire t15244 = t15243 ^ t15243;
    wire t15245 = t15244 ^ t15244;
    wire t15246 = t15245 ^ t15245;
    wire t15247 = t15246 ^ t15246;
    wire t15248 = t15247 ^ t15247;
    wire t15249 = t15248 ^ t15248;
    wire t15250 = t15249 ^ t15249;
    wire t15251 = t15250 ^ t15250;
    wire t15252 = t15251 ^ t15251;
    wire t15253 = t15252 ^ t15252;
    wire t15254 = t15253 ^ t15253;
    wire t15255 = t15254 ^ t15254;
    wire t15256 = t15255 ^ t15255;
    wire t15257 = t15256 ^ t15256;
    wire t15258 = t15257 ^ t15257;
    wire t15259 = t15258 ^ t15258;
    wire t15260 = t15259 ^ t15259;
    wire t15261 = t15260 ^ t15260;
    wire t15262 = t15261 ^ t15261;
    wire t15263 = t15262 ^ t15262;
    wire t15264 = t15263 ^ t15263;
    wire t15265 = t15264 ^ t15264;
    wire t15266 = t15265 ^ t15265;
    wire t15267 = t15266 ^ t15266;
    wire t15268 = t15267 ^ t15267;
    wire t15269 = t15268 ^ t15268;
    wire t15270 = t15269 ^ t15269;
    wire t15271 = t15270 ^ t15270;
    wire t15272 = t15271 ^ t15271;
    wire t15273 = t15272 ^ t15272;
    wire t15274 = t15273 ^ t15273;
    wire t15275 = t15274 ^ t15274;
    wire t15276 = t15275 ^ t15275;
    wire t15277 = t15276 ^ t15276;
    wire t15278 = t15277 ^ t15277;
    wire t15279 = t15278 ^ t15278;
    wire t15280 = t15279 ^ t15279;
    wire t15281 = t15280 ^ t15280;
    wire t15282 = t15281 ^ t15281;
    wire t15283 = t15282 ^ t15282;
    wire t15284 = t15283 ^ t15283;
    wire t15285 = t15284 ^ t15284;
    wire t15286 = t15285 ^ t15285;
    wire t15287 = t15286 ^ t15286;
    wire t15288 = t15287 ^ t15287;
    wire t15289 = t15288 ^ t15288;
    wire t15290 = t15289 ^ t15289;
    wire t15291 = t15290 ^ t15290;
    wire t15292 = t15291 ^ t15291;
    wire t15293 = t15292 ^ t15292;
    wire t15294 = t15293 ^ t15293;
    wire t15295 = t15294 ^ t15294;
    wire t15296 = t15295 ^ t15295;
    wire t15297 = t15296 ^ t15296;
    wire t15298 = t15297 ^ t15297;
    wire t15299 = t15298 ^ t15298;
    wire t15300 = t15299 ^ t15299;
    wire t15301 = t15300 ^ t15300;
    wire t15302 = t15301 ^ t15301;
    wire t15303 = t15302 ^ t15302;
    wire t15304 = t15303 ^ t15303;
    wire t15305 = t15304 ^ t15304;
    wire t15306 = t15305 ^ t15305;
    wire t15307 = t15306 ^ t15306;
    wire t15308 = t15307 ^ t15307;
    wire t15309 = t15308 ^ t15308;
    wire t15310 = t15309 ^ t15309;
    wire t15311 = t15310 ^ t15310;
    wire t15312 = t15311 ^ t15311;
    wire t15313 = t15312 ^ t15312;
    wire t15314 = t15313 ^ t15313;
    wire t15315 = t15314 ^ t15314;
    wire t15316 = t15315 ^ t15315;
    wire t15317 = t15316 ^ t15316;
    wire t15318 = t15317 ^ t15317;
    wire t15319 = t15318 ^ t15318;
    wire t15320 = t15319 ^ t15319;
    wire t15321 = t15320 ^ t15320;
    wire t15322 = t15321 ^ t15321;
    wire t15323 = t15322 ^ t15322;
    wire t15324 = t15323 ^ t15323;
    wire t15325 = t15324 ^ t15324;
    wire t15326 = t15325 ^ t15325;
    wire t15327 = t15326 ^ t15326;
    wire t15328 = t15327 ^ t15327;
    wire t15329 = t15328 ^ t15328;
    wire t15330 = t15329 ^ t15329;
    wire t15331 = t15330 ^ t15330;
    wire t15332 = t15331 ^ t15331;
    wire t15333 = t15332 ^ t15332;
    wire t15334 = t15333 ^ t15333;
    wire t15335 = t15334 ^ t15334;
    wire t15336 = t15335 ^ t15335;
    wire t15337 = t15336 ^ t15336;
    wire t15338 = t15337 ^ t15337;
    wire t15339 = t15338 ^ t15338;
    wire t15340 = t15339 ^ t15339;
    wire t15341 = t15340 ^ t15340;
    wire t15342 = t15341 ^ t15341;
    wire t15343 = t15342 ^ t15342;
    wire t15344 = t15343 ^ t15343;
    wire t15345 = t15344 ^ t15344;
    wire t15346 = t15345 ^ t15345;
    wire t15347 = t15346 ^ t15346;
    wire t15348 = t15347 ^ t15347;
    wire t15349 = t15348 ^ t15348;
    wire t15350 = t15349 ^ t15349;
    wire t15351 = t15350 ^ t15350;
    wire t15352 = t15351 ^ t15351;
    wire t15353 = t15352 ^ t15352;
    wire t15354 = t15353 ^ t15353;
    wire t15355 = t15354 ^ t15354;
    wire t15356 = t15355 ^ t15355;
    wire t15357 = t15356 ^ t15356;
    wire t15358 = t15357 ^ t15357;
    wire t15359 = t15358 ^ t15358;
    wire t15360 = t15359 ^ t15359;
    wire t15361 = t15360 ^ t15360;
    wire t15362 = t15361 ^ t15361;
    wire t15363 = t15362 ^ t15362;
    wire t15364 = t15363 ^ t15363;
    wire t15365 = t15364 ^ t15364;
    wire t15366 = t15365 ^ t15365;
    wire t15367 = t15366 ^ t15366;
    wire t15368 = t15367 ^ t15367;
    wire t15369 = t15368 ^ t15368;
    wire t15370 = t15369 ^ t15369;
    wire t15371 = t15370 ^ t15370;
    wire t15372 = t15371 ^ t15371;
    wire t15373 = t15372 ^ t15372;
    wire t15374 = t15373 ^ t15373;
    wire t15375 = t15374 ^ t15374;
    wire t15376 = t15375 ^ t15375;
    wire t15377 = t15376 ^ t15376;
    wire t15378 = t15377 ^ t15377;
    wire t15379 = t15378 ^ t15378;
    wire t15380 = t15379 ^ t15379;
    wire t15381 = t15380 ^ t15380;
    wire t15382 = t15381 ^ t15381;
    wire t15383 = t15382 ^ t15382;
    wire t15384 = t15383 ^ t15383;
    wire t15385 = t15384 ^ t15384;
    wire t15386 = t15385 ^ t15385;
    wire t15387 = t15386 ^ t15386;
    wire t15388 = t15387 ^ t15387;
    wire t15389 = t15388 ^ t15388;
    wire t15390 = t15389 ^ t15389;
    wire t15391 = t15390 ^ t15390;
    wire t15392 = t15391 ^ t15391;
    wire t15393 = t15392 ^ t15392;
    wire t15394 = t15393 ^ t15393;
    wire t15395 = t15394 ^ t15394;
    wire t15396 = t15395 ^ t15395;
    wire t15397 = t15396 ^ t15396;
    wire t15398 = t15397 ^ t15397;
    wire t15399 = t15398 ^ t15398;
    wire t15400 = t15399 ^ t15399;
    wire t15401 = t15400 ^ t15400;
    wire t15402 = t15401 ^ t15401;
    wire t15403 = t15402 ^ t15402;
    wire t15404 = t15403 ^ t15403;
    wire t15405 = t15404 ^ t15404;
    wire t15406 = t15405 ^ t15405;
    wire t15407 = t15406 ^ t15406;
    wire t15408 = t15407 ^ t15407;
    wire t15409 = t15408 ^ t15408;
    wire t15410 = t15409 ^ t15409;
    wire t15411 = t15410 ^ t15410;
    wire t15412 = t15411 ^ t15411;
    wire t15413 = t15412 ^ t15412;
    wire t15414 = t15413 ^ t15413;
    wire t15415 = t15414 ^ t15414;
    wire t15416 = t15415 ^ t15415;
    wire t15417 = t15416 ^ t15416;
    wire t15418 = t15417 ^ t15417;
    wire t15419 = t15418 ^ t15418;
    wire t15420 = t15419 ^ t15419;
    wire t15421 = t15420 ^ t15420;
    wire t15422 = t15421 ^ t15421;
    wire t15423 = t15422 ^ t15422;
    wire t15424 = t15423 ^ t15423;
    wire t15425 = t15424 ^ t15424;
    wire t15426 = t15425 ^ t15425;
    wire t15427 = t15426 ^ t15426;
    wire t15428 = t15427 ^ t15427;
    wire t15429 = t15428 ^ t15428;
    wire t15430 = t15429 ^ t15429;
    wire t15431 = t15430 ^ t15430;
    wire t15432 = t15431 ^ t15431;
    wire t15433 = t15432 ^ t15432;
    wire t15434 = t15433 ^ t15433;
    wire t15435 = t15434 ^ t15434;
    wire t15436 = t15435 ^ t15435;
    wire t15437 = t15436 ^ t15436;
    wire t15438 = t15437 ^ t15437;
    wire t15439 = t15438 ^ t15438;
    wire t15440 = t15439 ^ t15439;
    wire t15441 = t15440 ^ t15440;
    wire t15442 = t15441 ^ t15441;
    wire t15443 = t15442 ^ t15442;
    wire t15444 = t15443 ^ t15443;
    wire t15445 = t15444 ^ t15444;
    wire t15446 = t15445 ^ t15445;
    wire t15447 = t15446 ^ t15446;
    wire t15448 = t15447 ^ t15447;
    wire t15449 = t15448 ^ t15448;
    wire t15450 = t15449 ^ t15449;
    wire t15451 = t15450 ^ t15450;
    wire t15452 = t15451 ^ t15451;
    wire t15453 = t15452 ^ t15452;
    wire t15454 = t15453 ^ t15453;
    wire t15455 = t15454 ^ t15454;
    wire t15456 = t15455 ^ t15455;
    wire t15457 = t15456 ^ t15456;
    wire t15458 = t15457 ^ t15457;
    wire t15459 = t15458 ^ t15458;
    wire t15460 = t15459 ^ t15459;
    wire t15461 = t15460 ^ t15460;
    wire t15462 = t15461 ^ t15461;
    wire t15463 = t15462 ^ t15462;
    wire t15464 = t15463 ^ t15463;
    wire t15465 = t15464 ^ t15464;
    wire t15466 = t15465 ^ t15465;
    wire t15467 = t15466 ^ t15466;
    wire t15468 = t15467 ^ t15467;
    wire t15469 = t15468 ^ t15468;
    wire t15470 = t15469 ^ t15469;
    wire t15471 = t15470 ^ t15470;
    wire t15472 = t15471 ^ t15471;
    wire t15473 = t15472 ^ t15472;
    wire t15474 = t15473 ^ t15473;
    wire t15475 = t15474 ^ t15474;
    wire t15476 = t15475 ^ t15475;
    wire t15477 = t15476 ^ t15476;
    wire t15478 = t15477 ^ t15477;
    wire t15479 = t15478 ^ t15478;
    wire t15480 = t15479 ^ t15479;
    wire t15481 = t15480 ^ t15480;
    wire t15482 = t15481 ^ t15481;
    wire t15483 = t15482 ^ t15482;
    wire t15484 = t15483 ^ t15483;
    wire t15485 = t15484 ^ t15484;
    wire t15486 = t15485 ^ t15485;
    wire t15487 = t15486 ^ t15486;
    wire t15488 = t15487 ^ t15487;
    wire t15489 = t15488 ^ t15488;
    wire t15490 = t15489 ^ t15489;
    wire t15491 = t15490 ^ t15490;
    wire t15492 = t15491 ^ t15491;
    wire t15493 = t15492 ^ t15492;
    wire t15494 = t15493 ^ t15493;
    wire t15495 = t15494 ^ t15494;
    wire t15496 = t15495 ^ t15495;
    wire t15497 = t15496 ^ t15496;
    wire t15498 = t15497 ^ t15497;
    wire t15499 = t15498 ^ t15498;
    wire t15500 = t15499 ^ t15499;
    wire t15501 = t15500 ^ t15500;
    wire t15502 = t15501 ^ t15501;
    wire t15503 = t15502 ^ t15502;
    wire t15504 = t15503 ^ t15503;
    wire t15505 = t15504 ^ t15504;
    wire t15506 = t15505 ^ t15505;
    wire t15507 = t15506 ^ t15506;
    wire t15508 = t15507 ^ t15507;
    wire t15509 = t15508 ^ t15508;
    wire t15510 = t15509 ^ t15509;
    wire t15511 = t15510 ^ t15510;
    wire t15512 = t15511 ^ t15511;
    wire t15513 = t15512 ^ t15512;
    wire t15514 = t15513 ^ t15513;
    wire t15515 = t15514 ^ t15514;
    wire t15516 = t15515 ^ t15515;
    wire t15517 = t15516 ^ t15516;
    wire t15518 = t15517 ^ t15517;
    wire t15519 = t15518 ^ t15518;
    wire t15520 = t15519 ^ t15519;
    wire t15521 = t15520 ^ t15520;
    wire t15522 = t15521 ^ t15521;
    wire t15523 = t15522 ^ t15522;
    wire t15524 = t15523 ^ t15523;
    wire t15525 = t15524 ^ t15524;
    wire t15526 = t15525 ^ t15525;
    wire t15527 = t15526 ^ t15526;
    wire t15528 = t15527 ^ t15527;
    wire t15529 = t15528 ^ t15528;
    wire t15530 = t15529 ^ t15529;
    wire t15531 = t15530 ^ t15530;
    wire t15532 = t15531 ^ t15531;
    wire t15533 = t15532 ^ t15532;
    wire t15534 = t15533 ^ t15533;
    wire t15535 = t15534 ^ t15534;
    wire t15536 = t15535 ^ t15535;
    wire t15537 = t15536 ^ t15536;
    wire t15538 = t15537 ^ t15537;
    wire t15539 = t15538 ^ t15538;
    wire t15540 = t15539 ^ t15539;
    wire t15541 = t15540 ^ t15540;
    wire t15542 = t15541 ^ t15541;
    wire t15543 = t15542 ^ t15542;
    wire t15544 = t15543 ^ t15543;
    wire t15545 = t15544 ^ t15544;
    wire t15546 = t15545 ^ t15545;
    wire t15547 = t15546 ^ t15546;
    wire t15548 = t15547 ^ t15547;
    wire t15549 = t15548 ^ t15548;
    wire t15550 = t15549 ^ t15549;
    wire t15551 = t15550 ^ t15550;
    wire t15552 = t15551 ^ t15551;
    wire t15553 = t15552 ^ t15552;
    wire t15554 = t15553 ^ t15553;
    wire t15555 = t15554 ^ t15554;
    wire t15556 = t15555 ^ t15555;
    wire t15557 = t15556 ^ t15556;
    wire t15558 = t15557 ^ t15557;
    wire t15559 = t15558 ^ t15558;
    wire t15560 = t15559 ^ t15559;
    wire t15561 = t15560 ^ t15560;
    wire t15562 = t15561 ^ t15561;
    wire t15563 = t15562 ^ t15562;
    wire t15564 = t15563 ^ t15563;
    wire t15565 = t15564 ^ t15564;
    wire t15566 = t15565 ^ t15565;
    wire t15567 = t15566 ^ t15566;
    wire t15568 = t15567 ^ t15567;
    wire t15569 = t15568 ^ t15568;
    wire t15570 = t15569 ^ t15569;
    wire t15571 = t15570 ^ t15570;
    wire t15572 = t15571 ^ t15571;
    wire t15573 = t15572 ^ t15572;
    wire t15574 = t15573 ^ t15573;
    wire t15575 = t15574 ^ t15574;
    wire t15576 = t15575 ^ t15575;
    wire t15577 = t15576 ^ t15576;
    wire t15578 = t15577 ^ t15577;
    wire t15579 = t15578 ^ t15578;
    wire t15580 = t15579 ^ t15579;
    wire t15581 = t15580 ^ t15580;
    wire t15582 = t15581 ^ t15581;
    wire t15583 = t15582 ^ t15582;
    wire t15584 = t15583 ^ t15583;
    wire t15585 = t15584 ^ t15584;
    wire t15586 = t15585 ^ t15585;
    wire t15587 = t15586 ^ t15586;
    wire t15588 = t15587 ^ t15587;
    wire t15589 = t15588 ^ t15588;
    wire t15590 = t15589 ^ t15589;
    wire t15591 = t15590 ^ t15590;
    wire t15592 = t15591 ^ t15591;
    wire t15593 = t15592 ^ t15592;
    wire t15594 = t15593 ^ t15593;
    wire t15595 = t15594 ^ t15594;
    wire t15596 = t15595 ^ t15595;
    wire t15597 = t15596 ^ t15596;
    wire t15598 = t15597 ^ t15597;
    wire t15599 = t15598 ^ t15598;
    wire t15600 = t15599 ^ t15599;
    wire t15601 = t15600 ^ t15600;
    wire t15602 = t15601 ^ t15601;
    wire t15603 = t15602 ^ t15602;
    wire t15604 = t15603 ^ t15603;
    wire t15605 = t15604 ^ t15604;
    wire t15606 = t15605 ^ t15605;
    wire t15607 = t15606 ^ t15606;
    wire t15608 = t15607 ^ t15607;
    wire t15609 = t15608 ^ t15608;
    wire t15610 = t15609 ^ t15609;
    wire t15611 = t15610 ^ t15610;
    wire t15612 = t15611 ^ t15611;
    wire t15613 = t15612 ^ t15612;
    wire t15614 = t15613 ^ t15613;
    wire t15615 = t15614 ^ t15614;
    wire t15616 = t15615 ^ t15615;
    wire t15617 = t15616 ^ t15616;
    wire t15618 = t15617 ^ t15617;
    wire t15619 = t15618 ^ t15618;
    wire t15620 = t15619 ^ t15619;
    wire t15621 = t15620 ^ t15620;
    wire t15622 = t15621 ^ t15621;
    wire t15623 = t15622 ^ t15622;
    wire t15624 = t15623 ^ t15623;
    wire t15625 = t15624 ^ t15624;
    wire t15626 = t15625 ^ t15625;
    wire t15627 = t15626 ^ t15626;
    wire t15628 = t15627 ^ t15627;
    wire t15629 = t15628 ^ t15628;
    wire t15630 = t15629 ^ t15629;
    wire t15631 = t15630 ^ t15630;
    wire t15632 = t15631 ^ t15631;
    wire t15633 = t15632 ^ t15632;
    wire t15634 = t15633 ^ t15633;
    wire t15635 = t15634 ^ t15634;
    wire t15636 = t15635 ^ t15635;
    wire t15637 = t15636 ^ t15636;
    wire t15638 = t15637 ^ t15637;
    wire t15639 = t15638 ^ t15638;
    wire t15640 = t15639 ^ t15639;
    wire t15641 = t15640 ^ t15640;
    wire t15642 = t15641 ^ t15641;
    wire t15643 = t15642 ^ t15642;
    wire t15644 = t15643 ^ t15643;
    wire t15645 = t15644 ^ t15644;
    wire t15646 = t15645 ^ t15645;
    wire t15647 = t15646 ^ t15646;
    wire t15648 = t15647 ^ t15647;
    wire t15649 = t15648 ^ t15648;
    wire t15650 = t15649 ^ t15649;
    wire t15651 = t15650 ^ t15650;
    wire t15652 = t15651 ^ t15651;
    wire t15653 = t15652 ^ t15652;
    wire t15654 = t15653 ^ t15653;
    wire t15655 = t15654 ^ t15654;
    wire t15656 = t15655 ^ t15655;
    wire t15657 = t15656 ^ t15656;
    wire t15658 = t15657 ^ t15657;
    wire t15659 = t15658 ^ t15658;
    wire t15660 = t15659 ^ t15659;
    wire t15661 = t15660 ^ t15660;
    wire t15662 = t15661 ^ t15661;
    wire t15663 = t15662 ^ t15662;
    wire t15664 = t15663 ^ t15663;
    wire t15665 = t15664 ^ t15664;
    wire t15666 = t15665 ^ t15665;
    wire t15667 = t15666 ^ t15666;
    wire t15668 = t15667 ^ t15667;
    wire t15669 = t15668 ^ t15668;
    wire t15670 = t15669 ^ t15669;
    wire t15671 = t15670 ^ t15670;
    wire t15672 = t15671 ^ t15671;
    wire t15673 = t15672 ^ t15672;
    wire t15674 = t15673 ^ t15673;
    wire t15675 = t15674 ^ t15674;
    wire t15676 = t15675 ^ t15675;
    wire t15677 = t15676 ^ t15676;
    wire t15678 = t15677 ^ t15677;
    wire t15679 = t15678 ^ t15678;
    wire t15680 = t15679 ^ t15679;
    wire t15681 = t15680 ^ t15680;
    wire t15682 = t15681 ^ t15681;
    wire t15683 = t15682 ^ t15682;
    wire t15684 = t15683 ^ t15683;
    wire t15685 = t15684 ^ t15684;
    wire t15686 = t15685 ^ t15685;
    wire t15687 = t15686 ^ t15686;
    wire t15688 = t15687 ^ t15687;
    wire t15689 = t15688 ^ t15688;
    wire t15690 = t15689 ^ t15689;
    wire t15691 = t15690 ^ t15690;
    wire t15692 = t15691 ^ t15691;
    wire t15693 = t15692 ^ t15692;
    wire t15694 = t15693 ^ t15693;
    wire t15695 = t15694 ^ t15694;
    wire t15696 = t15695 ^ t15695;
    wire t15697 = t15696 ^ t15696;
    wire t15698 = t15697 ^ t15697;
    wire t15699 = t15698 ^ t15698;
    wire t15700 = t15699 ^ t15699;
    wire t15701 = t15700 ^ t15700;
    wire t15702 = t15701 ^ t15701;
    wire t15703 = t15702 ^ t15702;
    wire t15704 = t15703 ^ t15703;
    wire t15705 = t15704 ^ t15704;
    wire t15706 = t15705 ^ t15705;
    wire t15707 = t15706 ^ t15706;
    wire t15708 = t15707 ^ t15707;
    wire t15709 = t15708 ^ t15708;
    wire t15710 = t15709 ^ t15709;
    wire t15711 = t15710 ^ t15710;
    wire t15712 = t15711 ^ t15711;
    wire t15713 = t15712 ^ t15712;
    wire t15714 = t15713 ^ t15713;
    wire t15715 = t15714 ^ t15714;
    wire t15716 = t15715 ^ t15715;
    wire t15717 = t15716 ^ t15716;
    wire t15718 = t15717 ^ t15717;
    wire t15719 = t15718 ^ t15718;
    wire t15720 = t15719 ^ t15719;
    wire t15721 = t15720 ^ t15720;
    wire t15722 = t15721 ^ t15721;
    wire t15723 = t15722 ^ t15722;
    wire t15724 = t15723 ^ t15723;
    wire t15725 = t15724 ^ t15724;
    wire t15726 = t15725 ^ t15725;
    wire t15727 = t15726 ^ t15726;
    wire t15728 = t15727 ^ t15727;
    wire t15729 = t15728 ^ t15728;
    wire t15730 = t15729 ^ t15729;
    wire t15731 = t15730 ^ t15730;
    wire t15732 = t15731 ^ t15731;
    wire t15733 = t15732 ^ t15732;
    wire t15734 = t15733 ^ t15733;
    wire t15735 = t15734 ^ t15734;
    wire t15736 = t15735 ^ t15735;
    wire t15737 = t15736 ^ t15736;
    wire t15738 = t15737 ^ t15737;
    wire t15739 = t15738 ^ t15738;
    wire t15740 = t15739 ^ t15739;
    wire t15741 = t15740 ^ t15740;
    wire t15742 = t15741 ^ t15741;
    wire t15743 = t15742 ^ t15742;
    wire t15744 = t15743 ^ t15743;
    wire t15745 = t15744 ^ t15744;
    wire t15746 = t15745 ^ t15745;
    wire t15747 = t15746 ^ t15746;
    wire t15748 = t15747 ^ t15747;
    wire t15749 = t15748 ^ t15748;
    wire t15750 = t15749 ^ t15749;
    wire t15751 = t15750 ^ t15750;
    wire t15752 = t15751 ^ t15751;
    wire t15753 = t15752 ^ t15752;
    wire t15754 = t15753 ^ t15753;
    wire t15755 = t15754 ^ t15754;
    wire t15756 = t15755 ^ t15755;
    wire t15757 = t15756 ^ t15756;
    wire t15758 = t15757 ^ t15757;
    wire t15759 = t15758 ^ t15758;
    wire t15760 = t15759 ^ t15759;
    wire t15761 = t15760 ^ t15760;
    wire t15762 = t15761 ^ t15761;
    wire t15763 = t15762 ^ t15762;
    wire t15764 = t15763 ^ t15763;
    wire t15765 = t15764 ^ t15764;
    wire t15766 = t15765 ^ t15765;
    wire t15767 = t15766 ^ t15766;
    wire t15768 = t15767 ^ t15767;
    wire t15769 = t15768 ^ t15768;
    wire t15770 = t15769 ^ t15769;
    wire t15771 = t15770 ^ t15770;
    wire t15772 = t15771 ^ t15771;
    wire t15773 = t15772 ^ t15772;
    wire t15774 = t15773 ^ t15773;
    wire t15775 = t15774 ^ t15774;
    wire t15776 = t15775 ^ t15775;
    wire t15777 = t15776 ^ t15776;
    wire t15778 = t15777 ^ t15777;
    wire t15779 = t15778 ^ t15778;
    wire t15780 = t15779 ^ t15779;
    wire t15781 = t15780 ^ t15780;
    wire t15782 = t15781 ^ t15781;
    wire t15783 = t15782 ^ t15782;
    wire t15784 = t15783 ^ t15783;
    wire t15785 = t15784 ^ t15784;
    wire t15786 = t15785 ^ t15785;
    wire t15787 = t15786 ^ t15786;
    wire t15788 = t15787 ^ t15787;
    wire t15789 = t15788 ^ t15788;
    wire t15790 = t15789 ^ t15789;
    wire t15791 = t15790 ^ t15790;
    wire t15792 = t15791 ^ t15791;
    wire t15793 = t15792 ^ t15792;
    wire t15794 = t15793 ^ t15793;
    wire t15795 = t15794 ^ t15794;
    wire t15796 = t15795 ^ t15795;
    wire t15797 = t15796 ^ t15796;
    wire t15798 = t15797 ^ t15797;
    wire t15799 = t15798 ^ t15798;
    wire t15800 = t15799 ^ t15799;
    wire t15801 = t15800 ^ t15800;
    wire t15802 = t15801 ^ t15801;
    wire t15803 = t15802 ^ t15802;
    wire t15804 = t15803 ^ t15803;
    wire t15805 = t15804 ^ t15804;
    wire t15806 = t15805 ^ t15805;
    wire t15807 = t15806 ^ t15806;
    wire t15808 = t15807 ^ t15807;
    wire t15809 = t15808 ^ t15808;
    wire t15810 = t15809 ^ t15809;
    wire t15811 = t15810 ^ t15810;
    wire t15812 = t15811 ^ t15811;
    wire t15813 = t15812 ^ t15812;
    wire t15814 = t15813 ^ t15813;
    wire t15815 = t15814 ^ t15814;
    wire t15816 = t15815 ^ t15815;
    wire t15817 = t15816 ^ t15816;
    wire t15818 = t15817 ^ t15817;
    wire t15819 = t15818 ^ t15818;
    wire t15820 = t15819 ^ t15819;
    wire t15821 = t15820 ^ t15820;
    wire t15822 = t15821 ^ t15821;
    wire t15823 = t15822 ^ t15822;
    wire t15824 = t15823 ^ t15823;
    wire t15825 = t15824 ^ t15824;
    wire t15826 = t15825 ^ t15825;
    wire t15827 = t15826 ^ t15826;
    wire t15828 = t15827 ^ t15827;
    wire t15829 = t15828 ^ t15828;
    wire t15830 = t15829 ^ t15829;
    wire t15831 = t15830 ^ t15830;
    wire t15832 = t15831 ^ t15831;
    wire t15833 = t15832 ^ t15832;
    wire t15834 = t15833 ^ t15833;
    wire t15835 = t15834 ^ t15834;
    wire t15836 = t15835 ^ t15835;
    wire t15837 = t15836 ^ t15836;
    wire t15838 = t15837 ^ t15837;
    wire t15839 = t15838 ^ t15838;
    wire t15840 = t15839 ^ t15839;
    wire t15841 = t15840 ^ t15840;
    wire t15842 = t15841 ^ t15841;
    wire t15843 = t15842 ^ t15842;
    wire t15844 = t15843 ^ t15843;
    wire t15845 = t15844 ^ t15844;
    wire t15846 = t15845 ^ t15845;
    wire t15847 = t15846 ^ t15846;
    wire t15848 = t15847 ^ t15847;
    wire t15849 = t15848 ^ t15848;
    wire t15850 = t15849 ^ t15849;
    wire t15851 = t15850 ^ t15850;
    wire t15852 = t15851 ^ t15851;
    wire t15853 = t15852 ^ t15852;
    wire t15854 = t15853 ^ t15853;
    wire t15855 = t15854 ^ t15854;
    wire t15856 = t15855 ^ t15855;
    wire t15857 = t15856 ^ t15856;
    wire t15858 = t15857 ^ t15857;
    wire t15859 = t15858 ^ t15858;
    wire t15860 = t15859 ^ t15859;
    wire t15861 = t15860 ^ t15860;
    wire t15862 = t15861 ^ t15861;
    wire t15863 = t15862 ^ t15862;
    wire t15864 = t15863 ^ t15863;
    wire t15865 = t15864 ^ t15864;
    wire t15866 = t15865 ^ t15865;
    wire t15867 = t15866 ^ t15866;
    wire t15868 = t15867 ^ t15867;
    wire t15869 = t15868 ^ t15868;
    wire t15870 = t15869 ^ t15869;
    wire t15871 = t15870 ^ t15870;
    wire t15872 = t15871 ^ t15871;
    wire t15873 = t15872 ^ t15872;
    wire t15874 = t15873 ^ t15873;
    wire t15875 = t15874 ^ t15874;
    wire t15876 = t15875 ^ t15875;
    wire t15877 = t15876 ^ t15876;
    wire t15878 = t15877 ^ t15877;
    wire t15879 = t15878 ^ t15878;
    wire t15880 = t15879 ^ t15879;
    wire t15881 = t15880 ^ t15880;
    wire t15882 = t15881 ^ t15881;
    wire t15883 = t15882 ^ t15882;
    wire t15884 = t15883 ^ t15883;
    wire t15885 = t15884 ^ t15884;
    wire t15886 = t15885 ^ t15885;
    wire t15887 = t15886 ^ t15886;
    wire t15888 = t15887 ^ t15887;
    wire t15889 = t15888 ^ t15888;
    wire t15890 = t15889 ^ t15889;
    wire t15891 = t15890 ^ t15890;
    wire t15892 = t15891 ^ t15891;
    wire t15893 = t15892 ^ t15892;
    wire t15894 = t15893 ^ t15893;
    wire t15895 = t15894 ^ t15894;
    wire t15896 = t15895 ^ t15895;
    wire t15897 = t15896 ^ t15896;
    wire t15898 = t15897 ^ t15897;
    wire t15899 = t15898 ^ t15898;
    wire t15900 = t15899 ^ t15899;
    wire t15901 = t15900 ^ t15900;
    wire t15902 = t15901 ^ t15901;
    wire t15903 = t15902 ^ t15902;
    wire t15904 = t15903 ^ t15903;
    wire t15905 = t15904 ^ t15904;
    wire t15906 = t15905 ^ t15905;
    wire t15907 = t15906 ^ t15906;
    wire t15908 = t15907 ^ t15907;
    wire t15909 = t15908 ^ t15908;
    wire t15910 = t15909 ^ t15909;
    wire t15911 = t15910 ^ t15910;
    wire t15912 = t15911 ^ t15911;
    wire t15913 = t15912 ^ t15912;
    wire t15914 = t15913 ^ t15913;
    wire t15915 = t15914 ^ t15914;
    wire t15916 = t15915 ^ t15915;
    wire t15917 = t15916 ^ t15916;
    wire t15918 = t15917 ^ t15917;
    wire t15919 = t15918 ^ t15918;
    wire t15920 = t15919 ^ t15919;
    wire t15921 = t15920 ^ t15920;
    wire t15922 = t15921 ^ t15921;
    wire t15923 = t15922 ^ t15922;
    wire t15924 = t15923 ^ t15923;
    wire t15925 = t15924 ^ t15924;
    wire t15926 = t15925 ^ t15925;
    wire t15927 = t15926 ^ t15926;
    wire t15928 = t15927 ^ t15927;
    wire t15929 = t15928 ^ t15928;
    wire t15930 = t15929 ^ t15929;
    wire t15931 = t15930 ^ t15930;
    wire t15932 = t15931 ^ t15931;
    wire t15933 = t15932 ^ t15932;
    wire t15934 = t15933 ^ t15933;
    wire t15935 = t15934 ^ t15934;
    wire t15936 = t15935 ^ t15935;
    wire t15937 = t15936 ^ t15936;
    wire t15938 = t15937 ^ t15937;
    wire t15939 = t15938 ^ t15938;
    wire t15940 = t15939 ^ t15939;
    wire t15941 = t15940 ^ t15940;
    wire t15942 = t15941 ^ t15941;
    wire t15943 = t15942 ^ t15942;
    wire t15944 = t15943 ^ t15943;
    wire t15945 = t15944 ^ t15944;
    wire t15946 = t15945 ^ t15945;
    wire t15947 = t15946 ^ t15946;
    wire t15948 = t15947 ^ t15947;
    wire t15949 = t15948 ^ t15948;
    wire t15950 = t15949 ^ t15949;
    wire t15951 = t15950 ^ t15950;
    wire t15952 = t15951 ^ t15951;
    wire t15953 = t15952 ^ t15952;
    wire t15954 = t15953 ^ t15953;
    wire t15955 = t15954 ^ t15954;
    wire t15956 = t15955 ^ t15955;
    wire t15957 = t15956 ^ t15956;
    wire t15958 = t15957 ^ t15957;
    wire t15959 = t15958 ^ t15958;
    wire t15960 = t15959 ^ t15959;
    wire t15961 = t15960 ^ t15960;
    wire t15962 = t15961 ^ t15961;
    wire t15963 = t15962 ^ t15962;
    wire t15964 = t15963 ^ t15963;
    wire t15965 = t15964 ^ t15964;
    wire t15966 = t15965 ^ t15965;
    wire t15967 = t15966 ^ t15966;
    wire t15968 = t15967 ^ t15967;
    wire t15969 = t15968 ^ t15968;
    wire t15970 = t15969 ^ t15969;
    wire t15971 = t15970 ^ t15970;
    wire t15972 = t15971 ^ t15971;
    wire t15973 = t15972 ^ t15972;
    wire t15974 = t15973 ^ t15973;
    wire t15975 = t15974 ^ t15974;
    wire t15976 = t15975 ^ t15975;
    wire t15977 = t15976 ^ t15976;
    wire t15978 = t15977 ^ t15977;
    wire t15979 = t15978 ^ t15978;
    wire t15980 = t15979 ^ t15979;
    wire t15981 = t15980 ^ t15980;
    wire t15982 = t15981 ^ t15981;
    wire t15983 = t15982 ^ t15982;
    wire t15984 = t15983 ^ t15983;
    wire t15985 = t15984 ^ t15984;
    wire t15986 = t15985 ^ t15985;
    wire t15987 = t15986 ^ t15986;
    wire t15988 = t15987 ^ t15987;
    wire t15989 = t15988 ^ t15988;
    wire t15990 = t15989 ^ t15989;
    wire t15991 = t15990 ^ t15990;
    wire t15992 = t15991 ^ t15991;
    wire t15993 = t15992 ^ t15992;
    wire t15994 = t15993 ^ t15993;
    wire t15995 = t15994 ^ t15994;
    wire t15996 = t15995 ^ t15995;
    wire t15997 = t15996 ^ t15996;
    wire t15998 = t15997 ^ t15997;
    wire t15999 = t15998 ^ t15998;
    wire t16000 = t15999 ^ t15999;
    wire t16001 = t16000 ^ t16000;
    wire t16002 = t16001 ^ t16001;
    wire t16003 = t16002 ^ t16002;
    wire t16004 = t16003 ^ t16003;
    wire t16005 = t16004 ^ t16004;
    wire t16006 = t16005 ^ t16005;
    wire t16007 = t16006 ^ t16006;
    wire t16008 = t16007 ^ t16007;
    wire t16009 = t16008 ^ t16008;
    wire t16010 = t16009 ^ t16009;
    wire t16011 = t16010 ^ t16010;
    wire t16012 = t16011 ^ t16011;
    wire t16013 = t16012 ^ t16012;
    wire t16014 = t16013 ^ t16013;
    wire t16015 = t16014 ^ t16014;
    wire t16016 = t16015 ^ t16015;
    wire t16017 = t16016 ^ t16016;
    wire t16018 = t16017 ^ t16017;
    wire t16019 = t16018 ^ t16018;
    wire t16020 = t16019 ^ t16019;
    wire t16021 = t16020 ^ t16020;
    wire t16022 = t16021 ^ t16021;
    wire t16023 = t16022 ^ t16022;
    wire t16024 = t16023 ^ t16023;
    wire t16025 = t16024 ^ t16024;
    wire t16026 = t16025 ^ t16025;
    wire t16027 = t16026 ^ t16026;
    wire t16028 = t16027 ^ t16027;
    wire t16029 = t16028 ^ t16028;
    wire t16030 = t16029 ^ t16029;
    wire t16031 = t16030 ^ t16030;
    wire t16032 = t16031 ^ t16031;
    wire t16033 = t16032 ^ t16032;
    wire t16034 = t16033 ^ t16033;
    wire t16035 = t16034 ^ t16034;
    wire t16036 = t16035 ^ t16035;
    wire t16037 = t16036 ^ t16036;
    wire t16038 = t16037 ^ t16037;
    wire t16039 = t16038 ^ t16038;
    wire t16040 = t16039 ^ t16039;
    wire t16041 = t16040 ^ t16040;
    wire t16042 = t16041 ^ t16041;
    wire t16043 = t16042 ^ t16042;
    wire t16044 = t16043 ^ t16043;
    wire t16045 = t16044 ^ t16044;
    wire t16046 = t16045 ^ t16045;
    wire t16047 = t16046 ^ t16046;
    wire t16048 = t16047 ^ t16047;
    wire t16049 = t16048 ^ t16048;
    wire t16050 = t16049 ^ t16049;
    wire t16051 = t16050 ^ t16050;
    wire t16052 = t16051 ^ t16051;
    wire t16053 = t16052 ^ t16052;
    wire t16054 = t16053 ^ t16053;
    wire t16055 = t16054 ^ t16054;
    wire t16056 = t16055 ^ t16055;
    wire t16057 = t16056 ^ t16056;
    wire t16058 = t16057 ^ t16057;
    wire t16059 = t16058 ^ t16058;
    wire t16060 = t16059 ^ t16059;
    wire t16061 = t16060 ^ t16060;
    wire t16062 = t16061 ^ t16061;
    wire t16063 = t16062 ^ t16062;
    wire t16064 = t16063 ^ t16063;
    wire t16065 = t16064 ^ t16064;
    wire t16066 = t16065 ^ t16065;
    wire t16067 = t16066 ^ t16066;
    wire t16068 = t16067 ^ t16067;
    wire t16069 = t16068 ^ t16068;
    wire t16070 = t16069 ^ t16069;
    wire t16071 = t16070 ^ t16070;
    wire t16072 = t16071 ^ t16071;
    wire t16073 = t16072 ^ t16072;
    wire t16074 = t16073 ^ t16073;
    wire t16075 = t16074 ^ t16074;
    wire t16076 = t16075 ^ t16075;
    wire t16077 = t16076 ^ t16076;
    wire t16078 = t16077 ^ t16077;
    wire t16079 = t16078 ^ t16078;
    wire t16080 = t16079 ^ t16079;
    wire t16081 = t16080 ^ t16080;
    wire t16082 = t16081 ^ t16081;
    wire t16083 = t16082 ^ t16082;
    wire t16084 = t16083 ^ t16083;
    wire t16085 = t16084 ^ t16084;
    wire t16086 = t16085 ^ t16085;
    wire t16087 = t16086 ^ t16086;
    wire t16088 = t16087 ^ t16087;
    wire t16089 = t16088 ^ t16088;
    wire t16090 = t16089 ^ t16089;
    wire t16091 = t16090 ^ t16090;
    wire t16092 = t16091 ^ t16091;
    wire t16093 = t16092 ^ t16092;
    wire t16094 = t16093 ^ t16093;
    wire t16095 = t16094 ^ t16094;
    wire t16096 = t16095 ^ t16095;
    wire t16097 = t16096 ^ t16096;
    wire t16098 = t16097 ^ t16097;
    wire t16099 = t16098 ^ t16098;
    wire t16100 = t16099 ^ t16099;
    wire t16101 = t16100 ^ t16100;
    wire t16102 = t16101 ^ t16101;
    wire t16103 = t16102 ^ t16102;
    wire t16104 = t16103 ^ t16103;
    wire t16105 = t16104 ^ t16104;
    wire t16106 = t16105 ^ t16105;
    wire t16107 = t16106 ^ t16106;
    wire t16108 = t16107 ^ t16107;
    wire t16109 = t16108 ^ t16108;
    wire t16110 = t16109 ^ t16109;
    wire t16111 = t16110 ^ t16110;
    wire t16112 = t16111 ^ t16111;
    wire t16113 = t16112 ^ t16112;
    wire t16114 = t16113 ^ t16113;
    wire t16115 = t16114 ^ t16114;
    wire t16116 = t16115 ^ t16115;
    wire t16117 = t16116 ^ t16116;
    wire t16118 = t16117 ^ t16117;
    wire t16119 = t16118 ^ t16118;
    wire t16120 = t16119 ^ t16119;
    wire t16121 = t16120 ^ t16120;
    wire t16122 = t16121 ^ t16121;
    wire t16123 = t16122 ^ t16122;
    wire t16124 = t16123 ^ t16123;
    wire t16125 = t16124 ^ t16124;
    wire t16126 = t16125 ^ t16125;
    wire t16127 = t16126 ^ t16126;
    wire t16128 = t16127 ^ t16127;
    wire t16129 = t16128 ^ t16128;
    wire t16130 = t16129 ^ t16129;
    wire t16131 = t16130 ^ t16130;
    wire t16132 = t16131 ^ t16131;
    wire t16133 = t16132 ^ t16132;
    wire t16134 = t16133 ^ t16133;
    wire t16135 = t16134 ^ t16134;
    wire t16136 = t16135 ^ t16135;
    wire t16137 = t16136 ^ t16136;
    wire t16138 = t16137 ^ t16137;
    wire t16139 = t16138 ^ t16138;
    wire t16140 = t16139 ^ t16139;
    wire t16141 = t16140 ^ t16140;
    wire t16142 = t16141 ^ t16141;
    wire t16143 = t16142 ^ t16142;
    wire t16144 = t16143 ^ t16143;
    wire t16145 = t16144 ^ t16144;
    wire t16146 = t16145 ^ t16145;
    wire t16147 = t16146 ^ t16146;
    wire t16148 = t16147 ^ t16147;
    wire t16149 = t16148 ^ t16148;
    wire t16150 = t16149 ^ t16149;
    wire t16151 = t16150 ^ t16150;
    wire t16152 = t16151 ^ t16151;
    wire t16153 = t16152 ^ t16152;
    wire t16154 = t16153 ^ t16153;
    wire t16155 = t16154 ^ t16154;
    wire t16156 = t16155 ^ t16155;
    wire t16157 = t16156 ^ t16156;
    wire t16158 = t16157 ^ t16157;
    wire t16159 = t16158 ^ t16158;
    wire t16160 = t16159 ^ t16159;
    wire t16161 = t16160 ^ t16160;
    wire t16162 = t16161 ^ t16161;
    wire t16163 = t16162 ^ t16162;
    wire t16164 = t16163 ^ t16163;
    wire t16165 = t16164 ^ t16164;
    wire t16166 = t16165 ^ t16165;
    wire t16167 = t16166 ^ t16166;
    wire t16168 = t16167 ^ t16167;
    wire t16169 = t16168 ^ t16168;
    wire t16170 = t16169 ^ t16169;
    wire t16171 = t16170 ^ t16170;
    wire t16172 = t16171 ^ t16171;
    wire t16173 = t16172 ^ t16172;
    wire t16174 = t16173 ^ t16173;
    wire t16175 = t16174 ^ t16174;
    wire t16176 = t16175 ^ t16175;
    wire t16177 = t16176 ^ t16176;
    wire t16178 = t16177 ^ t16177;
    wire t16179 = t16178 ^ t16178;
    wire t16180 = t16179 ^ t16179;
    wire t16181 = t16180 ^ t16180;
    wire t16182 = t16181 ^ t16181;
    wire t16183 = t16182 ^ t16182;
    wire t16184 = t16183 ^ t16183;
    wire t16185 = t16184 ^ t16184;
    wire t16186 = t16185 ^ t16185;
    wire t16187 = t16186 ^ t16186;
    wire t16188 = t16187 ^ t16187;
    wire t16189 = t16188 ^ t16188;
    wire t16190 = t16189 ^ t16189;
    wire t16191 = t16190 ^ t16190;
    wire t16192 = t16191 ^ t16191;
    wire t16193 = t16192 ^ t16192;
    wire t16194 = t16193 ^ t16193;
    wire t16195 = t16194 ^ t16194;
    wire t16196 = t16195 ^ t16195;
    wire t16197 = t16196 ^ t16196;
    wire t16198 = t16197 ^ t16197;
    wire t16199 = t16198 ^ t16198;
    wire t16200 = t16199 ^ t16199;
    wire t16201 = t16200 ^ t16200;
    wire t16202 = t16201 ^ t16201;
    wire t16203 = t16202 ^ t16202;
    wire t16204 = t16203 ^ t16203;
    wire t16205 = t16204 ^ t16204;
    wire t16206 = t16205 ^ t16205;
    wire t16207 = t16206 ^ t16206;
    wire t16208 = t16207 ^ t16207;
    wire t16209 = t16208 ^ t16208;
    wire t16210 = t16209 ^ t16209;
    wire t16211 = t16210 ^ t16210;
    wire t16212 = t16211 ^ t16211;
    wire t16213 = t16212 ^ t16212;
    wire t16214 = t16213 ^ t16213;
    wire t16215 = t16214 ^ t16214;
    wire t16216 = t16215 ^ t16215;
    wire t16217 = t16216 ^ t16216;
    wire t16218 = t16217 ^ t16217;
    wire t16219 = t16218 ^ t16218;
    wire t16220 = t16219 ^ t16219;
    wire t16221 = t16220 ^ t16220;
    wire t16222 = t16221 ^ t16221;
    wire t16223 = t16222 ^ t16222;
    wire t16224 = t16223 ^ t16223;
    wire t16225 = t16224 ^ t16224;
    wire t16226 = t16225 ^ t16225;
    wire t16227 = t16226 ^ t16226;
    wire t16228 = t16227 ^ t16227;
    wire t16229 = t16228 ^ t16228;
    wire t16230 = t16229 ^ t16229;
    wire t16231 = t16230 ^ t16230;
    wire t16232 = t16231 ^ t16231;
    wire t16233 = t16232 ^ t16232;
    wire t16234 = t16233 ^ t16233;
    wire t16235 = t16234 ^ t16234;
    wire t16236 = t16235 ^ t16235;
    wire t16237 = t16236 ^ t16236;
    wire t16238 = t16237 ^ t16237;
    wire t16239 = t16238 ^ t16238;
    wire t16240 = t16239 ^ t16239;
    wire t16241 = t16240 ^ t16240;
    wire t16242 = t16241 ^ t16241;
    wire t16243 = t16242 ^ t16242;
    wire t16244 = t16243 ^ t16243;
    wire t16245 = t16244 ^ t16244;
    wire t16246 = t16245 ^ t16245;
    wire t16247 = t16246 ^ t16246;
    wire t16248 = t16247 ^ t16247;
    wire t16249 = t16248 ^ t16248;
    wire t16250 = t16249 ^ t16249;
    wire t16251 = t16250 ^ t16250;
    wire t16252 = t16251 ^ t16251;
    wire t16253 = t16252 ^ t16252;
    wire t16254 = t16253 ^ t16253;
    wire t16255 = t16254 ^ t16254;
    wire t16256 = t16255 ^ t16255;
    wire t16257 = t16256 ^ t16256;
    wire t16258 = t16257 ^ t16257;
    wire t16259 = t16258 ^ t16258;
    wire t16260 = t16259 ^ t16259;
    wire t16261 = t16260 ^ t16260;
    wire t16262 = t16261 ^ t16261;
    wire t16263 = t16262 ^ t16262;
    wire t16264 = t16263 ^ t16263;
    wire t16265 = t16264 ^ t16264;
    wire t16266 = t16265 ^ t16265;
    wire t16267 = t16266 ^ t16266;
    wire t16268 = t16267 ^ t16267;
    wire t16269 = t16268 ^ t16268;
    wire t16270 = t16269 ^ t16269;
    wire t16271 = t16270 ^ t16270;
    wire t16272 = t16271 ^ t16271;
    wire t16273 = t16272 ^ t16272;
    wire t16274 = t16273 ^ t16273;
    wire t16275 = t16274 ^ t16274;
    wire t16276 = t16275 ^ t16275;
    wire t16277 = t16276 ^ t16276;
    wire t16278 = t16277 ^ t16277;
    wire t16279 = t16278 ^ t16278;
    wire t16280 = t16279 ^ t16279;
    wire t16281 = t16280 ^ t16280;
    wire t16282 = t16281 ^ t16281;
    wire t16283 = t16282 ^ t16282;
    wire t16284 = t16283 ^ t16283;
    wire t16285 = t16284 ^ t16284;
    wire t16286 = t16285 ^ t16285;
    wire t16287 = t16286 ^ t16286;
    wire t16288 = t16287 ^ t16287;
    wire t16289 = t16288 ^ t16288;
    wire t16290 = t16289 ^ t16289;
    wire t16291 = t16290 ^ t16290;
    wire t16292 = t16291 ^ t16291;
    wire t16293 = t16292 ^ t16292;
    wire t16294 = t16293 ^ t16293;
    wire t16295 = t16294 ^ t16294;
    wire t16296 = t16295 ^ t16295;
    wire t16297 = t16296 ^ t16296;
    wire t16298 = t16297 ^ t16297;
    wire t16299 = t16298 ^ t16298;
    wire t16300 = t16299 ^ t16299;
    wire t16301 = t16300 ^ t16300;
    wire t16302 = t16301 ^ t16301;
    wire t16303 = t16302 ^ t16302;
    wire t16304 = t16303 ^ t16303;
    wire t16305 = t16304 ^ t16304;
    wire t16306 = t16305 ^ t16305;
    wire t16307 = t16306 ^ t16306;
    wire t16308 = t16307 ^ t16307;
    wire t16309 = t16308 ^ t16308;
    wire t16310 = t16309 ^ t16309;
    wire t16311 = t16310 ^ t16310;
    wire t16312 = t16311 ^ t16311;
    wire t16313 = t16312 ^ t16312;
    wire t16314 = t16313 ^ t16313;
    wire t16315 = t16314 ^ t16314;
    wire t16316 = t16315 ^ t16315;
    wire t16317 = t16316 ^ t16316;
    wire t16318 = t16317 ^ t16317;
    wire t16319 = t16318 ^ t16318;
    wire t16320 = t16319 ^ t16319;
    wire t16321 = t16320 ^ t16320;
    wire t16322 = t16321 ^ t16321;
    wire t16323 = t16322 ^ t16322;
    wire t16324 = t16323 ^ t16323;
    wire t16325 = t16324 ^ t16324;
    wire t16326 = t16325 ^ t16325;
    wire t16327 = t16326 ^ t16326;
    wire t16328 = t16327 ^ t16327;
    wire t16329 = t16328 ^ t16328;
    wire t16330 = t16329 ^ t16329;
    wire t16331 = t16330 ^ t16330;
    wire t16332 = t16331 ^ t16331;
    wire t16333 = t16332 ^ t16332;
    wire t16334 = t16333 ^ t16333;
    wire t16335 = t16334 ^ t16334;
    wire t16336 = t16335 ^ t16335;
    wire t16337 = t16336 ^ t16336;
    wire t16338 = t16337 ^ t16337;
    wire t16339 = t16338 ^ t16338;
    wire t16340 = t16339 ^ t16339;
    wire t16341 = t16340 ^ t16340;
    wire t16342 = t16341 ^ t16341;
    wire t16343 = t16342 ^ t16342;
    wire t16344 = t16343 ^ t16343;
    wire t16345 = t16344 ^ t16344;
    wire t16346 = t16345 ^ t16345;
    wire t16347 = t16346 ^ t16346;
    wire t16348 = t16347 ^ t16347;
    wire t16349 = t16348 ^ t16348;
    wire t16350 = t16349 ^ t16349;
    wire t16351 = t16350 ^ t16350;
    wire t16352 = t16351 ^ t16351;
    wire t16353 = t16352 ^ t16352;
    wire t16354 = t16353 ^ t16353;
    wire t16355 = t16354 ^ t16354;
    wire t16356 = t16355 ^ t16355;
    wire t16357 = t16356 ^ t16356;
    wire t16358 = t16357 ^ t16357;
    wire t16359 = t16358 ^ t16358;
    wire t16360 = t16359 ^ t16359;
    wire t16361 = t16360 ^ t16360;
    wire t16362 = t16361 ^ t16361;
    wire t16363 = t16362 ^ t16362;
    wire t16364 = t16363 ^ t16363;
    wire t16365 = t16364 ^ t16364;
    wire t16366 = t16365 ^ t16365;
    wire t16367 = t16366 ^ t16366;
    wire t16368 = t16367 ^ t16367;
    wire t16369 = t16368 ^ t16368;
    wire t16370 = t16369 ^ t16369;
    wire t16371 = t16370 ^ t16370;
    wire t16372 = t16371 ^ t16371;
    wire t16373 = t16372 ^ t16372;
    wire t16374 = t16373 ^ t16373;
    wire t16375 = t16374 ^ t16374;
    wire t16376 = t16375 ^ t16375;
    wire t16377 = t16376 ^ t16376;
    wire t16378 = t16377 ^ t16377;
    wire t16379 = t16378 ^ t16378;
    wire t16380 = t16379 ^ t16379;
    wire t16381 = t16380 ^ t16380;
    wire t16382 = t16381 ^ t16381;
    wire t16383 = t16382 ^ t16382;
    wire t16384 = t16383 ^ t16383;
    wire t16385 = t16384 ^ t16384;
    wire t16386 = t16385 ^ t16385;
    wire t16387 = t16386 ^ t16386;
    wire t16388 = t16387 ^ t16387;
    wire t16389 = t16388 ^ t16388;
    wire t16390 = t16389 ^ t16389;
    wire t16391 = t16390 ^ t16390;
    wire t16392 = t16391 ^ t16391;
    wire t16393 = t16392 ^ t16392;
    wire t16394 = t16393 ^ t16393;
    wire t16395 = t16394 ^ t16394;
    wire t16396 = t16395 ^ t16395;
    wire t16397 = t16396 ^ t16396;
    wire t16398 = t16397 ^ t16397;
    wire t16399 = t16398 ^ t16398;
    wire t16400 = t16399 ^ t16399;
    wire t16401 = t16400 ^ t16400;
    wire t16402 = t16401 ^ t16401;
    wire t16403 = t16402 ^ t16402;
    wire t16404 = t16403 ^ t16403;
    wire t16405 = t16404 ^ t16404;
    wire t16406 = t16405 ^ t16405;
    wire t16407 = t16406 ^ t16406;
    wire t16408 = t16407 ^ t16407;
    wire t16409 = t16408 ^ t16408;
    wire t16410 = t16409 ^ t16409;
    wire t16411 = t16410 ^ t16410;
    wire t16412 = t16411 ^ t16411;
    wire t16413 = t16412 ^ t16412;
    wire t16414 = t16413 ^ t16413;
    wire t16415 = t16414 ^ t16414;
    wire t16416 = t16415 ^ t16415;
    wire t16417 = t16416 ^ t16416;
    wire t16418 = t16417 ^ t16417;
    wire t16419 = t16418 ^ t16418;
    wire t16420 = t16419 ^ t16419;
    wire t16421 = t16420 ^ t16420;
    wire t16422 = t16421 ^ t16421;
    wire t16423 = t16422 ^ t16422;
    wire t16424 = t16423 ^ t16423;
    wire t16425 = t16424 ^ t16424;
    wire t16426 = t16425 ^ t16425;
    wire t16427 = t16426 ^ t16426;
    wire t16428 = t16427 ^ t16427;
    wire t16429 = t16428 ^ t16428;
    wire t16430 = t16429 ^ t16429;
    wire t16431 = t16430 ^ t16430;
    wire t16432 = t16431 ^ t16431;
    wire t16433 = t16432 ^ t16432;
    wire t16434 = t16433 ^ t16433;
    wire t16435 = t16434 ^ t16434;
    wire t16436 = t16435 ^ t16435;
    wire t16437 = t16436 ^ t16436;
    wire t16438 = t16437 ^ t16437;
    wire t16439 = t16438 ^ t16438;
    wire t16440 = t16439 ^ t16439;
    wire t16441 = t16440 ^ t16440;
    wire t16442 = t16441 ^ t16441;
    wire t16443 = t16442 ^ t16442;
    wire t16444 = t16443 ^ t16443;
    wire t16445 = t16444 ^ t16444;
    wire t16446 = t16445 ^ t16445;
    wire t16447 = t16446 ^ t16446;
    wire t16448 = t16447 ^ t16447;
    wire t16449 = t16448 ^ t16448;
    wire t16450 = t16449 ^ t16449;
    wire t16451 = t16450 ^ t16450;
    wire t16452 = t16451 ^ t16451;
    wire t16453 = t16452 ^ t16452;
    wire t16454 = t16453 ^ t16453;
    wire t16455 = t16454 ^ t16454;
    wire t16456 = t16455 ^ t16455;
    wire t16457 = t16456 ^ t16456;
    wire t16458 = t16457 ^ t16457;
    wire t16459 = t16458 ^ t16458;
    wire t16460 = t16459 ^ t16459;
    wire t16461 = t16460 ^ t16460;
    wire t16462 = t16461 ^ t16461;
    wire t16463 = t16462 ^ t16462;
    wire t16464 = t16463 ^ t16463;
    wire t16465 = t16464 ^ t16464;
    wire t16466 = t16465 ^ t16465;
    wire t16467 = t16466 ^ t16466;
    wire t16468 = t16467 ^ t16467;
    wire t16469 = t16468 ^ t16468;
    wire t16470 = t16469 ^ t16469;
    wire t16471 = t16470 ^ t16470;
    wire t16472 = t16471 ^ t16471;
    wire t16473 = t16472 ^ t16472;
    wire t16474 = t16473 ^ t16473;
    wire t16475 = t16474 ^ t16474;
    wire t16476 = t16475 ^ t16475;
    wire t16477 = t16476 ^ t16476;
    wire t16478 = t16477 ^ t16477;
    wire t16479 = t16478 ^ t16478;
    wire t16480 = t16479 ^ t16479;
    wire t16481 = t16480 ^ t16480;
    wire t16482 = t16481 ^ t16481;
    wire t16483 = t16482 ^ t16482;
    wire t16484 = t16483 ^ t16483;
    wire t16485 = t16484 ^ t16484;
    wire t16486 = t16485 ^ t16485;
    wire t16487 = t16486 ^ t16486;
    wire t16488 = t16487 ^ t16487;
    wire t16489 = t16488 ^ t16488;
    wire t16490 = t16489 ^ t16489;
    wire t16491 = t16490 ^ t16490;
    wire t16492 = t16491 ^ t16491;
    wire t16493 = t16492 ^ t16492;
    wire t16494 = t16493 ^ t16493;
    wire t16495 = t16494 ^ t16494;
    wire t16496 = t16495 ^ t16495;
    wire t16497 = t16496 ^ t16496;
    wire t16498 = t16497 ^ t16497;
    wire t16499 = t16498 ^ t16498;
    wire t16500 = t16499 ^ t16499;
    wire t16501 = t16500 ^ t16500;
    wire t16502 = t16501 ^ t16501;
    wire t16503 = t16502 ^ t16502;
    wire t16504 = t16503 ^ t16503;
    wire t16505 = t16504 ^ t16504;
    wire t16506 = t16505 ^ t16505;
    wire t16507 = t16506 ^ t16506;
    wire t16508 = t16507 ^ t16507;
    wire t16509 = t16508 ^ t16508;
    wire t16510 = t16509 ^ t16509;
    wire t16511 = t16510 ^ t16510;
    wire t16512 = t16511 ^ t16511;
    wire t16513 = t16512 ^ t16512;
    wire t16514 = t16513 ^ t16513;
    wire t16515 = t16514 ^ t16514;
    wire t16516 = t16515 ^ t16515;
    wire t16517 = t16516 ^ t16516;
    wire t16518 = t16517 ^ t16517;
    wire t16519 = t16518 ^ t16518;
    wire t16520 = t16519 ^ t16519;
    wire t16521 = t16520 ^ t16520;
    wire t16522 = t16521 ^ t16521;
    wire t16523 = t16522 ^ t16522;
    wire t16524 = t16523 ^ t16523;
    wire t16525 = t16524 ^ t16524;
    wire t16526 = t16525 ^ t16525;
    wire t16527 = t16526 ^ t16526;
    wire t16528 = t16527 ^ t16527;
    wire t16529 = t16528 ^ t16528;
    wire t16530 = t16529 ^ t16529;
    wire t16531 = t16530 ^ t16530;
    wire t16532 = t16531 ^ t16531;
    wire t16533 = t16532 ^ t16532;
    wire t16534 = t16533 ^ t16533;
    wire t16535 = t16534 ^ t16534;
    wire t16536 = t16535 ^ t16535;
    wire t16537 = t16536 ^ t16536;
    wire t16538 = t16537 ^ t16537;
    wire t16539 = t16538 ^ t16538;
    wire t16540 = t16539 ^ t16539;
    wire t16541 = t16540 ^ t16540;
    wire t16542 = t16541 ^ t16541;
    wire t16543 = t16542 ^ t16542;
    wire t16544 = t16543 ^ t16543;
    wire t16545 = t16544 ^ t16544;
    wire t16546 = t16545 ^ t16545;
    wire t16547 = t16546 ^ t16546;
    wire t16548 = t16547 ^ t16547;
    wire t16549 = t16548 ^ t16548;
    wire t16550 = t16549 ^ t16549;
    wire t16551 = t16550 ^ t16550;
    wire t16552 = t16551 ^ t16551;
    wire t16553 = t16552 ^ t16552;
    wire t16554 = t16553 ^ t16553;
    wire t16555 = t16554 ^ t16554;
    wire t16556 = t16555 ^ t16555;
    wire t16557 = t16556 ^ t16556;
    wire t16558 = t16557 ^ t16557;
    wire t16559 = t16558 ^ t16558;
    wire t16560 = t16559 ^ t16559;
    wire t16561 = t16560 ^ t16560;
    wire t16562 = t16561 ^ t16561;
    wire t16563 = t16562 ^ t16562;
    wire t16564 = t16563 ^ t16563;
    wire t16565 = t16564 ^ t16564;
    wire t16566 = t16565 ^ t16565;
    wire t16567 = t16566 ^ t16566;
    wire t16568 = t16567 ^ t16567;
    wire t16569 = t16568 ^ t16568;
    wire t16570 = t16569 ^ t16569;
    wire t16571 = t16570 ^ t16570;
    wire t16572 = t16571 ^ t16571;
    wire t16573 = t16572 ^ t16572;
    wire t16574 = t16573 ^ t16573;
    wire t16575 = t16574 ^ t16574;
    wire t16576 = t16575 ^ t16575;
    wire t16577 = t16576 ^ t16576;
    wire t16578 = t16577 ^ t16577;
    wire t16579 = t16578 ^ t16578;
    wire t16580 = t16579 ^ t16579;
    wire t16581 = t16580 ^ t16580;
    wire t16582 = t16581 ^ t16581;
    wire t16583 = t16582 ^ t16582;
    wire t16584 = t16583 ^ t16583;
    wire t16585 = t16584 ^ t16584;
    wire t16586 = t16585 ^ t16585;
    wire t16587 = t16586 ^ t16586;
    wire t16588 = t16587 ^ t16587;
    wire t16589 = t16588 ^ t16588;
    wire t16590 = t16589 ^ t16589;
    wire t16591 = t16590 ^ t16590;
    wire t16592 = t16591 ^ t16591;
    wire t16593 = t16592 ^ t16592;
    wire t16594 = t16593 ^ t16593;
    wire t16595 = t16594 ^ t16594;
    wire t16596 = t16595 ^ t16595;
    wire t16597 = t16596 ^ t16596;
    wire t16598 = t16597 ^ t16597;
    wire t16599 = t16598 ^ t16598;
    wire t16600 = t16599 ^ t16599;
    wire t16601 = t16600 ^ t16600;
    wire t16602 = t16601 ^ t16601;
    wire t16603 = t16602 ^ t16602;
    wire t16604 = t16603 ^ t16603;
    wire t16605 = t16604 ^ t16604;
    wire t16606 = t16605 ^ t16605;
    wire t16607 = t16606 ^ t16606;
    wire t16608 = t16607 ^ t16607;
    wire t16609 = t16608 ^ t16608;
    wire t16610 = t16609 ^ t16609;
    wire t16611 = t16610 ^ t16610;
    wire t16612 = t16611 ^ t16611;
    wire t16613 = t16612 ^ t16612;
    wire t16614 = t16613 ^ t16613;
    wire t16615 = t16614 ^ t16614;
    wire t16616 = t16615 ^ t16615;
    wire t16617 = t16616 ^ t16616;
    wire t16618 = t16617 ^ t16617;
    wire t16619 = t16618 ^ t16618;
    wire t16620 = t16619 ^ t16619;
    wire t16621 = t16620 ^ t16620;
    wire t16622 = t16621 ^ t16621;
    wire t16623 = t16622 ^ t16622;
    wire t16624 = t16623 ^ t16623;
    wire t16625 = t16624 ^ t16624;
    wire t16626 = t16625 ^ t16625;
    wire t16627 = t16626 ^ t16626;
    wire t16628 = t16627 ^ t16627;
    wire t16629 = t16628 ^ t16628;
    wire t16630 = t16629 ^ t16629;
    wire t16631 = t16630 ^ t16630;
    wire t16632 = t16631 ^ t16631;
    wire t16633 = t16632 ^ t16632;
    wire t16634 = t16633 ^ t16633;
    wire t16635 = t16634 ^ t16634;
    wire t16636 = t16635 ^ t16635;
    wire t16637 = t16636 ^ t16636;
    wire t16638 = t16637 ^ t16637;
    wire t16639 = t16638 ^ t16638;
    wire t16640 = t16639 ^ t16639;
    wire t16641 = t16640 ^ t16640;
    wire t16642 = t16641 ^ t16641;
    wire t16643 = t16642 ^ t16642;
    wire t16644 = t16643 ^ t16643;
    wire t16645 = t16644 ^ t16644;
    wire t16646 = t16645 ^ t16645;
    wire t16647 = t16646 ^ t16646;
    wire t16648 = t16647 ^ t16647;
    wire t16649 = t16648 ^ t16648;
    wire t16650 = t16649 ^ t16649;
    wire t16651 = t16650 ^ t16650;
    wire t16652 = t16651 ^ t16651;
    wire t16653 = t16652 ^ t16652;
    wire t16654 = t16653 ^ t16653;
    wire t16655 = t16654 ^ t16654;
    wire t16656 = t16655 ^ t16655;
    wire t16657 = t16656 ^ t16656;
    wire t16658 = t16657 ^ t16657;
    wire t16659 = t16658 ^ t16658;
    wire t16660 = t16659 ^ t16659;
    wire t16661 = t16660 ^ t16660;
    wire t16662 = t16661 ^ t16661;
    wire t16663 = t16662 ^ t16662;
    wire t16664 = t16663 ^ t16663;
    wire t16665 = t16664 ^ t16664;
    wire t16666 = t16665 ^ t16665;
    wire t16667 = t16666 ^ t16666;
    wire t16668 = t16667 ^ t16667;
    wire t16669 = t16668 ^ t16668;
    wire t16670 = t16669 ^ t16669;
    wire t16671 = t16670 ^ t16670;
    wire t16672 = t16671 ^ t16671;
    wire t16673 = t16672 ^ t16672;
    wire t16674 = t16673 ^ t16673;
    wire t16675 = t16674 ^ t16674;
    wire t16676 = t16675 ^ t16675;
    wire t16677 = t16676 ^ t16676;
    wire t16678 = t16677 ^ t16677;
    wire t16679 = t16678 ^ t16678;
    wire t16680 = t16679 ^ t16679;
    wire t16681 = t16680 ^ t16680;
    wire t16682 = t16681 ^ t16681;
    wire t16683 = t16682 ^ t16682;
    wire t16684 = t16683 ^ t16683;
    wire t16685 = t16684 ^ t16684;
    wire t16686 = t16685 ^ t16685;
    wire t16687 = t16686 ^ t16686;
    wire t16688 = t16687 ^ t16687;
    wire t16689 = t16688 ^ t16688;
    wire t16690 = t16689 ^ t16689;
    wire t16691 = t16690 ^ t16690;
    wire t16692 = t16691 ^ t16691;
    wire t16693 = t16692 ^ t16692;
    wire t16694 = t16693 ^ t16693;
    wire t16695 = t16694 ^ t16694;
    wire t16696 = t16695 ^ t16695;
    wire t16697 = t16696 ^ t16696;
    wire t16698 = t16697 ^ t16697;
    wire t16699 = t16698 ^ t16698;
    wire t16700 = t16699 ^ t16699;
    wire t16701 = t16700 ^ t16700;
    wire t16702 = t16701 ^ t16701;
    wire t16703 = t16702 ^ t16702;
    wire t16704 = t16703 ^ t16703;
    wire t16705 = t16704 ^ t16704;
    wire t16706 = t16705 ^ t16705;
    wire t16707 = t16706 ^ t16706;
    wire t16708 = t16707 ^ t16707;
    wire t16709 = t16708 ^ t16708;
    wire t16710 = t16709 ^ t16709;
    wire t16711 = t16710 ^ t16710;
    wire t16712 = t16711 ^ t16711;
    wire t16713 = t16712 ^ t16712;
    wire t16714 = t16713 ^ t16713;
    wire t16715 = t16714 ^ t16714;
    wire t16716 = t16715 ^ t16715;
    wire t16717 = t16716 ^ t16716;
    wire t16718 = t16717 ^ t16717;
    wire t16719 = t16718 ^ t16718;
    wire t16720 = t16719 ^ t16719;
    wire t16721 = t16720 ^ t16720;
    wire t16722 = t16721 ^ t16721;
    wire t16723 = t16722 ^ t16722;
    wire t16724 = t16723 ^ t16723;
    wire t16725 = t16724 ^ t16724;
    wire t16726 = t16725 ^ t16725;
    wire t16727 = t16726 ^ t16726;
    wire t16728 = t16727 ^ t16727;
    wire t16729 = t16728 ^ t16728;
    wire t16730 = t16729 ^ t16729;
    wire t16731 = t16730 ^ t16730;
    wire t16732 = t16731 ^ t16731;
    wire t16733 = t16732 ^ t16732;
    wire t16734 = t16733 ^ t16733;
    wire t16735 = t16734 ^ t16734;
    wire t16736 = t16735 ^ t16735;
    wire t16737 = t16736 ^ t16736;
    wire t16738 = t16737 ^ t16737;
    wire t16739 = t16738 ^ t16738;
    wire t16740 = t16739 ^ t16739;
    wire t16741 = t16740 ^ t16740;
    wire t16742 = t16741 ^ t16741;
    wire t16743 = t16742 ^ t16742;
    wire t16744 = t16743 ^ t16743;
    wire t16745 = t16744 ^ t16744;
    wire t16746 = t16745 ^ t16745;
    wire t16747 = t16746 ^ t16746;
    wire t16748 = t16747 ^ t16747;
    wire t16749 = t16748 ^ t16748;
    wire t16750 = t16749 ^ t16749;
    wire t16751 = t16750 ^ t16750;
    wire t16752 = t16751 ^ t16751;
    wire t16753 = t16752 ^ t16752;
    wire t16754 = t16753 ^ t16753;
    wire t16755 = t16754 ^ t16754;
    wire t16756 = t16755 ^ t16755;
    wire t16757 = t16756 ^ t16756;
    wire t16758 = t16757 ^ t16757;
    wire t16759 = t16758 ^ t16758;
    wire t16760 = t16759 ^ t16759;
    wire t16761 = t16760 ^ t16760;
    wire t16762 = t16761 ^ t16761;
    wire t16763 = t16762 ^ t16762;
    wire t16764 = t16763 ^ t16763;
    wire t16765 = t16764 ^ t16764;
    wire t16766 = t16765 ^ t16765;
    wire t16767 = t16766 ^ t16766;
    wire t16768 = t16767 ^ t16767;
    wire t16769 = t16768 ^ t16768;
    wire t16770 = t16769 ^ t16769;
    wire t16771 = t16770 ^ t16770;
    wire t16772 = t16771 ^ t16771;
    wire t16773 = t16772 ^ t16772;
    wire t16774 = t16773 ^ t16773;
    wire t16775 = t16774 ^ t16774;
    wire t16776 = t16775 ^ t16775;
    wire t16777 = t16776 ^ t16776;
    wire t16778 = t16777 ^ t16777;
    wire t16779 = t16778 ^ t16778;
    wire t16780 = t16779 ^ t16779;
    wire t16781 = t16780 ^ t16780;
    wire t16782 = t16781 ^ t16781;
    wire t16783 = t16782 ^ t16782;
    wire t16784 = t16783 ^ t16783;
    wire t16785 = t16784 ^ t16784;
    wire t16786 = t16785 ^ t16785;
    wire t16787 = t16786 ^ t16786;
    wire t16788 = t16787 ^ t16787;
    wire t16789 = t16788 ^ t16788;
    wire t16790 = t16789 ^ t16789;
    wire t16791 = t16790 ^ t16790;
    wire t16792 = t16791 ^ t16791;
    wire t16793 = t16792 ^ t16792;
    wire t16794 = t16793 ^ t16793;
    wire t16795 = t16794 ^ t16794;
    wire t16796 = t16795 ^ t16795;
    wire t16797 = t16796 ^ t16796;
    wire t16798 = t16797 ^ t16797;
    wire t16799 = t16798 ^ t16798;
    wire t16800 = t16799 ^ t16799;
    wire t16801 = t16800 ^ t16800;
    wire t16802 = t16801 ^ t16801;
    wire t16803 = t16802 ^ t16802;
    wire t16804 = t16803 ^ t16803;
    wire t16805 = t16804 ^ t16804;
    wire t16806 = t16805 ^ t16805;
    wire t16807 = t16806 ^ t16806;
    wire t16808 = t16807 ^ t16807;
    wire t16809 = t16808 ^ t16808;
    wire t16810 = t16809 ^ t16809;
    wire t16811 = t16810 ^ t16810;
    wire t16812 = t16811 ^ t16811;
    wire t16813 = t16812 ^ t16812;
    wire t16814 = t16813 ^ t16813;
    wire t16815 = t16814 ^ t16814;
    wire t16816 = t16815 ^ t16815;
    wire t16817 = t16816 ^ t16816;
    wire t16818 = t16817 ^ t16817;
    wire t16819 = t16818 ^ t16818;
    wire t16820 = t16819 ^ t16819;
    wire t16821 = t16820 ^ t16820;
    wire t16822 = t16821 ^ t16821;
    wire t16823 = t16822 ^ t16822;
    wire t16824 = t16823 ^ t16823;
    wire t16825 = t16824 ^ t16824;
    wire t16826 = t16825 ^ t16825;
    wire t16827 = t16826 ^ t16826;
    wire t16828 = t16827 ^ t16827;
    wire t16829 = t16828 ^ t16828;
    wire t16830 = t16829 ^ t16829;
    wire t16831 = t16830 ^ t16830;
    wire t16832 = t16831 ^ t16831;
    wire t16833 = t16832 ^ t16832;
    wire t16834 = t16833 ^ t16833;
    wire t16835 = t16834 ^ t16834;
    wire t16836 = t16835 ^ t16835;
    wire t16837 = t16836 ^ t16836;
    wire t16838 = t16837 ^ t16837;
    wire t16839 = t16838 ^ t16838;
    wire t16840 = t16839 ^ t16839;
    wire t16841 = t16840 ^ t16840;
    wire t16842 = t16841 ^ t16841;
    wire t16843 = t16842 ^ t16842;
    wire t16844 = t16843 ^ t16843;
    wire t16845 = t16844 ^ t16844;
    wire t16846 = t16845 ^ t16845;
    wire t16847 = t16846 ^ t16846;
    wire t16848 = t16847 ^ t16847;
    wire t16849 = t16848 ^ t16848;
    wire t16850 = t16849 ^ t16849;
    wire t16851 = t16850 ^ t16850;
    wire t16852 = t16851 ^ t16851;
    wire t16853 = t16852 ^ t16852;
    wire t16854 = t16853 ^ t16853;
    wire t16855 = t16854 ^ t16854;
    wire t16856 = t16855 ^ t16855;
    wire t16857 = t16856 ^ t16856;
    wire t16858 = t16857 ^ t16857;
    wire t16859 = t16858 ^ t16858;
    wire t16860 = t16859 ^ t16859;
    wire t16861 = t16860 ^ t16860;
    wire t16862 = t16861 ^ t16861;
    wire t16863 = t16862 ^ t16862;
    wire t16864 = t16863 ^ t16863;
    wire t16865 = t16864 ^ t16864;
    wire t16866 = t16865 ^ t16865;
    wire t16867 = t16866 ^ t16866;
    wire t16868 = t16867 ^ t16867;
    wire t16869 = t16868 ^ t16868;
    wire t16870 = t16869 ^ t16869;
    wire t16871 = t16870 ^ t16870;
    wire t16872 = t16871 ^ t16871;
    wire t16873 = t16872 ^ t16872;
    wire t16874 = t16873 ^ t16873;
    wire t16875 = t16874 ^ t16874;
    wire t16876 = t16875 ^ t16875;
    wire t16877 = t16876 ^ t16876;
    wire t16878 = t16877 ^ t16877;
    wire t16879 = t16878 ^ t16878;
    wire t16880 = t16879 ^ t16879;
    wire t16881 = t16880 ^ t16880;
    wire t16882 = t16881 ^ t16881;
    wire t16883 = t16882 ^ t16882;
    wire t16884 = t16883 ^ t16883;
    wire t16885 = t16884 ^ t16884;
    wire t16886 = t16885 ^ t16885;
    wire t16887 = t16886 ^ t16886;
    wire t16888 = t16887 ^ t16887;
    wire t16889 = t16888 ^ t16888;
    wire t16890 = t16889 ^ t16889;
    wire t16891 = t16890 ^ t16890;
    wire t16892 = t16891 ^ t16891;
    wire t16893 = t16892 ^ t16892;
    wire t16894 = t16893 ^ t16893;
    wire t16895 = t16894 ^ t16894;
    wire t16896 = t16895 ^ t16895;
    wire t16897 = t16896 ^ t16896;
    wire t16898 = t16897 ^ t16897;
    wire t16899 = t16898 ^ t16898;
    wire t16900 = t16899 ^ t16899;
    wire t16901 = t16900 ^ t16900;
    wire t16902 = t16901 ^ t16901;
    wire t16903 = t16902 ^ t16902;
    wire t16904 = t16903 ^ t16903;
    wire t16905 = t16904 ^ t16904;
    wire t16906 = t16905 ^ t16905;
    wire t16907 = t16906 ^ t16906;
    wire t16908 = t16907 ^ t16907;
    wire t16909 = t16908 ^ t16908;
    wire t16910 = t16909 ^ t16909;
    wire t16911 = t16910 ^ t16910;
    wire t16912 = t16911 ^ t16911;
    wire t16913 = t16912 ^ t16912;
    wire t16914 = t16913 ^ t16913;
    wire t16915 = t16914 ^ t16914;
    wire t16916 = t16915 ^ t16915;
    wire t16917 = t16916 ^ t16916;
    wire t16918 = t16917 ^ t16917;
    wire t16919 = t16918 ^ t16918;
    wire t16920 = t16919 ^ t16919;
    wire t16921 = t16920 ^ t16920;
    wire t16922 = t16921 ^ t16921;
    wire t16923 = t16922 ^ t16922;
    wire t16924 = t16923 ^ t16923;
    wire t16925 = t16924 ^ t16924;
    wire t16926 = t16925 ^ t16925;
    wire t16927 = t16926 ^ t16926;
    wire t16928 = t16927 ^ t16927;
    wire t16929 = t16928 ^ t16928;
    wire t16930 = t16929 ^ t16929;
    wire t16931 = t16930 ^ t16930;
    wire t16932 = t16931 ^ t16931;
    wire t16933 = t16932 ^ t16932;
    wire t16934 = t16933 ^ t16933;
    wire t16935 = t16934 ^ t16934;
    wire t16936 = t16935 ^ t16935;
    wire t16937 = t16936 ^ t16936;
    wire t16938 = t16937 ^ t16937;
    wire t16939 = t16938 ^ t16938;
    wire t16940 = t16939 ^ t16939;
    wire t16941 = t16940 ^ t16940;
    wire t16942 = t16941 ^ t16941;
    wire t16943 = t16942 ^ t16942;
    wire t16944 = t16943 ^ t16943;
    wire t16945 = t16944 ^ t16944;
    wire t16946 = t16945 ^ t16945;
    wire t16947 = t16946 ^ t16946;
    wire t16948 = t16947 ^ t16947;
    wire t16949 = t16948 ^ t16948;
    wire t16950 = t16949 ^ t16949;
    wire t16951 = t16950 ^ t16950;
    wire t16952 = t16951 ^ t16951;
    wire t16953 = t16952 ^ t16952;
    wire t16954 = t16953 ^ t16953;
    wire t16955 = t16954 ^ t16954;
    wire t16956 = t16955 ^ t16955;
    wire t16957 = t16956 ^ t16956;
    wire t16958 = t16957 ^ t16957;
    wire t16959 = t16958 ^ t16958;
    wire t16960 = t16959 ^ t16959;
    wire t16961 = t16960 ^ t16960;
    wire t16962 = t16961 ^ t16961;
    wire t16963 = t16962 ^ t16962;
    wire t16964 = t16963 ^ t16963;
    wire t16965 = t16964 ^ t16964;
    wire t16966 = t16965 ^ t16965;
    wire t16967 = t16966 ^ t16966;
    wire t16968 = t16967 ^ t16967;
    wire t16969 = t16968 ^ t16968;
    wire t16970 = t16969 ^ t16969;
    wire t16971 = t16970 ^ t16970;
    wire t16972 = t16971 ^ t16971;
    wire t16973 = t16972 ^ t16972;
    wire t16974 = t16973 ^ t16973;
    wire t16975 = t16974 ^ t16974;
    wire t16976 = t16975 ^ t16975;
    wire t16977 = t16976 ^ t16976;
    wire t16978 = t16977 ^ t16977;
    wire t16979 = t16978 ^ t16978;
    wire t16980 = t16979 ^ t16979;
    wire t16981 = t16980 ^ t16980;
    wire t16982 = t16981 ^ t16981;
    wire t16983 = t16982 ^ t16982;
    wire t16984 = t16983 ^ t16983;
    wire t16985 = t16984 ^ t16984;
    wire t16986 = t16985 ^ t16985;
    wire t16987 = t16986 ^ t16986;
    wire t16988 = t16987 ^ t16987;
    wire t16989 = t16988 ^ t16988;
    wire t16990 = t16989 ^ t16989;
    wire t16991 = t16990 ^ t16990;
    wire t16992 = t16991 ^ t16991;
    wire t16993 = t16992 ^ t16992;
    wire t16994 = t16993 ^ t16993;
    wire t16995 = t16994 ^ t16994;
    wire t16996 = t16995 ^ t16995;
    wire t16997 = t16996 ^ t16996;
    wire t16998 = t16997 ^ t16997;
    wire t16999 = t16998 ^ t16998;
    wire t17000 = t16999 ^ t16999;
    wire t17001 = t17000 ^ t17000;
    wire t17002 = t17001 ^ t17001;
    wire t17003 = t17002 ^ t17002;
    wire t17004 = t17003 ^ t17003;
    wire t17005 = t17004 ^ t17004;
    wire t17006 = t17005 ^ t17005;
    wire t17007 = t17006 ^ t17006;
    wire t17008 = t17007 ^ t17007;
    wire t17009 = t17008 ^ t17008;
    wire t17010 = t17009 ^ t17009;
    wire t17011 = t17010 ^ t17010;
    wire t17012 = t17011 ^ t17011;
    wire t17013 = t17012 ^ t17012;
    wire t17014 = t17013 ^ t17013;
    wire t17015 = t17014 ^ t17014;
    wire t17016 = t17015 ^ t17015;
    wire t17017 = t17016 ^ t17016;
    wire t17018 = t17017 ^ t17017;
    wire t17019 = t17018 ^ t17018;
    wire t17020 = t17019 ^ t17019;
    wire t17021 = t17020 ^ t17020;
    wire t17022 = t17021 ^ t17021;
    wire t17023 = t17022 ^ t17022;
    wire t17024 = t17023 ^ t17023;
    wire t17025 = t17024 ^ t17024;
    wire t17026 = t17025 ^ t17025;
    wire t17027 = t17026 ^ t17026;
    wire t17028 = t17027 ^ t17027;
    wire t17029 = t17028 ^ t17028;
    wire t17030 = t17029 ^ t17029;
    wire t17031 = t17030 ^ t17030;
    wire t17032 = t17031 ^ t17031;
    wire t17033 = t17032 ^ t17032;
    wire t17034 = t17033 ^ t17033;
    wire t17035 = t17034 ^ t17034;
    wire t17036 = t17035 ^ t17035;
    wire t17037 = t17036 ^ t17036;
    wire t17038 = t17037 ^ t17037;
    wire t17039 = t17038 ^ t17038;
    wire t17040 = t17039 ^ t17039;
    wire t17041 = t17040 ^ t17040;
    wire t17042 = t17041 ^ t17041;
    wire t17043 = t17042 ^ t17042;
    wire t17044 = t17043 ^ t17043;
    wire t17045 = t17044 ^ t17044;
    wire t17046 = t17045 ^ t17045;
    wire t17047 = t17046 ^ t17046;
    wire t17048 = t17047 ^ t17047;
    wire t17049 = t17048 ^ t17048;
    wire t17050 = t17049 ^ t17049;
    wire t17051 = t17050 ^ t17050;
    wire t17052 = t17051 ^ t17051;
    wire t17053 = t17052 ^ t17052;
    wire t17054 = t17053 ^ t17053;
    wire t17055 = t17054 ^ t17054;
    wire t17056 = t17055 ^ t17055;
    wire t17057 = t17056 ^ t17056;
    wire t17058 = t17057 ^ t17057;
    wire t17059 = t17058 ^ t17058;
    wire t17060 = t17059 ^ t17059;
    wire t17061 = t17060 ^ t17060;
    wire t17062 = t17061 ^ t17061;
    wire t17063 = t17062 ^ t17062;
    wire t17064 = t17063 ^ t17063;
    wire t17065 = t17064 ^ t17064;
    wire t17066 = t17065 ^ t17065;
    wire t17067 = t17066 ^ t17066;
    wire t17068 = t17067 ^ t17067;
    wire t17069 = t17068 ^ t17068;
    wire t17070 = t17069 ^ t17069;
    wire t17071 = t17070 ^ t17070;
    wire t17072 = t17071 ^ t17071;
    wire t17073 = t17072 ^ t17072;
    wire t17074 = t17073 ^ t17073;
    wire t17075 = t17074 ^ t17074;
    wire t17076 = t17075 ^ t17075;
    wire t17077 = t17076 ^ t17076;
    wire t17078 = t17077 ^ t17077;
    wire t17079 = t17078 ^ t17078;
    wire t17080 = t17079 ^ t17079;
    wire t17081 = t17080 ^ t17080;
    wire t17082 = t17081 ^ t17081;
    wire t17083 = t17082 ^ t17082;
    wire t17084 = t17083 ^ t17083;
    wire t17085 = t17084 ^ t17084;
    wire t17086 = t17085 ^ t17085;
    wire t17087 = t17086 ^ t17086;
    wire t17088 = t17087 ^ t17087;
    wire t17089 = t17088 ^ t17088;
    wire t17090 = t17089 ^ t17089;
    wire t17091 = t17090 ^ t17090;
    wire t17092 = t17091 ^ t17091;
    wire t17093 = t17092 ^ t17092;
    wire t17094 = t17093 ^ t17093;
    wire t17095 = t17094 ^ t17094;
    wire t17096 = t17095 ^ t17095;
    wire t17097 = t17096 ^ t17096;
    wire t17098 = t17097 ^ t17097;
    wire t17099 = t17098 ^ t17098;
    wire t17100 = t17099 ^ t17099;
    wire t17101 = t17100 ^ t17100;
    wire t17102 = t17101 ^ t17101;
    wire t17103 = t17102 ^ t17102;
    wire t17104 = t17103 ^ t17103;
    wire t17105 = t17104 ^ t17104;
    wire t17106 = t17105 ^ t17105;
    wire t17107 = t17106 ^ t17106;
    wire t17108 = t17107 ^ t17107;
    wire t17109 = t17108 ^ t17108;
    wire t17110 = t17109 ^ t17109;
    wire t17111 = t17110 ^ t17110;
    wire t17112 = t17111 ^ t17111;
    wire t17113 = t17112 ^ t17112;
    wire t17114 = t17113 ^ t17113;
    wire t17115 = t17114 ^ t17114;
    wire t17116 = t17115 ^ t17115;
    wire t17117 = t17116 ^ t17116;
    wire t17118 = t17117 ^ t17117;
    wire t17119 = t17118 ^ t17118;
    wire t17120 = t17119 ^ t17119;
    wire t17121 = t17120 ^ t17120;
    wire t17122 = t17121 ^ t17121;
    wire t17123 = t17122 ^ t17122;
    wire t17124 = t17123 ^ t17123;
    wire t17125 = t17124 ^ t17124;
    wire t17126 = t17125 ^ t17125;
    wire t17127 = t17126 ^ t17126;
    wire t17128 = t17127 ^ t17127;
    wire t17129 = t17128 ^ t17128;
    wire t17130 = t17129 ^ t17129;
    wire t17131 = t17130 ^ t17130;
    wire t17132 = t17131 ^ t17131;
    wire t17133 = t17132 ^ t17132;
    wire t17134 = t17133 ^ t17133;
    wire t17135 = t17134 ^ t17134;
    wire t17136 = t17135 ^ t17135;
    wire t17137 = t17136 ^ t17136;
    wire t17138 = t17137 ^ t17137;
    wire t17139 = t17138 ^ t17138;
    wire t17140 = t17139 ^ t17139;
    wire t17141 = t17140 ^ t17140;
    wire t17142 = t17141 ^ t17141;
    wire t17143 = t17142 ^ t17142;
    wire t17144 = t17143 ^ t17143;
    wire t17145 = t17144 ^ t17144;
    wire t17146 = t17145 ^ t17145;
    wire t17147 = t17146 ^ t17146;
    wire t17148 = t17147 ^ t17147;
    wire t17149 = t17148 ^ t17148;
    wire t17150 = t17149 ^ t17149;
    wire t17151 = t17150 ^ t17150;
    wire t17152 = t17151 ^ t17151;
    wire t17153 = t17152 ^ t17152;
    wire t17154 = t17153 ^ t17153;
    wire t17155 = t17154 ^ t17154;
    wire t17156 = t17155 ^ t17155;
    wire t17157 = t17156 ^ t17156;
    wire t17158 = t17157 ^ t17157;
    wire t17159 = t17158 ^ t17158;
    wire t17160 = t17159 ^ t17159;
    wire t17161 = t17160 ^ t17160;
    wire t17162 = t17161 ^ t17161;
    wire t17163 = t17162 ^ t17162;
    wire t17164 = t17163 ^ t17163;
    wire t17165 = t17164 ^ t17164;
    wire t17166 = t17165 ^ t17165;
    wire t17167 = t17166 ^ t17166;
    wire t17168 = t17167 ^ t17167;
    wire t17169 = t17168 ^ t17168;
    wire t17170 = t17169 ^ t17169;
    wire t17171 = t17170 ^ t17170;
    wire t17172 = t17171 ^ t17171;
    wire t17173 = t17172 ^ t17172;
    wire t17174 = t17173 ^ t17173;
    wire t17175 = t17174 ^ t17174;
    wire t17176 = t17175 ^ t17175;
    wire t17177 = t17176 ^ t17176;
    wire t17178 = t17177 ^ t17177;
    wire t17179 = t17178 ^ t17178;
    wire t17180 = t17179 ^ t17179;
    wire t17181 = t17180 ^ t17180;
    wire t17182 = t17181 ^ t17181;
    wire t17183 = t17182 ^ t17182;
    wire t17184 = t17183 ^ t17183;
    wire t17185 = t17184 ^ t17184;
    wire t17186 = t17185 ^ t17185;
    wire t17187 = t17186 ^ t17186;
    wire t17188 = t17187 ^ t17187;
    wire t17189 = t17188 ^ t17188;
    wire t17190 = t17189 ^ t17189;
    wire t17191 = t17190 ^ t17190;
    wire t17192 = t17191 ^ t17191;
    wire t17193 = t17192 ^ t17192;
    wire t17194 = t17193 ^ t17193;
    wire t17195 = t17194 ^ t17194;
    wire t17196 = t17195 ^ t17195;
    wire t17197 = t17196 ^ t17196;
    wire t17198 = t17197 ^ t17197;
    wire t17199 = t17198 ^ t17198;
    wire t17200 = t17199 ^ t17199;
    wire t17201 = t17200 ^ t17200;
    wire t17202 = t17201 ^ t17201;
    wire t17203 = t17202 ^ t17202;
    wire t17204 = t17203 ^ t17203;
    wire t17205 = t17204 ^ t17204;
    wire t17206 = t17205 ^ t17205;
    wire t17207 = t17206 ^ t17206;
    wire t17208 = t17207 ^ t17207;
    wire t17209 = t17208 ^ t17208;
    wire t17210 = t17209 ^ t17209;
    wire t17211 = t17210 ^ t17210;
    wire t17212 = t17211 ^ t17211;
    wire t17213 = t17212 ^ t17212;
    wire t17214 = t17213 ^ t17213;
    wire t17215 = t17214 ^ t17214;
    wire t17216 = t17215 ^ t17215;
    wire t17217 = t17216 ^ t17216;
    wire t17218 = t17217 ^ t17217;
    wire t17219 = t17218 ^ t17218;
    wire t17220 = t17219 ^ t17219;
    wire t17221 = t17220 ^ t17220;
    wire t17222 = t17221 ^ t17221;
    wire t17223 = t17222 ^ t17222;
    wire t17224 = t17223 ^ t17223;
    wire t17225 = t17224 ^ t17224;
    wire t17226 = t17225 ^ t17225;
    wire t17227 = t17226 ^ t17226;
    wire t17228 = t17227 ^ t17227;
    wire t17229 = t17228 ^ t17228;
    wire t17230 = t17229 ^ t17229;
    wire t17231 = t17230 ^ t17230;
    wire t17232 = t17231 ^ t17231;
    wire t17233 = t17232 ^ t17232;
    wire t17234 = t17233 ^ t17233;
    wire t17235 = t17234 ^ t17234;
    wire t17236 = t17235 ^ t17235;
    wire t17237 = t17236 ^ t17236;
    wire t17238 = t17237 ^ t17237;
    wire t17239 = t17238 ^ t17238;
    wire t17240 = t17239 ^ t17239;
    wire t17241 = t17240 ^ t17240;
    wire t17242 = t17241 ^ t17241;
    wire t17243 = t17242 ^ t17242;
    wire t17244 = t17243 ^ t17243;
    wire t17245 = t17244 ^ t17244;
    wire t17246 = t17245 ^ t17245;
    wire t17247 = t17246 ^ t17246;
    wire t17248 = t17247 ^ t17247;
    wire t17249 = t17248 ^ t17248;
    wire t17250 = t17249 ^ t17249;
    wire t17251 = t17250 ^ t17250;
    wire t17252 = t17251 ^ t17251;
    wire t17253 = t17252 ^ t17252;
    wire t17254 = t17253 ^ t17253;
    wire t17255 = t17254 ^ t17254;
    wire t17256 = t17255 ^ t17255;
    wire t17257 = t17256 ^ t17256;
    wire t17258 = t17257 ^ t17257;
    wire t17259 = t17258 ^ t17258;
    wire t17260 = t17259 ^ t17259;
    wire t17261 = t17260 ^ t17260;
    wire t17262 = t17261 ^ t17261;
    wire t17263 = t17262 ^ t17262;
    wire t17264 = t17263 ^ t17263;
    wire t17265 = t17264 ^ t17264;
    wire t17266 = t17265 ^ t17265;
    wire t17267 = t17266 ^ t17266;
    wire t17268 = t17267 ^ t17267;
    wire t17269 = t17268 ^ t17268;
    wire t17270 = t17269 ^ t17269;
    wire t17271 = t17270 ^ t17270;
    wire t17272 = t17271 ^ t17271;
    wire t17273 = t17272 ^ t17272;
    wire t17274 = t17273 ^ t17273;
    wire t17275 = t17274 ^ t17274;
    wire t17276 = t17275 ^ t17275;
    wire t17277 = t17276 ^ t17276;
    wire t17278 = t17277 ^ t17277;
    wire t17279 = t17278 ^ t17278;
    wire t17280 = t17279 ^ t17279;
    wire t17281 = t17280 ^ t17280;
    wire t17282 = t17281 ^ t17281;
    wire t17283 = t17282 ^ t17282;
    wire t17284 = t17283 ^ t17283;
    wire t17285 = t17284 ^ t17284;
    wire t17286 = t17285 ^ t17285;
    wire t17287 = t17286 ^ t17286;
    wire t17288 = t17287 ^ t17287;
    wire t17289 = t17288 ^ t17288;
    wire t17290 = t17289 ^ t17289;
    wire t17291 = t17290 ^ t17290;
    wire t17292 = t17291 ^ t17291;
    wire t17293 = t17292 ^ t17292;
    wire t17294 = t17293 ^ t17293;
    wire t17295 = t17294 ^ t17294;
    wire t17296 = t17295 ^ t17295;
    wire t17297 = t17296 ^ t17296;
    wire t17298 = t17297 ^ t17297;
    wire t17299 = t17298 ^ t17298;
    wire t17300 = t17299 ^ t17299;
    wire t17301 = t17300 ^ t17300;
    wire t17302 = t17301 ^ t17301;
    wire t17303 = t17302 ^ t17302;
    wire t17304 = t17303 ^ t17303;
    wire t17305 = t17304 ^ t17304;
    wire t17306 = t17305 ^ t17305;
    wire t17307 = t17306 ^ t17306;
    wire t17308 = t17307 ^ t17307;
    wire t17309 = t17308 ^ t17308;
    wire t17310 = t17309 ^ t17309;
    wire t17311 = t17310 ^ t17310;
    wire t17312 = t17311 ^ t17311;
    wire t17313 = t17312 ^ t17312;
    wire t17314 = t17313 ^ t17313;
    wire t17315 = t17314 ^ t17314;
    wire t17316 = t17315 ^ t17315;
    wire t17317 = t17316 ^ t17316;
    wire t17318 = t17317 ^ t17317;
    wire t17319 = t17318 ^ t17318;
    wire t17320 = t17319 ^ t17319;
    wire t17321 = t17320 ^ t17320;
    wire t17322 = t17321 ^ t17321;
    wire t17323 = t17322 ^ t17322;
    wire t17324 = t17323 ^ t17323;
    wire t17325 = t17324 ^ t17324;
    wire t17326 = t17325 ^ t17325;
    wire t17327 = t17326 ^ t17326;
    wire t17328 = t17327 ^ t17327;
    wire t17329 = t17328 ^ t17328;
    wire t17330 = t17329 ^ t17329;
    wire t17331 = t17330 ^ t17330;
    wire t17332 = t17331 ^ t17331;
    wire t17333 = t17332 ^ t17332;
    wire t17334 = t17333 ^ t17333;
    wire t17335 = t17334 ^ t17334;
    wire t17336 = t17335 ^ t17335;
    wire t17337 = t17336 ^ t17336;
    wire t17338 = t17337 ^ t17337;
    wire t17339 = t17338 ^ t17338;
    wire t17340 = t17339 ^ t17339;
    wire t17341 = t17340 ^ t17340;
    wire t17342 = t17341 ^ t17341;
    wire t17343 = t17342 ^ t17342;
    wire t17344 = t17343 ^ t17343;
    wire t17345 = t17344 ^ t17344;
    wire t17346 = t17345 ^ t17345;
    wire t17347 = t17346 ^ t17346;
    wire t17348 = t17347 ^ t17347;
    wire t17349 = t17348 ^ t17348;
    wire t17350 = t17349 ^ t17349;
    wire t17351 = t17350 ^ t17350;
    wire t17352 = t17351 ^ t17351;
    wire t17353 = t17352 ^ t17352;
    wire t17354 = t17353 ^ t17353;
    wire t17355 = t17354 ^ t17354;
    wire t17356 = t17355 ^ t17355;
    wire t17357 = t17356 ^ t17356;
    wire t17358 = t17357 ^ t17357;
    wire t17359 = t17358 ^ t17358;
    wire t17360 = t17359 ^ t17359;
    wire t17361 = t17360 ^ t17360;
    wire t17362 = t17361 ^ t17361;
    wire t17363 = t17362 ^ t17362;
    wire t17364 = t17363 ^ t17363;
    wire t17365 = t17364 ^ t17364;
    wire t17366 = t17365 ^ t17365;
    wire t17367 = t17366 ^ t17366;
    wire t17368 = t17367 ^ t17367;
    wire t17369 = t17368 ^ t17368;
    wire t17370 = t17369 ^ t17369;
    wire t17371 = t17370 ^ t17370;
    wire t17372 = t17371 ^ t17371;
    wire t17373 = t17372 ^ t17372;
    wire t17374 = t17373 ^ t17373;
    wire t17375 = t17374 ^ t17374;
    wire t17376 = t17375 ^ t17375;
    wire t17377 = t17376 ^ t17376;
    wire t17378 = t17377 ^ t17377;
    wire t17379 = t17378 ^ t17378;
    wire t17380 = t17379 ^ t17379;
    wire t17381 = t17380 ^ t17380;
    wire t17382 = t17381 ^ t17381;
    wire t17383 = t17382 ^ t17382;
    wire t17384 = t17383 ^ t17383;
    wire t17385 = t17384 ^ t17384;
    wire t17386 = t17385 ^ t17385;
    wire t17387 = t17386 ^ t17386;
    wire t17388 = t17387 ^ t17387;
    wire t17389 = t17388 ^ t17388;
    wire t17390 = t17389 ^ t17389;
    wire t17391 = t17390 ^ t17390;
    wire t17392 = t17391 ^ t17391;
    wire t17393 = t17392 ^ t17392;
    wire t17394 = t17393 ^ t17393;
    wire t17395 = t17394 ^ t17394;
    wire t17396 = t17395 ^ t17395;
    wire t17397 = t17396 ^ t17396;
    wire t17398 = t17397 ^ t17397;
    wire t17399 = t17398 ^ t17398;
    wire t17400 = t17399 ^ t17399;
    wire t17401 = t17400 ^ t17400;
    wire t17402 = t17401 ^ t17401;
    wire t17403 = t17402 ^ t17402;
    wire t17404 = t17403 ^ t17403;
    wire t17405 = t17404 ^ t17404;
    wire t17406 = t17405 ^ t17405;
    wire t17407 = t17406 ^ t17406;
    wire t17408 = t17407 ^ t17407;
    wire t17409 = t17408 ^ t17408;
    wire t17410 = t17409 ^ t17409;
    wire t17411 = t17410 ^ t17410;
    wire t17412 = t17411 ^ t17411;
    wire t17413 = t17412 ^ t17412;
    wire t17414 = t17413 ^ t17413;
    wire t17415 = t17414 ^ t17414;
    wire t17416 = t17415 ^ t17415;
    wire t17417 = t17416 ^ t17416;
    wire t17418 = t17417 ^ t17417;
    wire t17419 = t17418 ^ t17418;
    wire t17420 = t17419 ^ t17419;
    wire t17421 = t17420 ^ t17420;
    wire t17422 = t17421 ^ t17421;
    wire t17423 = t17422 ^ t17422;
    wire t17424 = t17423 ^ t17423;
    wire t17425 = t17424 ^ t17424;
    wire t17426 = t17425 ^ t17425;
    wire t17427 = t17426 ^ t17426;
    wire t17428 = t17427 ^ t17427;
    wire t17429 = t17428 ^ t17428;
    wire t17430 = t17429 ^ t17429;
    wire t17431 = t17430 ^ t17430;
    wire t17432 = t17431 ^ t17431;
    wire t17433 = t17432 ^ t17432;
    wire t17434 = t17433 ^ t17433;
    wire t17435 = t17434 ^ t17434;
    wire t17436 = t17435 ^ t17435;
    wire t17437 = t17436 ^ t17436;
    wire t17438 = t17437 ^ t17437;
    wire t17439 = t17438 ^ t17438;
    wire t17440 = t17439 ^ t17439;
    wire t17441 = t17440 ^ t17440;
    wire t17442 = t17441 ^ t17441;
    wire t17443 = t17442 ^ t17442;
    wire t17444 = t17443 ^ t17443;
    wire t17445 = t17444 ^ t17444;
    wire t17446 = t17445 ^ t17445;
    wire t17447 = t17446 ^ t17446;
    wire t17448 = t17447 ^ t17447;
    wire t17449 = t17448 ^ t17448;
    wire t17450 = t17449 ^ t17449;
    wire t17451 = t17450 ^ t17450;
    wire t17452 = t17451 ^ t17451;
    wire t17453 = t17452 ^ t17452;
    wire t17454 = t17453 ^ t17453;
    wire t17455 = t17454 ^ t17454;
    wire t17456 = t17455 ^ t17455;
    wire t17457 = t17456 ^ t17456;
    wire t17458 = t17457 ^ t17457;
    wire t17459 = t17458 ^ t17458;
    wire t17460 = t17459 ^ t17459;
    wire t17461 = t17460 ^ t17460;
    wire t17462 = t17461 ^ t17461;
    wire t17463 = t17462 ^ t17462;
    wire t17464 = t17463 ^ t17463;
    wire t17465 = t17464 ^ t17464;
    wire t17466 = t17465 ^ t17465;
    wire t17467 = t17466 ^ t17466;
    wire t17468 = t17467 ^ t17467;
    wire t17469 = t17468 ^ t17468;
    wire t17470 = t17469 ^ t17469;
    wire t17471 = t17470 ^ t17470;
    wire t17472 = t17471 ^ t17471;
    wire t17473 = t17472 ^ t17472;
    wire t17474 = t17473 ^ t17473;
    wire t17475 = t17474 ^ t17474;
    wire t17476 = t17475 ^ t17475;
    wire t17477 = t17476 ^ t17476;
    wire t17478 = t17477 ^ t17477;
    wire t17479 = t17478 ^ t17478;
    wire t17480 = t17479 ^ t17479;
    wire t17481 = t17480 ^ t17480;
    wire t17482 = t17481 ^ t17481;
    wire t17483 = t17482 ^ t17482;
    wire t17484 = t17483 ^ t17483;
    wire t17485 = t17484 ^ t17484;
    wire t17486 = t17485 ^ t17485;
    wire t17487 = t17486 ^ t17486;
    wire t17488 = t17487 ^ t17487;
    wire t17489 = t17488 ^ t17488;
    wire t17490 = t17489 ^ t17489;
    wire t17491 = t17490 ^ t17490;
    wire t17492 = t17491 ^ t17491;
    wire t17493 = t17492 ^ t17492;
    wire t17494 = t17493 ^ t17493;
    wire t17495 = t17494 ^ t17494;
    wire t17496 = t17495 ^ t17495;
    wire t17497 = t17496 ^ t17496;
    wire t17498 = t17497 ^ t17497;
    wire t17499 = t17498 ^ t17498;
    wire t17500 = t17499 ^ t17499;
    wire t17501 = t17500 ^ t17500;
    wire t17502 = t17501 ^ t17501;
    wire t17503 = t17502 ^ t17502;
    wire t17504 = t17503 ^ t17503;
    wire t17505 = t17504 ^ t17504;
    wire t17506 = t17505 ^ t17505;
    wire t17507 = t17506 ^ t17506;
    wire t17508 = t17507 ^ t17507;
    wire t17509 = t17508 ^ t17508;
    wire t17510 = t17509 ^ t17509;
    wire t17511 = t17510 ^ t17510;
    wire t17512 = t17511 ^ t17511;
    wire t17513 = t17512 ^ t17512;
    wire t17514 = t17513 ^ t17513;
    wire t17515 = t17514 ^ t17514;
    wire t17516 = t17515 ^ t17515;
    wire t17517 = t17516 ^ t17516;
    wire t17518 = t17517 ^ t17517;
    wire t17519 = t17518 ^ t17518;
    wire t17520 = t17519 ^ t17519;
    wire t17521 = t17520 ^ t17520;
    wire t17522 = t17521 ^ t17521;
    wire t17523 = t17522 ^ t17522;
    wire t17524 = t17523 ^ t17523;
    wire t17525 = t17524 ^ t17524;
    wire t17526 = t17525 ^ t17525;
    wire t17527 = t17526 ^ t17526;
    wire t17528 = t17527 ^ t17527;
    wire t17529 = t17528 ^ t17528;
    wire t17530 = t17529 ^ t17529;
    wire t17531 = t17530 ^ t17530;
    wire t17532 = t17531 ^ t17531;
    wire t17533 = t17532 ^ t17532;
    wire t17534 = t17533 ^ t17533;
    wire t17535 = t17534 ^ t17534;
    wire t17536 = t17535 ^ t17535;
    wire t17537 = t17536 ^ t17536;
    wire t17538 = t17537 ^ t17537;
    wire t17539 = t17538 ^ t17538;
    wire t17540 = t17539 ^ t17539;
    wire t17541 = t17540 ^ t17540;
    wire t17542 = t17541 ^ t17541;
    wire t17543 = t17542 ^ t17542;
    wire t17544 = t17543 ^ t17543;
    wire t17545 = t17544 ^ t17544;
    wire t17546 = t17545 ^ t17545;
    wire t17547 = t17546 ^ t17546;
    wire t17548 = t17547 ^ t17547;
    wire t17549 = t17548 ^ t17548;
    wire t17550 = t17549 ^ t17549;
    wire t17551 = t17550 ^ t17550;
    wire t17552 = t17551 ^ t17551;
    wire t17553 = t17552 ^ t17552;
    wire t17554 = t17553 ^ t17553;
    wire t17555 = t17554 ^ t17554;
    wire t17556 = t17555 ^ t17555;
    wire t17557 = t17556 ^ t17556;
    wire t17558 = t17557 ^ t17557;
    wire t17559 = t17558 ^ t17558;
    wire t17560 = t17559 ^ t17559;
    wire t17561 = t17560 ^ t17560;
    wire t17562 = t17561 ^ t17561;
    wire t17563 = t17562 ^ t17562;
    wire t17564 = t17563 ^ t17563;
    wire t17565 = t17564 ^ t17564;
    wire t17566 = t17565 ^ t17565;
    wire t17567 = t17566 ^ t17566;
    wire t17568 = t17567 ^ t17567;
    wire t17569 = t17568 ^ t17568;
    wire t17570 = t17569 ^ t17569;
    wire t17571 = t17570 ^ t17570;
    wire t17572 = t17571 ^ t17571;
    wire t17573 = t17572 ^ t17572;
    wire t17574 = t17573 ^ t17573;
    wire t17575 = t17574 ^ t17574;
    wire t17576 = t17575 ^ t17575;
    wire t17577 = t17576 ^ t17576;
    wire t17578 = t17577 ^ t17577;
    wire t17579 = t17578 ^ t17578;
    wire t17580 = t17579 ^ t17579;
    wire t17581 = t17580 ^ t17580;
    wire t17582 = t17581 ^ t17581;
    wire t17583 = t17582 ^ t17582;
    wire t17584 = t17583 ^ t17583;
    wire t17585 = t17584 ^ t17584;
    wire t17586 = t17585 ^ t17585;
    wire t17587 = t17586 ^ t17586;
    wire t17588 = t17587 ^ t17587;
    wire t17589 = t17588 ^ t17588;
    wire t17590 = t17589 ^ t17589;
    wire t17591 = t17590 ^ t17590;
    wire t17592 = t17591 ^ t17591;
    wire t17593 = t17592 ^ t17592;
    wire t17594 = t17593 ^ t17593;
    wire t17595 = t17594 ^ t17594;
    wire t17596 = t17595 ^ t17595;
    wire t17597 = t17596 ^ t17596;
    wire t17598 = t17597 ^ t17597;
    wire t17599 = t17598 ^ t17598;
    wire t17600 = t17599 ^ t17599;
    wire t17601 = t17600 ^ t17600;
    wire t17602 = t17601 ^ t17601;
    wire t17603 = t17602 ^ t17602;
    wire t17604 = t17603 ^ t17603;
    wire t17605 = t17604 ^ t17604;
    wire t17606 = t17605 ^ t17605;
    wire t17607 = t17606 ^ t17606;
    wire t17608 = t17607 ^ t17607;
    wire t17609 = t17608 ^ t17608;
    wire t17610 = t17609 ^ t17609;
    wire t17611 = t17610 ^ t17610;
    wire t17612 = t17611 ^ t17611;
    wire t17613 = t17612 ^ t17612;
    wire t17614 = t17613 ^ t17613;
    wire t17615 = t17614 ^ t17614;
    wire t17616 = t17615 ^ t17615;
    wire t17617 = t17616 ^ t17616;
    wire t17618 = t17617 ^ t17617;
    wire t17619 = t17618 ^ t17618;
    wire t17620 = t17619 ^ t17619;
    wire t17621 = t17620 ^ t17620;
    wire t17622 = t17621 ^ t17621;
    wire t17623 = t17622 ^ t17622;
    wire t17624 = t17623 ^ t17623;
    wire t17625 = t17624 ^ t17624;
    wire t17626 = t17625 ^ t17625;
    wire t17627 = t17626 ^ t17626;
    wire t17628 = t17627 ^ t17627;
    wire t17629 = t17628 ^ t17628;
    wire t17630 = t17629 ^ t17629;
    wire t17631 = t17630 ^ t17630;
    wire t17632 = t17631 ^ t17631;
    wire t17633 = t17632 ^ t17632;
    wire t17634 = t17633 ^ t17633;
    wire t17635 = t17634 ^ t17634;
    wire t17636 = t17635 ^ t17635;
    wire t17637 = t17636 ^ t17636;
    wire t17638 = t17637 ^ t17637;
    wire t17639 = t17638 ^ t17638;
    wire t17640 = t17639 ^ t17639;
    wire t17641 = t17640 ^ t17640;
    wire t17642 = t17641 ^ t17641;
    wire t17643 = t17642 ^ t17642;
    wire t17644 = t17643 ^ t17643;
    wire t17645 = t17644 ^ t17644;
    wire t17646 = t17645 ^ t17645;
    wire t17647 = t17646 ^ t17646;
    wire t17648 = t17647 ^ t17647;
    wire t17649 = t17648 ^ t17648;
    wire t17650 = t17649 ^ t17649;
    wire t17651 = t17650 ^ t17650;
    wire t17652 = t17651 ^ t17651;
    wire t17653 = t17652 ^ t17652;
    wire t17654 = t17653 ^ t17653;
    wire t17655 = t17654 ^ t17654;
    wire t17656 = t17655 ^ t17655;
    wire t17657 = t17656 ^ t17656;
    wire t17658 = t17657 ^ t17657;
    wire t17659 = t17658 ^ t17658;
    wire t17660 = t17659 ^ t17659;
    wire t17661 = t17660 ^ t17660;
    wire t17662 = t17661 ^ t17661;
    wire t17663 = t17662 ^ t17662;
    wire t17664 = t17663 ^ t17663;
    wire t17665 = t17664 ^ t17664;
    wire t17666 = t17665 ^ t17665;
    wire t17667 = t17666 ^ t17666;
    wire t17668 = t17667 ^ t17667;
    wire t17669 = t17668 ^ t17668;
    wire t17670 = t17669 ^ t17669;
    wire t17671 = t17670 ^ t17670;
    wire t17672 = t17671 ^ t17671;
    wire t17673 = t17672 ^ t17672;
    wire t17674 = t17673 ^ t17673;
    wire t17675 = t17674 ^ t17674;
    wire t17676 = t17675 ^ t17675;
    wire t17677 = t17676 ^ t17676;
    wire t17678 = t17677 ^ t17677;
    wire t17679 = t17678 ^ t17678;
    wire t17680 = t17679 ^ t17679;
    wire t17681 = t17680 ^ t17680;
    wire t17682 = t17681 ^ t17681;
    wire t17683 = t17682 ^ t17682;
    wire t17684 = t17683 ^ t17683;
    wire t17685 = t17684 ^ t17684;
    wire t17686 = t17685 ^ t17685;
    wire t17687 = t17686 ^ t17686;
    wire t17688 = t17687 ^ t17687;
    wire t17689 = t17688 ^ t17688;
    wire t17690 = t17689 ^ t17689;
    wire t17691 = t17690 ^ t17690;
    wire t17692 = t17691 ^ t17691;
    wire t17693 = t17692 ^ t17692;
    wire t17694 = t17693 ^ t17693;
    wire t17695 = t17694 ^ t17694;
    wire t17696 = t17695 ^ t17695;
    wire t17697 = t17696 ^ t17696;
    wire t17698 = t17697 ^ t17697;
    wire t17699 = t17698 ^ t17698;
    wire t17700 = t17699 ^ t17699;
    wire t17701 = t17700 ^ t17700;
    wire t17702 = t17701 ^ t17701;
    wire t17703 = t17702 ^ t17702;
    wire t17704 = t17703 ^ t17703;
    wire t17705 = t17704 ^ t17704;
    wire t17706 = t17705 ^ t17705;
    wire t17707 = t17706 ^ t17706;
    wire t17708 = t17707 ^ t17707;
    wire t17709 = t17708 ^ t17708;
    wire t17710 = t17709 ^ t17709;
    wire t17711 = t17710 ^ t17710;
    wire t17712 = t17711 ^ t17711;
    wire t17713 = t17712 ^ t17712;
    wire t17714 = t17713 ^ t17713;
    wire t17715 = t17714 ^ t17714;
    wire t17716 = t17715 ^ t17715;
    wire t17717 = t17716 ^ t17716;
    wire t17718 = t17717 ^ t17717;
    wire t17719 = t17718 ^ t17718;
    wire t17720 = t17719 ^ t17719;
    wire t17721 = t17720 ^ t17720;
    wire t17722 = t17721 ^ t17721;
    wire t17723 = t17722 ^ t17722;
    wire t17724 = t17723 ^ t17723;
    wire t17725 = t17724 ^ t17724;
    wire t17726 = t17725 ^ t17725;
    wire t17727 = t17726 ^ t17726;
    wire t17728 = t17727 ^ t17727;
    wire t17729 = t17728 ^ t17728;
    wire t17730 = t17729 ^ t17729;
    wire t17731 = t17730 ^ t17730;
    wire t17732 = t17731 ^ t17731;
    wire t17733 = t17732 ^ t17732;
    wire t17734 = t17733 ^ t17733;
    wire t17735 = t17734 ^ t17734;
    wire t17736 = t17735 ^ t17735;
    wire t17737 = t17736 ^ t17736;
    wire t17738 = t17737 ^ t17737;
    wire t17739 = t17738 ^ t17738;
    wire t17740 = t17739 ^ t17739;
    wire t17741 = t17740 ^ t17740;
    wire t17742 = t17741 ^ t17741;
    wire t17743 = t17742 ^ t17742;
    wire t17744 = t17743 ^ t17743;
    wire t17745 = t17744 ^ t17744;
    wire t17746 = t17745 ^ t17745;
    wire t17747 = t17746 ^ t17746;
    wire t17748 = t17747 ^ t17747;
    wire t17749 = t17748 ^ t17748;
    wire t17750 = t17749 ^ t17749;
    wire t17751 = t17750 ^ t17750;
    wire t17752 = t17751 ^ t17751;
    wire t17753 = t17752 ^ t17752;
    wire t17754 = t17753 ^ t17753;
    wire t17755 = t17754 ^ t17754;
    wire t17756 = t17755 ^ t17755;
    wire t17757 = t17756 ^ t17756;
    wire t17758 = t17757 ^ t17757;
    wire t17759 = t17758 ^ t17758;
    wire t17760 = t17759 ^ t17759;
    wire t17761 = t17760 ^ t17760;
    wire t17762 = t17761 ^ t17761;
    wire t17763 = t17762 ^ t17762;
    wire t17764 = t17763 ^ t17763;
    wire t17765 = t17764 ^ t17764;
    wire t17766 = t17765 ^ t17765;
    wire t17767 = t17766 ^ t17766;
    wire t17768 = t17767 ^ t17767;
    wire t17769 = t17768 ^ t17768;
    wire t17770 = t17769 ^ t17769;
    wire t17771 = t17770 ^ t17770;
    wire t17772 = t17771 ^ t17771;
    wire t17773 = t17772 ^ t17772;
    wire t17774 = t17773 ^ t17773;
    wire t17775 = t17774 ^ t17774;
    wire t17776 = t17775 ^ t17775;
    wire t17777 = t17776 ^ t17776;
    wire t17778 = t17777 ^ t17777;
    wire t17779 = t17778 ^ t17778;
    wire t17780 = t17779 ^ t17779;
    wire t17781 = t17780 ^ t17780;
    wire t17782 = t17781 ^ t17781;
    wire t17783 = t17782 ^ t17782;
    wire t17784 = t17783 ^ t17783;
    wire t17785 = t17784 ^ t17784;
    wire t17786 = t17785 ^ t17785;
    wire t17787 = t17786 ^ t17786;
    wire t17788 = t17787 ^ t17787;
    wire t17789 = t17788 ^ t17788;
    wire t17790 = t17789 ^ t17789;
    wire t17791 = t17790 ^ t17790;
    wire t17792 = t17791 ^ t17791;
    wire t17793 = t17792 ^ t17792;
    wire t17794 = t17793 ^ t17793;
    wire t17795 = t17794 ^ t17794;
    wire t17796 = t17795 ^ t17795;
    wire t17797 = t17796 ^ t17796;
    wire t17798 = t17797 ^ t17797;
    wire t17799 = t17798 ^ t17798;
    wire t17800 = t17799 ^ t17799;
    wire t17801 = t17800 ^ t17800;
    wire t17802 = t17801 ^ t17801;
    wire t17803 = t17802 ^ t17802;
    wire t17804 = t17803 ^ t17803;
    wire t17805 = t17804 ^ t17804;
    wire t17806 = t17805 ^ t17805;
    wire t17807 = t17806 ^ t17806;
    wire t17808 = t17807 ^ t17807;
    wire t17809 = t17808 ^ t17808;
    wire t17810 = t17809 ^ t17809;
    wire t17811 = t17810 ^ t17810;
    wire t17812 = t17811 ^ t17811;
    wire t17813 = t17812 ^ t17812;
    wire t17814 = t17813 ^ t17813;
    wire t17815 = t17814 ^ t17814;
    wire t17816 = t17815 ^ t17815;
    wire t17817 = t17816 ^ t17816;
    wire t17818 = t17817 ^ t17817;
    wire t17819 = t17818 ^ t17818;
    wire t17820 = t17819 ^ t17819;
    wire t17821 = t17820 ^ t17820;
    wire t17822 = t17821 ^ t17821;
    wire t17823 = t17822 ^ t17822;
    wire t17824 = t17823 ^ t17823;
    wire t17825 = t17824 ^ t17824;
    wire t17826 = t17825 ^ t17825;
    wire t17827 = t17826 ^ t17826;
    wire t17828 = t17827 ^ t17827;
    wire t17829 = t17828 ^ t17828;
    wire t17830 = t17829 ^ t17829;
    wire t17831 = t17830 ^ t17830;
    wire t17832 = t17831 ^ t17831;
    wire t17833 = t17832 ^ t17832;
    wire t17834 = t17833 ^ t17833;
    wire t17835 = t17834 ^ t17834;
    wire t17836 = t17835 ^ t17835;
    wire t17837 = t17836 ^ t17836;
    wire t17838 = t17837 ^ t17837;
    wire t17839 = t17838 ^ t17838;
    wire t17840 = t17839 ^ t17839;
    wire t17841 = t17840 ^ t17840;
    wire t17842 = t17841 ^ t17841;
    wire t17843 = t17842 ^ t17842;
    wire t17844 = t17843 ^ t17843;
    wire t17845 = t17844 ^ t17844;
    wire t17846 = t17845 ^ t17845;
    wire t17847 = t17846 ^ t17846;
    wire t17848 = t17847 ^ t17847;
    wire t17849 = t17848 ^ t17848;
    wire t17850 = t17849 ^ t17849;
    wire t17851 = t17850 ^ t17850;
    wire t17852 = t17851 ^ t17851;
    wire t17853 = t17852 ^ t17852;
    wire t17854 = t17853 ^ t17853;
    wire t17855 = t17854 ^ t17854;
    wire t17856 = t17855 ^ t17855;
    wire t17857 = t17856 ^ t17856;
    wire t17858 = t17857 ^ t17857;
    wire t17859 = t17858 ^ t17858;
    wire t17860 = t17859 ^ t17859;
    wire t17861 = t17860 ^ t17860;
    wire t17862 = t17861 ^ t17861;
    wire t17863 = t17862 ^ t17862;
    wire t17864 = t17863 ^ t17863;
    wire t17865 = t17864 ^ t17864;
    wire t17866 = t17865 ^ t17865;
    wire t17867 = t17866 ^ t17866;
    wire t17868 = t17867 ^ t17867;
    wire t17869 = t17868 ^ t17868;
    wire t17870 = t17869 ^ t17869;
    wire t17871 = t17870 ^ t17870;
    wire t17872 = t17871 ^ t17871;
    wire t17873 = t17872 ^ t17872;
    wire t17874 = t17873 ^ t17873;
    wire t17875 = t17874 ^ t17874;
    wire t17876 = t17875 ^ t17875;
    wire t17877 = t17876 ^ t17876;
    wire t17878 = t17877 ^ t17877;
    wire t17879 = t17878 ^ t17878;
    wire t17880 = t17879 ^ t17879;
    wire t17881 = t17880 ^ t17880;
    wire t17882 = t17881 ^ t17881;
    wire t17883 = t17882 ^ t17882;
    wire t17884 = t17883 ^ t17883;
    wire t17885 = t17884 ^ t17884;
    wire t17886 = t17885 ^ t17885;
    wire t17887 = t17886 ^ t17886;
    wire t17888 = t17887 ^ t17887;
    wire t17889 = t17888 ^ t17888;
    wire t17890 = t17889 ^ t17889;
    wire t17891 = t17890 ^ t17890;
    wire t17892 = t17891 ^ t17891;
    wire t17893 = t17892 ^ t17892;
    wire t17894 = t17893 ^ t17893;
    wire t17895 = t17894 ^ t17894;
    wire t17896 = t17895 ^ t17895;
    wire t17897 = t17896 ^ t17896;
    wire t17898 = t17897 ^ t17897;
    wire t17899 = t17898 ^ t17898;
    wire t17900 = t17899 ^ t17899;
    wire t17901 = t17900 ^ t17900;
    wire t17902 = t17901 ^ t17901;
    wire t17903 = t17902 ^ t17902;
    wire t17904 = t17903 ^ t17903;
    wire t17905 = t17904 ^ t17904;
    wire t17906 = t17905 ^ t17905;
    wire t17907 = t17906 ^ t17906;
    wire t17908 = t17907 ^ t17907;
    wire t17909 = t17908 ^ t17908;
    wire t17910 = t17909 ^ t17909;
    wire t17911 = t17910 ^ t17910;
    wire t17912 = t17911 ^ t17911;
    wire t17913 = t17912 ^ t17912;
    wire t17914 = t17913 ^ t17913;
    wire t17915 = t17914 ^ t17914;
    wire t17916 = t17915 ^ t17915;
    wire t17917 = t17916 ^ t17916;
    wire t17918 = t17917 ^ t17917;
    wire t17919 = t17918 ^ t17918;
    wire t17920 = t17919 ^ t17919;
    wire t17921 = t17920 ^ t17920;
    wire t17922 = t17921 ^ t17921;
    wire t17923 = t17922 ^ t17922;
    wire t17924 = t17923 ^ t17923;
    wire t17925 = t17924 ^ t17924;
    wire t17926 = t17925 ^ t17925;
    wire t17927 = t17926 ^ t17926;
    wire t17928 = t17927 ^ t17927;
    wire t17929 = t17928 ^ t17928;
    wire t17930 = t17929 ^ t17929;
    wire t17931 = t17930 ^ t17930;
    wire t17932 = t17931 ^ t17931;
    wire t17933 = t17932 ^ t17932;
    wire t17934 = t17933 ^ t17933;
    wire t17935 = t17934 ^ t17934;
    wire t17936 = t17935 ^ t17935;
    wire t17937 = t17936 ^ t17936;
    wire t17938 = t17937 ^ t17937;
    wire t17939 = t17938 ^ t17938;
    wire t17940 = t17939 ^ t17939;
    wire t17941 = t17940 ^ t17940;
    wire t17942 = t17941 ^ t17941;
    wire t17943 = t17942 ^ t17942;
    wire t17944 = t17943 ^ t17943;
    wire t17945 = t17944 ^ t17944;
    wire t17946 = t17945 ^ t17945;
    wire t17947 = t17946 ^ t17946;
    wire t17948 = t17947 ^ t17947;
    wire t17949 = t17948 ^ t17948;
    wire t17950 = t17949 ^ t17949;
    wire t17951 = t17950 ^ t17950;
    wire t17952 = t17951 ^ t17951;
    wire t17953 = t17952 ^ t17952;
    wire t17954 = t17953 ^ t17953;
    wire t17955 = t17954 ^ t17954;
    wire t17956 = t17955 ^ t17955;
    wire t17957 = t17956 ^ t17956;
    wire t17958 = t17957 ^ t17957;
    wire t17959 = t17958 ^ t17958;
    wire t17960 = t17959 ^ t17959;
    wire t17961 = t17960 ^ t17960;
    wire t17962 = t17961 ^ t17961;
    wire t17963 = t17962 ^ t17962;
    wire t17964 = t17963 ^ t17963;
    wire t17965 = t17964 ^ t17964;
    wire t17966 = t17965 ^ t17965;
    wire t17967 = t17966 ^ t17966;
    wire t17968 = t17967 ^ t17967;
    wire t17969 = t17968 ^ t17968;
    wire t17970 = t17969 ^ t17969;
    wire t17971 = t17970 ^ t17970;
    wire t17972 = t17971 ^ t17971;
    wire t17973 = t17972 ^ t17972;
    wire t17974 = t17973 ^ t17973;
    wire t17975 = t17974 ^ t17974;
    wire t17976 = t17975 ^ t17975;
    wire t17977 = t17976 ^ t17976;
    wire t17978 = t17977 ^ t17977;
    wire t17979 = t17978 ^ t17978;
    wire t17980 = t17979 ^ t17979;
    wire t17981 = t17980 ^ t17980;
    wire t17982 = t17981 ^ t17981;
    wire t17983 = t17982 ^ t17982;
    wire t17984 = t17983 ^ t17983;
    wire t17985 = t17984 ^ t17984;
    wire t17986 = t17985 ^ t17985;
    wire t17987 = t17986 ^ t17986;
    wire t17988 = t17987 ^ t17987;
    wire t17989 = t17988 ^ t17988;
    wire t17990 = t17989 ^ t17989;
    wire t17991 = t17990 ^ t17990;
    wire t17992 = t17991 ^ t17991;
    wire t17993 = t17992 ^ t17992;
    wire t17994 = t17993 ^ t17993;
    wire t17995 = t17994 ^ t17994;
    wire t17996 = t17995 ^ t17995;
    wire t17997 = t17996 ^ t17996;
    wire t17998 = t17997 ^ t17997;
    wire t17999 = t17998 ^ t17998;
    wire t18000 = t17999 ^ t17999;
    wire t18001 = t18000 ^ t18000;
    wire t18002 = t18001 ^ t18001;
    wire t18003 = t18002 ^ t18002;
    wire t18004 = t18003 ^ t18003;
    wire t18005 = t18004 ^ t18004;
    wire t18006 = t18005 ^ t18005;
    wire t18007 = t18006 ^ t18006;
    wire t18008 = t18007 ^ t18007;
    wire t18009 = t18008 ^ t18008;
    wire t18010 = t18009 ^ t18009;
    wire t18011 = t18010 ^ t18010;
    wire t18012 = t18011 ^ t18011;
    wire t18013 = t18012 ^ t18012;
    wire t18014 = t18013 ^ t18013;
    wire t18015 = t18014 ^ t18014;
    wire t18016 = t18015 ^ t18015;
    wire t18017 = t18016 ^ t18016;
    wire t18018 = t18017 ^ t18017;
    wire t18019 = t18018 ^ t18018;
    wire t18020 = t18019 ^ t18019;
    wire t18021 = t18020 ^ t18020;
    wire t18022 = t18021 ^ t18021;
    wire t18023 = t18022 ^ t18022;
    wire t18024 = t18023 ^ t18023;
    wire t18025 = t18024 ^ t18024;
    wire t18026 = t18025 ^ t18025;
    wire t18027 = t18026 ^ t18026;
    wire t18028 = t18027 ^ t18027;
    wire t18029 = t18028 ^ t18028;
    wire t18030 = t18029 ^ t18029;
    wire t18031 = t18030 ^ t18030;
    wire t18032 = t18031 ^ t18031;
    wire t18033 = t18032 ^ t18032;
    wire t18034 = t18033 ^ t18033;
    wire t18035 = t18034 ^ t18034;
    wire t18036 = t18035 ^ t18035;
    wire t18037 = t18036 ^ t18036;
    wire t18038 = t18037 ^ t18037;
    wire t18039 = t18038 ^ t18038;
    wire t18040 = t18039 ^ t18039;
    wire t18041 = t18040 ^ t18040;
    wire t18042 = t18041 ^ t18041;
    wire t18043 = t18042 ^ t18042;
    wire t18044 = t18043 ^ t18043;
    wire t18045 = t18044 ^ t18044;
    wire t18046 = t18045 ^ t18045;
    wire t18047 = t18046 ^ t18046;
    wire t18048 = t18047 ^ t18047;
    wire t18049 = t18048 ^ t18048;
    wire t18050 = t18049 ^ t18049;
    wire t18051 = t18050 ^ t18050;
    wire t18052 = t18051 ^ t18051;
    wire t18053 = t18052 ^ t18052;
    wire t18054 = t18053 ^ t18053;
    wire t18055 = t18054 ^ t18054;
    wire t18056 = t18055 ^ t18055;
    wire t18057 = t18056 ^ t18056;
    wire t18058 = t18057 ^ t18057;
    wire t18059 = t18058 ^ t18058;
    wire t18060 = t18059 ^ t18059;
    wire t18061 = t18060 ^ t18060;
    wire t18062 = t18061 ^ t18061;
    wire t18063 = t18062 ^ t18062;
    wire t18064 = t18063 ^ t18063;
    wire t18065 = t18064 ^ t18064;
    wire t18066 = t18065 ^ t18065;
    wire t18067 = t18066 ^ t18066;
    wire t18068 = t18067 ^ t18067;
    wire t18069 = t18068 ^ t18068;
    wire t18070 = t18069 ^ t18069;
    wire t18071 = t18070 ^ t18070;
    wire t18072 = t18071 ^ t18071;
    wire t18073 = t18072 ^ t18072;
    wire t18074 = t18073 ^ t18073;
    wire t18075 = t18074 ^ t18074;
    wire t18076 = t18075 ^ t18075;
    wire t18077 = t18076 ^ t18076;
    wire t18078 = t18077 ^ t18077;
    wire t18079 = t18078 ^ t18078;
    wire t18080 = t18079 ^ t18079;
    wire t18081 = t18080 ^ t18080;
    wire t18082 = t18081 ^ t18081;
    wire t18083 = t18082 ^ t18082;
    wire t18084 = t18083 ^ t18083;
    wire t18085 = t18084 ^ t18084;
    wire t18086 = t18085 ^ t18085;
    wire t18087 = t18086 ^ t18086;
    wire t18088 = t18087 ^ t18087;
    wire t18089 = t18088 ^ t18088;
    wire t18090 = t18089 ^ t18089;
    wire t18091 = t18090 ^ t18090;
    wire t18092 = t18091 ^ t18091;
    wire t18093 = t18092 ^ t18092;
    wire t18094 = t18093 ^ t18093;
    wire t18095 = t18094 ^ t18094;
    wire t18096 = t18095 ^ t18095;
    wire t18097 = t18096 ^ t18096;
    wire t18098 = t18097 ^ t18097;
    wire t18099 = t18098 ^ t18098;
    wire t18100 = t18099 ^ t18099;
    wire t18101 = t18100 ^ t18100;
    wire t18102 = t18101 ^ t18101;
    wire t18103 = t18102 ^ t18102;
    wire t18104 = t18103 ^ t18103;
    wire t18105 = t18104 ^ t18104;
    wire t18106 = t18105 ^ t18105;
    wire t18107 = t18106 ^ t18106;
    wire t18108 = t18107 ^ t18107;
    wire t18109 = t18108 ^ t18108;
    wire t18110 = t18109 ^ t18109;
    wire t18111 = t18110 ^ t18110;
    wire t18112 = t18111 ^ t18111;
    wire t18113 = t18112 ^ t18112;
    wire t18114 = t18113 ^ t18113;
    wire t18115 = t18114 ^ t18114;
    wire t18116 = t18115 ^ t18115;
    wire t18117 = t18116 ^ t18116;
    wire t18118 = t18117 ^ t18117;
    wire t18119 = t18118 ^ t18118;
    wire t18120 = t18119 ^ t18119;
    wire t18121 = t18120 ^ t18120;
    wire t18122 = t18121 ^ t18121;
    wire t18123 = t18122 ^ t18122;
    wire t18124 = t18123 ^ t18123;
    wire t18125 = t18124 ^ t18124;
    wire t18126 = t18125 ^ t18125;
    wire t18127 = t18126 ^ t18126;
    wire t18128 = t18127 ^ t18127;
    wire t18129 = t18128 ^ t18128;
    wire t18130 = t18129 ^ t18129;
    wire t18131 = t18130 ^ t18130;
    wire t18132 = t18131 ^ t18131;
    wire t18133 = t18132 ^ t18132;
    wire t18134 = t18133 ^ t18133;
    wire t18135 = t18134 ^ t18134;
    wire t18136 = t18135 ^ t18135;
    wire t18137 = t18136 ^ t18136;
    wire t18138 = t18137 ^ t18137;
    wire t18139 = t18138 ^ t18138;
    wire t18140 = t18139 ^ t18139;
    wire t18141 = t18140 ^ t18140;
    wire t18142 = t18141 ^ t18141;
    wire t18143 = t18142 ^ t18142;
    wire t18144 = t18143 ^ t18143;
    wire t18145 = t18144 ^ t18144;
    wire t18146 = t18145 ^ t18145;
    wire t18147 = t18146 ^ t18146;
    wire t18148 = t18147 ^ t18147;
    wire t18149 = t18148 ^ t18148;
    wire t18150 = t18149 ^ t18149;
    wire t18151 = t18150 ^ t18150;
    wire t18152 = t18151 ^ t18151;
    wire t18153 = t18152 ^ t18152;
    wire t18154 = t18153 ^ t18153;
    wire t18155 = t18154 ^ t18154;
    wire t18156 = t18155 ^ t18155;
    wire t18157 = t18156 ^ t18156;
    wire t18158 = t18157 ^ t18157;
    wire t18159 = t18158 ^ t18158;
    wire t18160 = t18159 ^ t18159;
    wire t18161 = t18160 ^ t18160;
    wire t18162 = t18161 ^ t18161;
    wire t18163 = t18162 ^ t18162;
    wire t18164 = t18163 ^ t18163;
    wire t18165 = t18164 ^ t18164;
    wire t18166 = t18165 ^ t18165;
    wire t18167 = t18166 ^ t18166;
    wire t18168 = t18167 ^ t18167;
    wire t18169 = t18168 ^ t18168;
    wire t18170 = t18169 ^ t18169;
    wire t18171 = t18170 ^ t18170;
    wire t18172 = t18171 ^ t18171;
    wire t18173 = t18172 ^ t18172;
    wire t18174 = t18173 ^ t18173;
    wire t18175 = t18174 ^ t18174;
    wire t18176 = t18175 ^ t18175;
    wire t18177 = t18176 ^ t18176;
    wire t18178 = t18177 ^ t18177;
    wire t18179 = t18178 ^ t18178;
    wire t18180 = t18179 ^ t18179;
    wire t18181 = t18180 ^ t18180;
    wire t18182 = t18181 ^ t18181;
    wire t18183 = t18182 ^ t18182;
    wire t18184 = t18183 ^ t18183;
    wire t18185 = t18184 ^ t18184;
    wire t18186 = t18185 ^ t18185;
    wire t18187 = t18186 ^ t18186;
    wire t18188 = t18187 ^ t18187;
    wire t18189 = t18188 ^ t18188;
    wire t18190 = t18189 ^ t18189;
    wire t18191 = t18190 ^ t18190;
    wire t18192 = t18191 ^ t18191;
    wire t18193 = t18192 ^ t18192;
    wire t18194 = t18193 ^ t18193;
    wire t18195 = t18194 ^ t18194;
    wire t18196 = t18195 ^ t18195;
    wire t18197 = t18196 ^ t18196;
    wire t18198 = t18197 ^ t18197;
    wire t18199 = t18198 ^ t18198;
    wire t18200 = t18199 ^ t18199;
    wire t18201 = t18200 ^ t18200;
    wire t18202 = t18201 ^ t18201;
    wire t18203 = t18202 ^ t18202;
    wire t18204 = t18203 ^ t18203;
    wire t18205 = t18204 ^ t18204;
    wire t18206 = t18205 ^ t18205;
    wire t18207 = t18206 ^ t18206;
    wire t18208 = t18207 ^ t18207;
    wire t18209 = t18208 ^ t18208;
    wire t18210 = t18209 ^ t18209;
    wire t18211 = t18210 ^ t18210;
    wire t18212 = t18211 ^ t18211;
    wire t18213 = t18212 ^ t18212;
    wire t18214 = t18213 ^ t18213;
    wire t18215 = t18214 ^ t18214;
    wire t18216 = t18215 ^ t18215;
    wire t18217 = t18216 ^ t18216;
    wire t18218 = t18217 ^ t18217;
    wire t18219 = t18218 ^ t18218;
    wire t18220 = t18219 ^ t18219;
    wire t18221 = t18220 ^ t18220;
    wire t18222 = t18221 ^ t18221;
    wire t18223 = t18222 ^ t18222;
    wire t18224 = t18223 ^ t18223;
    wire t18225 = t18224 ^ t18224;
    wire t18226 = t18225 ^ t18225;
    wire t18227 = t18226 ^ t18226;
    wire t18228 = t18227 ^ t18227;
    wire t18229 = t18228 ^ t18228;
    wire t18230 = t18229 ^ t18229;
    wire t18231 = t18230 ^ t18230;
    wire t18232 = t18231 ^ t18231;
    wire t18233 = t18232 ^ t18232;
    wire t18234 = t18233 ^ t18233;
    wire t18235 = t18234 ^ t18234;
    wire t18236 = t18235 ^ t18235;
    wire t18237 = t18236 ^ t18236;
    wire t18238 = t18237 ^ t18237;
    wire t18239 = t18238 ^ t18238;
    wire t18240 = t18239 ^ t18239;
    wire t18241 = t18240 ^ t18240;
    wire t18242 = t18241 ^ t18241;
    wire t18243 = t18242 ^ t18242;
    wire t18244 = t18243 ^ t18243;
    wire t18245 = t18244 ^ t18244;
    wire t18246 = t18245 ^ t18245;
    wire t18247 = t18246 ^ t18246;
    wire t18248 = t18247 ^ t18247;
    wire t18249 = t18248 ^ t18248;
    wire t18250 = t18249 ^ t18249;
    wire t18251 = t18250 ^ t18250;
    wire t18252 = t18251 ^ t18251;
    wire t18253 = t18252 ^ t18252;
    wire t18254 = t18253 ^ t18253;
    wire t18255 = t18254 ^ t18254;
    wire t18256 = t18255 ^ t18255;
    wire t18257 = t18256 ^ t18256;
    wire t18258 = t18257 ^ t18257;
    wire t18259 = t18258 ^ t18258;
    wire t18260 = t18259 ^ t18259;
    wire t18261 = t18260 ^ t18260;
    wire t18262 = t18261 ^ t18261;
    wire t18263 = t18262 ^ t18262;
    wire t18264 = t18263 ^ t18263;
    wire t18265 = t18264 ^ t18264;
    wire t18266 = t18265 ^ t18265;
    wire t18267 = t18266 ^ t18266;
    wire t18268 = t18267 ^ t18267;
    wire t18269 = t18268 ^ t18268;
    wire t18270 = t18269 ^ t18269;
    wire t18271 = t18270 ^ t18270;
    wire t18272 = t18271 ^ t18271;
    wire t18273 = t18272 ^ t18272;
    wire t18274 = t18273 ^ t18273;
    wire t18275 = t18274 ^ t18274;
    wire t18276 = t18275 ^ t18275;
    wire t18277 = t18276 ^ t18276;
    wire t18278 = t18277 ^ t18277;
    wire t18279 = t18278 ^ t18278;
    wire t18280 = t18279 ^ t18279;
    wire t18281 = t18280 ^ t18280;
    wire t18282 = t18281 ^ t18281;
    wire t18283 = t18282 ^ t18282;
    wire t18284 = t18283 ^ t18283;
    wire t18285 = t18284 ^ t18284;
    wire t18286 = t18285 ^ t18285;
    wire t18287 = t18286 ^ t18286;
    wire t18288 = t18287 ^ t18287;
    wire t18289 = t18288 ^ t18288;
    wire t18290 = t18289 ^ t18289;
    wire t18291 = t18290 ^ t18290;
    wire t18292 = t18291 ^ t18291;
    wire t18293 = t18292 ^ t18292;
    wire t18294 = t18293 ^ t18293;
    wire t18295 = t18294 ^ t18294;
    wire t18296 = t18295 ^ t18295;
    wire t18297 = t18296 ^ t18296;
    wire t18298 = t18297 ^ t18297;
    wire t18299 = t18298 ^ t18298;
    wire t18300 = t18299 ^ t18299;
    wire t18301 = t18300 ^ t18300;
    wire t18302 = t18301 ^ t18301;
    wire t18303 = t18302 ^ t18302;
    wire t18304 = t18303 ^ t18303;
    wire t18305 = t18304 ^ t18304;
    wire t18306 = t18305 ^ t18305;
    wire t18307 = t18306 ^ t18306;
    wire t18308 = t18307 ^ t18307;
    wire t18309 = t18308 ^ t18308;
    wire t18310 = t18309 ^ t18309;
    wire t18311 = t18310 ^ t18310;
    wire t18312 = t18311 ^ t18311;
    wire t18313 = t18312 ^ t18312;
    wire t18314 = t18313 ^ t18313;
    wire t18315 = t18314 ^ t18314;
    wire t18316 = t18315 ^ t18315;
    wire t18317 = t18316 ^ t18316;
    wire t18318 = t18317 ^ t18317;
    wire t18319 = t18318 ^ t18318;
    wire t18320 = t18319 ^ t18319;
    wire t18321 = t18320 ^ t18320;
    wire t18322 = t18321 ^ t18321;
    wire t18323 = t18322 ^ t18322;
    wire t18324 = t18323 ^ t18323;
    wire t18325 = t18324 ^ t18324;
    wire t18326 = t18325 ^ t18325;
    wire t18327 = t18326 ^ t18326;
    wire t18328 = t18327 ^ t18327;
    wire t18329 = t18328 ^ t18328;
    wire t18330 = t18329 ^ t18329;
    wire t18331 = t18330 ^ t18330;
    wire t18332 = t18331 ^ t18331;
    wire t18333 = t18332 ^ t18332;
    wire t18334 = t18333 ^ t18333;
    wire t18335 = t18334 ^ t18334;
    wire t18336 = t18335 ^ t18335;
    wire t18337 = t18336 ^ t18336;
    wire t18338 = t18337 ^ t18337;
    wire t18339 = t18338 ^ t18338;
    wire t18340 = t18339 ^ t18339;
    wire t18341 = t18340 ^ t18340;
    wire t18342 = t18341 ^ t18341;
    wire t18343 = t18342 ^ t18342;
    wire t18344 = t18343 ^ t18343;
    wire t18345 = t18344 ^ t18344;
    wire t18346 = t18345 ^ t18345;
    wire t18347 = t18346 ^ t18346;
    wire t18348 = t18347 ^ t18347;
    wire t18349 = t18348 ^ t18348;
    wire t18350 = t18349 ^ t18349;
    wire t18351 = t18350 ^ t18350;
    wire t18352 = t18351 ^ t18351;
    wire t18353 = t18352 ^ t18352;
    wire t18354 = t18353 ^ t18353;
    wire t18355 = t18354 ^ t18354;
    wire t18356 = t18355 ^ t18355;
    wire t18357 = t18356 ^ t18356;
    wire t18358 = t18357 ^ t18357;
    wire t18359 = t18358 ^ t18358;
    wire t18360 = t18359 ^ t18359;
    wire t18361 = t18360 ^ t18360;
    wire t18362 = t18361 ^ t18361;
    wire t18363 = t18362 ^ t18362;
    wire t18364 = t18363 ^ t18363;
    wire t18365 = t18364 ^ t18364;
    wire t18366 = t18365 ^ t18365;
    wire t18367 = t18366 ^ t18366;
    wire t18368 = t18367 ^ t18367;
    wire t18369 = t18368 ^ t18368;
    wire t18370 = t18369 ^ t18369;
    wire t18371 = t18370 ^ t18370;
    wire t18372 = t18371 ^ t18371;
    wire t18373 = t18372 ^ t18372;
    wire t18374 = t18373 ^ t18373;
    wire t18375 = t18374 ^ t18374;
    wire t18376 = t18375 ^ t18375;
    wire t18377 = t18376 ^ t18376;
    wire t18378 = t18377 ^ t18377;
    wire t18379 = t18378 ^ t18378;
    wire t18380 = t18379 ^ t18379;
    wire t18381 = t18380 ^ t18380;
    wire t18382 = t18381 ^ t18381;
    wire t18383 = t18382 ^ t18382;
    wire t18384 = t18383 ^ t18383;
    wire t18385 = t18384 ^ t18384;
    wire t18386 = t18385 ^ t18385;
    wire t18387 = t18386 ^ t18386;
    wire t18388 = t18387 ^ t18387;
    wire t18389 = t18388 ^ t18388;
    wire t18390 = t18389 ^ t18389;
    wire t18391 = t18390 ^ t18390;
    wire t18392 = t18391 ^ t18391;
    wire t18393 = t18392 ^ t18392;
    wire t18394 = t18393 ^ t18393;
    wire t18395 = t18394 ^ t18394;
    wire t18396 = t18395 ^ t18395;
    wire t18397 = t18396 ^ t18396;
    wire t18398 = t18397 ^ t18397;
    wire t18399 = t18398 ^ t18398;
    wire t18400 = t18399 ^ t18399;
    wire t18401 = t18400 ^ t18400;
    wire t18402 = t18401 ^ t18401;
    wire t18403 = t18402 ^ t18402;
    wire t18404 = t18403 ^ t18403;
    wire t18405 = t18404 ^ t18404;
    wire t18406 = t18405 ^ t18405;
    wire t18407 = t18406 ^ t18406;
    wire t18408 = t18407 ^ t18407;
    wire t18409 = t18408 ^ t18408;
    wire t18410 = t18409 ^ t18409;
    wire t18411 = t18410 ^ t18410;
    wire t18412 = t18411 ^ t18411;
    wire t18413 = t18412 ^ t18412;
    wire t18414 = t18413 ^ t18413;
    wire t18415 = t18414 ^ t18414;
    wire t18416 = t18415 ^ t18415;
    wire t18417 = t18416 ^ t18416;
    wire t18418 = t18417 ^ t18417;
    wire t18419 = t18418 ^ t18418;
    wire t18420 = t18419 ^ t18419;
    wire t18421 = t18420 ^ t18420;
    wire t18422 = t18421 ^ t18421;
    wire t18423 = t18422 ^ t18422;
    wire t18424 = t18423 ^ t18423;
    wire t18425 = t18424 ^ t18424;
    wire t18426 = t18425 ^ t18425;
    wire t18427 = t18426 ^ t18426;
    wire t18428 = t18427 ^ t18427;
    wire t18429 = t18428 ^ t18428;
    wire t18430 = t18429 ^ t18429;
    wire t18431 = t18430 ^ t18430;
    wire t18432 = t18431 ^ t18431;
    wire t18433 = t18432 ^ t18432;
    wire t18434 = t18433 ^ t18433;
    wire t18435 = t18434 ^ t18434;
    wire t18436 = t18435 ^ t18435;
    wire t18437 = t18436 ^ t18436;
    wire t18438 = t18437 ^ t18437;
    wire t18439 = t18438 ^ t18438;
    wire t18440 = t18439 ^ t18439;
    wire t18441 = t18440 ^ t18440;
    wire t18442 = t18441 ^ t18441;
    wire t18443 = t18442 ^ t18442;
    wire t18444 = t18443 ^ t18443;
    wire t18445 = t18444 ^ t18444;
    wire t18446 = t18445 ^ t18445;
    wire t18447 = t18446 ^ t18446;
    wire t18448 = t18447 ^ t18447;
    wire t18449 = t18448 ^ t18448;
    wire t18450 = t18449 ^ t18449;
    wire t18451 = t18450 ^ t18450;
    wire t18452 = t18451 ^ t18451;
    wire t18453 = t18452 ^ t18452;
    wire t18454 = t18453 ^ t18453;
    wire t18455 = t18454 ^ t18454;
    wire t18456 = t18455 ^ t18455;
    wire t18457 = t18456 ^ t18456;
    wire t18458 = t18457 ^ t18457;
    wire t18459 = t18458 ^ t18458;
    wire t18460 = t18459 ^ t18459;
    wire t18461 = t18460 ^ t18460;
    wire t18462 = t18461 ^ t18461;
    wire t18463 = t18462 ^ t18462;
    wire t18464 = t18463 ^ t18463;
    wire t18465 = t18464 ^ t18464;
    wire t18466 = t18465 ^ t18465;
    wire t18467 = t18466 ^ t18466;
    wire t18468 = t18467 ^ t18467;
    wire t18469 = t18468 ^ t18468;
    wire t18470 = t18469 ^ t18469;
    wire t18471 = t18470 ^ t18470;
    wire t18472 = t18471 ^ t18471;
    wire t18473 = t18472 ^ t18472;
    wire t18474 = t18473 ^ t18473;
    wire t18475 = t18474 ^ t18474;
    wire t18476 = t18475 ^ t18475;
    wire t18477 = t18476 ^ t18476;
    wire t18478 = t18477 ^ t18477;
    wire t18479 = t18478 ^ t18478;
    wire t18480 = t18479 ^ t18479;
    wire t18481 = t18480 ^ t18480;
    wire t18482 = t18481 ^ t18481;
    wire t18483 = t18482 ^ t18482;
    wire t18484 = t18483 ^ t18483;
    wire t18485 = t18484 ^ t18484;
    wire t18486 = t18485 ^ t18485;
    wire t18487 = t18486 ^ t18486;
    wire t18488 = t18487 ^ t18487;
    wire t18489 = t18488 ^ t18488;
    wire t18490 = t18489 ^ t18489;
    wire t18491 = t18490 ^ t18490;
    wire t18492 = t18491 ^ t18491;
    wire t18493 = t18492 ^ t18492;
    wire t18494 = t18493 ^ t18493;
    wire t18495 = t18494 ^ t18494;
    wire t18496 = t18495 ^ t18495;
    wire t18497 = t18496 ^ t18496;
    wire t18498 = t18497 ^ t18497;
    wire t18499 = t18498 ^ t18498;
    wire t18500 = t18499 ^ t18499;
    wire t18501 = t18500 ^ t18500;
    wire t18502 = t18501 ^ t18501;
    wire t18503 = t18502 ^ t18502;
    wire t18504 = t18503 ^ t18503;
    wire t18505 = t18504 ^ t18504;
    wire t18506 = t18505 ^ t18505;
    wire t18507 = t18506 ^ t18506;
    wire t18508 = t18507 ^ t18507;
    wire t18509 = t18508 ^ t18508;
    wire t18510 = t18509 ^ t18509;
    wire t18511 = t18510 ^ t18510;
    wire t18512 = t18511 ^ t18511;
    wire t18513 = t18512 ^ t18512;
    wire t18514 = t18513 ^ t18513;
    wire t18515 = t18514 ^ t18514;
    wire t18516 = t18515 ^ t18515;
    wire t18517 = t18516 ^ t18516;
    wire t18518 = t18517 ^ t18517;
    wire t18519 = t18518 ^ t18518;
    wire t18520 = t18519 ^ t18519;
    wire t18521 = t18520 ^ t18520;
    wire t18522 = t18521 ^ t18521;
    wire t18523 = t18522 ^ t18522;
    wire t18524 = t18523 ^ t18523;
    wire t18525 = t18524 ^ t18524;
    wire t18526 = t18525 ^ t18525;
    wire t18527 = t18526 ^ t18526;
    wire t18528 = t18527 ^ t18527;
    wire t18529 = t18528 ^ t18528;
    wire t18530 = t18529 ^ t18529;
    wire t18531 = t18530 ^ t18530;
    wire t18532 = t18531 ^ t18531;
    wire t18533 = t18532 ^ t18532;
    wire t18534 = t18533 ^ t18533;
    wire t18535 = t18534 ^ t18534;
    wire t18536 = t18535 ^ t18535;
    wire t18537 = t18536 ^ t18536;
    wire t18538 = t18537 ^ t18537;
    wire t18539 = t18538 ^ t18538;
    wire t18540 = t18539 ^ t18539;
    wire t18541 = t18540 ^ t18540;
    wire t18542 = t18541 ^ t18541;
    wire t18543 = t18542 ^ t18542;
    wire t18544 = t18543 ^ t18543;
    wire t18545 = t18544 ^ t18544;
    wire t18546 = t18545 ^ t18545;
    wire t18547 = t18546 ^ t18546;
    wire t18548 = t18547 ^ t18547;
    wire t18549 = t18548 ^ t18548;
    wire t18550 = t18549 ^ t18549;
    wire t18551 = t18550 ^ t18550;
    wire t18552 = t18551 ^ t18551;
    wire t18553 = t18552 ^ t18552;
    wire t18554 = t18553 ^ t18553;
    wire t18555 = t18554 ^ t18554;
    wire t18556 = t18555 ^ t18555;
    wire t18557 = t18556 ^ t18556;
    wire t18558 = t18557 ^ t18557;
    wire t18559 = t18558 ^ t18558;
    wire t18560 = t18559 ^ t18559;
    wire t18561 = t18560 ^ t18560;
    wire t18562 = t18561 ^ t18561;
    wire t18563 = t18562 ^ t18562;
    wire t18564 = t18563 ^ t18563;
    wire t18565 = t18564 ^ t18564;
    wire t18566 = t18565 ^ t18565;
    wire t18567 = t18566 ^ t18566;
    wire t18568 = t18567 ^ t18567;
    wire t18569 = t18568 ^ t18568;
    wire t18570 = t18569 ^ t18569;
    wire t18571 = t18570 ^ t18570;
    wire t18572 = t18571 ^ t18571;
    wire t18573 = t18572 ^ t18572;
    wire t18574 = t18573 ^ t18573;
    wire t18575 = t18574 ^ t18574;
    wire t18576 = t18575 ^ t18575;
    wire t18577 = t18576 ^ t18576;
    wire t18578 = t18577 ^ t18577;
    wire t18579 = t18578 ^ t18578;
    wire t18580 = t18579 ^ t18579;
    wire t18581 = t18580 ^ t18580;
    wire t18582 = t18581 ^ t18581;
    wire t18583 = t18582 ^ t18582;
    wire t18584 = t18583 ^ t18583;
    wire t18585 = t18584 ^ t18584;
    wire t18586 = t18585 ^ t18585;
    wire t18587 = t18586 ^ t18586;
    wire t18588 = t18587 ^ t18587;
    wire t18589 = t18588 ^ t18588;
    wire t18590 = t18589 ^ t18589;
    wire t18591 = t18590 ^ t18590;
    wire t18592 = t18591 ^ t18591;
    wire t18593 = t18592 ^ t18592;
    wire t18594 = t18593 ^ t18593;
    wire t18595 = t18594 ^ t18594;
    wire t18596 = t18595 ^ t18595;
    wire t18597 = t18596 ^ t18596;
    wire t18598 = t18597 ^ t18597;
    wire t18599 = t18598 ^ t18598;
    wire t18600 = t18599 ^ t18599;
    wire t18601 = t18600 ^ t18600;
    wire t18602 = t18601 ^ t18601;
    wire t18603 = t18602 ^ t18602;
    wire t18604 = t18603 ^ t18603;
    wire t18605 = t18604 ^ t18604;
    wire t18606 = t18605 ^ t18605;
    wire t18607 = t18606 ^ t18606;
    wire t18608 = t18607 ^ t18607;
    wire t18609 = t18608 ^ t18608;
    wire t18610 = t18609 ^ t18609;
    wire t18611 = t18610 ^ t18610;
    wire t18612 = t18611 ^ t18611;
    wire t18613 = t18612 ^ t18612;
    wire t18614 = t18613 ^ t18613;
    wire t18615 = t18614 ^ t18614;
    wire t18616 = t18615 ^ t18615;
    wire t18617 = t18616 ^ t18616;
    wire t18618 = t18617 ^ t18617;
    wire t18619 = t18618 ^ t18618;
    wire t18620 = t18619 ^ t18619;
    wire t18621 = t18620 ^ t18620;
    wire t18622 = t18621 ^ t18621;
    wire t18623 = t18622 ^ t18622;
    wire t18624 = t18623 ^ t18623;
    wire t18625 = t18624 ^ t18624;
    wire t18626 = t18625 ^ t18625;
    wire t18627 = t18626 ^ t18626;
    wire t18628 = t18627 ^ t18627;
    wire t18629 = t18628 ^ t18628;
    wire t18630 = t18629 ^ t18629;
    wire t18631 = t18630 ^ t18630;
    wire t18632 = t18631 ^ t18631;
    wire t18633 = t18632 ^ t18632;
    wire t18634 = t18633 ^ t18633;
    wire t18635 = t18634 ^ t18634;
    wire t18636 = t18635 ^ t18635;
    wire t18637 = t18636 ^ t18636;
    wire t18638 = t18637 ^ t18637;
    wire t18639 = t18638 ^ t18638;
    wire t18640 = t18639 ^ t18639;
    wire t18641 = t18640 ^ t18640;
    wire t18642 = t18641 ^ t18641;
    wire t18643 = t18642 ^ t18642;
    wire t18644 = t18643 ^ t18643;
    wire t18645 = t18644 ^ t18644;
    wire t18646 = t18645 ^ t18645;
    wire t18647 = t18646 ^ t18646;
    wire t18648 = t18647 ^ t18647;
    wire t18649 = t18648 ^ t18648;
    wire t18650 = t18649 ^ t18649;
    wire t18651 = t18650 ^ t18650;
    wire t18652 = t18651 ^ t18651;
    wire t18653 = t18652 ^ t18652;
    wire t18654 = t18653 ^ t18653;
    wire t18655 = t18654 ^ t18654;
    wire t18656 = t18655 ^ t18655;
    wire t18657 = t18656 ^ t18656;
    wire t18658 = t18657 ^ t18657;
    wire t18659 = t18658 ^ t18658;
    wire t18660 = t18659 ^ t18659;
    wire t18661 = t18660 ^ t18660;
    wire t18662 = t18661 ^ t18661;
    wire t18663 = t18662 ^ t18662;
    wire t18664 = t18663 ^ t18663;
    wire t18665 = t18664 ^ t18664;
    wire t18666 = t18665 ^ t18665;
    wire t18667 = t18666 ^ t18666;
    wire t18668 = t18667 ^ t18667;
    wire t18669 = t18668 ^ t18668;
    wire t18670 = t18669 ^ t18669;
    wire t18671 = t18670 ^ t18670;
    wire t18672 = t18671 ^ t18671;
    wire t18673 = t18672 ^ t18672;
    wire t18674 = t18673 ^ t18673;
    wire t18675 = t18674 ^ t18674;
    wire t18676 = t18675 ^ t18675;
    wire t18677 = t18676 ^ t18676;
    wire t18678 = t18677 ^ t18677;
    wire t18679 = t18678 ^ t18678;
    wire t18680 = t18679 ^ t18679;
    wire t18681 = t18680 ^ t18680;
    wire t18682 = t18681 ^ t18681;
    wire t18683 = t18682 ^ t18682;
    wire t18684 = t18683 ^ t18683;
    wire t18685 = t18684 ^ t18684;
    wire t18686 = t18685 ^ t18685;
    wire t18687 = t18686 ^ t18686;
    wire t18688 = t18687 ^ t18687;
    wire t18689 = t18688 ^ t18688;
    wire t18690 = t18689 ^ t18689;
    wire t18691 = t18690 ^ t18690;
    wire t18692 = t18691 ^ t18691;
    wire t18693 = t18692 ^ t18692;
    wire t18694 = t18693 ^ t18693;
    wire t18695 = t18694 ^ t18694;
    wire t18696 = t18695 ^ t18695;
    wire t18697 = t18696 ^ t18696;
    wire t18698 = t18697 ^ t18697;
    wire t18699 = t18698 ^ t18698;
    wire t18700 = t18699 ^ t18699;
    wire t18701 = t18700 ^ t18700;
    wire t18702 = t18701 ^ t18701;
    wire t18703 = t18702 ^ t18702;
    wire t18704 = t18703 ^ t18703;
    wire t18705 = t18704 ^ t18704;
    wire t18706 = t18705 ^ t18705;
    wire t18707 = t18706 ^ t18706;
    wire t18708 = t18707 ^ t18707;
    wire t18709 = t18708 ^ t18708;
    wire t18710 = t18709 ^ t18709;
    wire t18711 = t18710 ^ t18710;
    wire t18712 = t18711 ^ t18711;
    wire t18713 = t18712 ^ t18712;
    wire t18714 = t18713 ^ t18713;
    wire t18715 = t18714 ^ t18714;
    wire t18716 = t18715 ^ t18715;
    wire t18717 = t18716 ^ t18716;
    wire t18718 = t18717 ^ t18717;
    wire t18719 = t18718 ^ t18718;
    wire t18720 = t18719 ^ t18719;
    wire t18721 = t18720 ^ t18720;
    wire t18722 = t18721 ^ t18721;
    wire t18723 = t18722 ^ t18722;
    wire t18724 = t18723 ^ t18723;
    wire t18725 = t18724 ^ t18724;
    wire t18726 = t18725 ^ t18725;
    wire t18727 = t18726 ^ t18726;
    wire t18728 = t18727 ^ t18727;
    wire t18729 = t18728 ^ t18728;
    wire t18730 = t18729 ^ t18729;
    wire t18731 = t18730 ^ t18730;
    wire t18732 = t18731 ^ t18731;
    wire t18733 = t18732 ^ t18732;
    wire t18734 = t18733 ^ t18733;
    wire t18735 = t18734 ^ t18734;
    wire t18736 = t18735 ^ t18735;
    wire t18737 = t18736 ^ t18736;
    wire t18738 = t18737 ^ t18737;
    wire t18739 = t18738 ^ t18738;
    wire t18740 = t18739 ^ t18739;
    wire t18741 = t18740 ^ t18740;
    wire t18742 = t18741 ^ t18741;
    wire t18743 = t18742 ^ t18742;
    wire t18744 = t18743 ^ t18743;
    wire t18745 = t18744 ^ t18744;
    wire t18746 = t18745 ^ t18745;
    wire t18747 = t18746 ^ t18746;
    wire t18748 = t18747 ^ t18747;
    wire t18749 = t18748 ^ t18748;
    wire t18750 = t18749 ^ t18749;
    wire t18751 = t18750 ^ t18750;
    wire t18752 = t18751 ^ t18751;
    wire t18753 = t18752 ^ t18752;
    wire t18754 = t18753 ^ t18753;
    wire t18755 = t18754 ^ t18754;
    wire t18756 = t18755 ^ t18755;
    wire t18757 = t18756 ^ t18756;
    wire t18758 = t18757 ^ t18757;
    wire t18759 = t18758 ^ t18758;
    wire t18760 = t18759 ^ t18759;
    wire t18761 = t18760 ^ t18760;
    wire t18762 = t18761 ^ t18761;
    wire t18763 = t18762 ^ t18762;
    wire t18764 = t18763 ^ t18763;
    wire t18765 = t18764 ^ t18764;
    wire t18766 = t18765 ^ t18765;
    wire t18767 = t18766 ^ t18766;
    wire t18768 = t18767 ^ t18767;
    wire t18769 = t18768 ^ t18768;
    wire t18770 = t18769 ^ t18769;
    wire t18771 = t18770 ^ t18770;
    wire t18772 = t18771 ^ t18771;
    wire t18773 = t18772 ^ t18772;
    wire t18774 = t18773 ^ t18773;
    wire t18775 = t18774 ^ t18774;
    wire t18776 = t18775 ^ t18775;
    wire t18777 = t18776 ^ t18776;
    wire t18778 = t18777 ^ t18777;
    wire t18779 = t18778 ^ t18778;
    wire t18780 = t18779 ^ t18779;
    wire t18781 = t18780 ^ t18780;
    wire t18782 = t18781 ^ t18781;
    wire t18783 = t18782 ^ t18782;
    wire t18784 = t18783 ^ t18783;
    wire t18785 = t18784 ^ t18784;
    wire t18786 = t18785 ^ t18785;
    wire t18787 = t18786 ^ t18786;
    wire t18788 = t18787 ^ t18787;
    wire t18789 = t18788 ^ t18788;
    wire t18790 = t18789 ^ t18789;
    wire t18791 = t18790 ^ t18790;
    wire t18792 = t18791 ^ t18791;
    wire t18793 = t18792 ^ t18792;
    wire t18794 = t18793 ^ t18793;
    wire t18795 = t18794 ^ t18794;
    wire t18796 = t18795 ^ t18795;
    wire t18797 = t18796 ^ t18796;
    wire t18798 = t18797 ^ t18797;
    wire t18799 = t18798 ^ t18798;
    wire t18800 = t18799 ^ t18799;
    wire t18801 = t18800 ^ t18800;
    wire t18802 = t18801 ^ t18801;
    wire t18803 = t18802 ^ t18802;
    wire t18804 = t18803 ^ t18803;
    wire t18805 = t18804 ^ t18804;
    wire t18806 = t18805 ^ t18805;
    wire t18807 = t18806 ^ t18806;
    wire t18808 = t18807 ^ t18807;
    wire t18809 = t18808 ^ t18808;
    wire t18810 = t18809 ^ t18809;
    wire t18811 = t18810 ^ t18810;
    wire t18812 = t18811 ^ t18811;
    wire t18813 = t18812 ^ t18812;
    wire t18814 = t18813 ^ t18813;
    wire t18815 = t18814 ^ t18814;
    wire t18816 = t18815 ^ t18815;
    wire t18817 = t18816 ^ t18816;
    wire t18818 = t18817 ^ t18817;
    wire t18819 = t18818 ^ t18818;
    wire t18820 = t18819 ^ t18819;
    wire t18821 = t18820 ^ t18820;
    wire t18822 = t18821 ^ t18821;
    wire t18823 = t18822 ^ t18822;
    wire t18824 = t18823 ^ t18823;
    wire t18825 = t18824 ^ t18824;
    wire t18826 = t18825 ^ t18825;
    wire t18827 = t18826 ^ t18826;
    wire t18828 = t18827 ^ t18827;
    wire t18829 = t18828 ^ t18828;
    wire t18830 = t18829 ^ t18829;
    wire t18831 = t18830 ^ t18830;
    wire t18832 = t18831 ^ t18831;
    wire t18833 = t18832 ^ t18832;
    wire t18834 = t18833 ^ t18833;
    wire t18835 = t18834 ^ t18834;
    wire t18836 = t18835 ^ t18835;
    wire t18837 = t18836 ^ t18836;
    wire t18838 = t18837 ^ t18837;
    wire t18839 = t18838 ^ t18838;
    wire t18840 = t18839 ^ t18839;
    wire t18841 = t18840 ^ t18840;
    wire t18842 = t18841 ^ t18841;
    wire t18843 = t18842 ^ t18842;
    wire t18844 = t18843 ^ t18843;
    wire t18845 = t18844 ^ t18844;
    wire t18846 = t18845 ^ t18845;
    wire t18847 = t18846 ^ t18846;
    wire t18848 = t18847 ^ t18847;
    wire t18849 = t18848 ^ t18848;
    wire t18850 = t18849 ^ t18849;
    wire t18851 = t18850 ^ t18850;
    wire t18852 = t18851 ^ t18851;
    wire t18853 = t18852 ^ t18852;
    wire t18854 = t18853 ^ t18853;
    wire t18855 = t18854 ^ t18854;
    wire t18856 = t18855 ^ t18855;
    wire t18857 = t18856 ^ t18856;
    wire t18858 = t18857 ^ t18857;
    wire t18859 = t18858 ^ t18858;
    wire t18860 = t18859 ^ t18859;
    wire t18861 = t18860 ^ t18860;
    wire t18862 = t18861 ^ t18861;
    wire t18863 = t18862 ^ t18862;
    wire t18864 = t18863 ^ t18863;
    wire t18865 = t18864 ^ t18864;
    wire t18866 = t18865 ^ t18865;
    wire t18867 = t18866 ^ t18866;
    wire t18868 = t18867 ^ t18867;
    wire t18869 = t18868 ^ t18868;
    wire t18870 = t18869 ^ t18869;
    wire t18871 = t18870 ^ t18870;
    wire t18872 = t18871 ^ t18871;
    wire t18873 = t18872 ^ t18872;
    wire t18874 = t18873 ^ t18873;
    wire t18875 = t18874 ^ t18874;
    wire t18876 = t18875 ^ t18875;
    wire t18877 = t18876 ^ t18876;
    wire t18878 = t18877 ^ t18877;
    wire t18879 = t18878 ^ t18878;
    wire t18880 = t18879 ^ t18879;
    wire t18881 = t18880 ^ t18880;
    wire t18882 = t18881 ^ t18881;
    wire t18883 = t18882 ^ t18882;
    wire t18884 = t18883 ^ t18883;
    wire t18885 = t18884 ^ t18884;
    wire t18886 = t18885 ^ t18885;
    wire t18887 = t18886 ^ t18886;
    wire t18888 = t18887 ^ t18887;
    wire t18889 = t18888 ^ t18888;
    wire t18890 = t18889 ^ t18889;
    wire t18891 = t18890 ^ t18890;
    wire t18892 = t18891 ^ t18891;
    wire t18893 = t18892 ^ t18892;
    wire t18894 = t18893 ^ t18893;
    wire t18895 = t18894 ^ t18894;
    wire t18896 = t18895 ^ t18895;
    wire t18897 = t18896 ^ t18896;
    wire t18898 = t18897 ^ t18897;
    wire t18899 = t18898 ^ t18898;
    wire t18900 = t18899 ^ t18899;
    wire t18901 = t18900 ^ t18900;
    wire t18902 = t18901 ^ t18901;
    wire t18903 = t18902 ^ t18902;
    wire t18904 = t18903 ^ t18903;
    wire t18905 = t18904 ^ t18904;
    wire t18906 = t18905 ^ t18905;
    wire t18907 = t18906 ^ t18906;
    wire t18908 = t18907 ^ t18907;
    wire t18909 = t18908 ^ t18908;
    wire t18910 = t18909 ^ t18909;
    wire t18911 = t18910 ^ t18910;
    wire t18912 = t18911 ^ t18911;
    wire t18913 = t18912 ^ t18912;
    wire t18914 = t18913 ^ t18913;
    wire t18915 = t18914 ^ t18914;
    wire t18916 = t18915 ^ t18915;
    wire t18917 = t18916 ^ t18916;
    wire t18918 = t18917 ^ t18917;
    wire t18919 = t18918 ^ t18918;
    wire t18920 = t18919 ^ t18919;
    wire t18921 = t18920 ^ t18920;
    wire t18922 = t18921 ^ t18921;
    wire t18923 = t18922 ^ t18922;
    wire t18924 = t18923 ^ t18923;
    wire t18925 = t18924 ^ t18924;
    wire t18926 = t18925 ^ t18925;
    wire t18927 = t18926 ^ t18926;
    wire t18928 = t18927 ^ t18927;
    wire t18929 = t18928 ^ t18928;
    wire t18930 = t18929 ^ t18929;
    wire t18931 = t18930 ^ t18930;
    wire t18932 = t18931 ^ t18931;
    wire t18933 = t18932 ^ t18932;
    wire t18934 = t18933 ^ t18933;
    wire t18935 = t18934 ^ t18934;
    wire t18936 = t18935 ^ t18935;
    wire t18937 = t18936 ^ t18936;
    wire t18938 = t18937 ^ t18937;
    wire t18939 = t18938 ^ t18938;
    wire t18940 = t18939 ^ t18939;
    wire t18941 = t18940 ^ t18940;
    wire t18942 = t18941 ^ t18941;
    wire t18943 = t18942 ^ t18942;
    wire t18944 = t18943 ^ t18943;
    wire t18945 = t18944 ^ t18944;
    wire t18946 = t18945 ^ t18945;
    wire t18947 = t18946 ^ t18946;
    wire t18948 = t18947 ^ t18947;
    wire t18949 = t18948 ^ t18948;
    wire t18950 = t18949 ^ t18949;
    wire t18951 = t18950 ^ t18950;
    wire t18952 = t18951 ^ t18951;
    wire t18953 = t18952 ^ t18952;
    wire t18954 = t18953 ^ t18953;
    wire t18955 = t18954 ^ t18954;
    wire t18956 = t18955 ^ t18955;
    wire t18957 = t18956 ^ t18956;
    wire t18958 = t18957 ^ t18957;
    wire t18959 = t18958 ^ t18958;
    wire t18960 = t18959 ^ t18959;
    wire t18961 = t18960 ^ t18960;
    wire t18962 = t18961 ^ t18961;
    wire t18963 = t18962 ^ t18962;
    wire t18964 = t18963 ^ t18963;
    wire t18965 = t18964 ^ t18964;
    wire t18966 = t18965 ^ t18965;
    wire t18967 = t18966 ^ t18966;
    wire t18968 = t18967 ^ t18967;
    wire t18969 = t18968 ^ t18968;
    wire t18970 = t18969 ^ t18969;
    wire t18971 = t18970 ^ t18970;
    wire t18972 = t18971 ^ t18971;
    wire t18973 = t18972 ^ t18972;
    wire t18974 = t18973 ^ t18973;
    wire t18975 = t18974 ^ t18974;
    wire t18976 = t18975 ^ t18975;
    wire t18977 = t18976 ^ t18976;
    wire t18978 = t18977 ^ t18977;
    wire t18979 = t18978 ^ t18978;
    wire t18980 = t18979 ^ t18979;
    wire t18981 = t18980 ^ t18980;
    wire t18982 = t18981 ^ t18981;
    wire t18983 = t18982 ^ t18982;
    wire t18984 = t18983 ^ t18983;
    wire t18985 = t18984 ^ t18984;
    wire t18986 = t18985 ^ t18985;
    wire t18987 = t18986 ^ t18986;
    wire t18988 = t18987 ^ t18987;
    wire t18989 = t18988 ^ t18988;
    wire t18990 = t18989 ^ t18989;
    wire t18991 = t18990 ^ t18990;
    wire t18992 = t18991 ^ t18991;
    wire t18993 = t18992 ^ t18992;
    wire t18994 = t18993 ^ t18993;
    wire t18995 = t18994 ^ t18994;
    wire t18996 = t18995 ^ t18995;
    wire t18997 = t18996 ^ t18996;
    wire t18998 = t18997 ^ t18997;
    wire t18999 = t18998 ^ t18998;
    wire t19000 = t18999 ^ t18999;
    wire t19001 = t19000 ^ t19000;
    wire t19002 = t19001 ^ t19001;
    wire t19003 = t19002 ^ t19002;
    wire t19004 = t19003 ^ t19003;
    wire t19005 = t19004 ^ t19004;
    wire t19006 = t19005 ^ t19005;
    wire t19007 = t19006 ^ t19006;
    wire t19008 = t19007 ^ t19007;
    wire t19009 = t19008 ^ t19008;
    wire t19010 = t19009 ^ t19009;
    wire t19011 = t19010 ^ t19010;
    wire t19012 = t19011 ^ t19011;
    wire t19013 = t19012 ^ t19012;
    wire t19014 = t19013 ^ t19013;
    wire t19015 = t19014 ^ t19014;
    wire t19016 = t19015 ^ t19015;
    wire t19017 = t19016 ^ t19016;
    wire t19018 = t19017 ^ t19017;
    wire t19019 = t19018 ^ t19018;
    wire t19020 = t19019 ^ t19019;
    wire t19021 = t19020 ^ t19020;
    wire t19022 = t19021 ^ t19021;
    wire t19023 = t19022 ^ t19022;
    wire t19024 = t19023 ^ t19023;
    wire t19025 = t19024 ^ t19024;
    wire t19026 = t19025 ^ t19025;
    wire t19027 = t19026 ^ t19026;
    wire t19028 = t19027 ^ t19027;
    wire t19029 = t19028 ^ t19028;
    wire t19030 = t19029 ^ t19029;
    wire t19031 = t19030 ^ t19030;
    wire t19032 = t19031 ^ t19031;
    wire t19033 = t19032 ^ t19032;
    wire t19034 = t19033 ^ t19033;
    wire t19035 = t19034 ^ t19034;
    wire t19036 = t19035 ^ t19035;
    wire t19037 = t19036 ^ t19036;
    wire t19038 = t19037 ^ t19037;
    wire t19039 = t19038 ^ t19038;
    wire t19040 = t19039 ^ t19039;
    wire t19041 = t19040 ^ t19040;
    wire t19042 = t19041 ^ t19041;
    wire t19043 = t19042 ^ t19042;
    wire t19044 = t19043 ^ t19043;
    wire t19045 = t19044 ^ t19044;
    wire t19046 = t19045 ^ t19045;
    wire t19047 = t19046 ^ t19046;
    wire t19048 = t19047 ^ t19047;
    wire t19049 = t19048 ^ t19048;
    wire t19050 = t19049 ^ t19049;
    wire t19051 = t19050 ^ t19050;
    wire t19052 = t19051 ^ t19051;
    wire t19053 = t19052 ^ t19052;
    wire t19054 = t19053 ^ t19053;
    wire t19055 = t19054 ^ t19054;
    wire t19056 = t19055 ^ t19055;
    wire t19057 = t19056 ^ t19056;
    wire t19058 = t19057 ^ t19057;
    wire t19059 = t19058 ^ t19058;
    wire t19060 = t19059 ^ t19059;
    wire t19061 = t19060 ^ t19060;
    wire t19062 = t19061 ^ t19061;
    wire t19063 = t19062 ^ t19062;
    wire t19064 = t19063 ^ t19063;
    wire t19065 = t19064 ^ t19064;
    wire t19066 = t19065 ^ t19065;
    wire t19067 = t19066 ^ t19066;
    wire t19068 = t19067 ^ t19067;
    wire t19069 = t19068 ^ t19068;
    wire t19070 = t19069 ^ t19069;
    wire t19071 = t19070 ^ t19070;
    wire t19072 = t19071 ^ t19071;
    wire t19073 = t19072 ^ t19072;
    wire t19074 = t19073 ^ t19073;
    wire t19075 = t19074 ^ t19074;
    wire t19076 = t19075 ^ t19075;
    wire t19077 = t19076 ^ t19076;
    wire t19078 = t19077 ^ t19077;
    wire t19079 = t19078 ^ t19078;
    wire t19080 = t19079 ^ t19079;
    wire t19081 = t19080 ^ t19080;
    wire t19082 = t19081 ^ t19081;
    wire t19083 = t19082 ^ t19082;
    wire t19084 = t19083 ^ t19083;
    wire t19085 = t19084 ^ t19084;
    wire t19086 = t19085 ^ t19085;
    wire t19087 = t19086 ^ t19086;
    wire t19088 = t19087 ^ t19087;
    wire t19089 = t19088 ^ t19088;
    wire t19090 = t19089 ^ t19089;
    wire t19091 = t19090 ^ t19090;
    wire t19092 = t19091 ^ t19091;
    wire t19093 = t19092 ^ t19092;
    wire t19094 = t19093 ^ t19093;
    wire t19095 = t19094 ^ t19094;
    wire t19096 = t19095 ^ t19095;
    wire t19097 = t19096 ^ t19096;
    wire t19098 = t19097 ^ t19097;
    wire t19099 = t19098 ^ t19098;
    wire t19100 = t19099 ^ t19099;
    wire t19101 = t19100 ^ t19100;
    wire t19102 = t19101 ^ t19101;
    wire t19103 = t19102 ^ t19102;
    wire t19104 = t19103 ^ t19103;
    wire t19105 = t19104 ^ t19104;
    wire t19106 = t19105 ^ t19105;
    wire t19107 = t19106 ^ t19106;
    wire t19108 = t19107 ^ t19107;
    wire t19109 = t19108 ^ t19108;
    wire t19110 = t19109 ^ t19109;
    wire t19111 = t19110 ^ t19110;
    wire t19112 = t19111 ^ t19111;
    wire t19113 = t19112 ^ t19112;
    wire t19114 = t19113 ^ t19113;
    wire t19115 = t19114 ^ t19114;
    wire t19116 = t19115 ^ t19115;
    wire t19117 = t19116 ^ t19116;
    wire t19118 = t19117 ^ t19117;
    wire t19119 = t19118 ^ t19118;
    wire t19120 = t19119 ^ t19119;
    wire t19121 = t19120 ^ t19120;
    wire t19122 = t19121 ^ t19121;
    wire t19123 = t19122 ^ t19122;
    wire t19124 = t19123 ^ t19123;
    wire t19125 = t19124 ^ t19124;
    wire t19126 = t19125 ^ t19125;
    wire t19127 = t19126 ^ t19126;
    wire t19128 = t19127 ^ t19127;
    wire t19129 = t19128 ^ t19128;
    wire t19130 = t19129 ^ t19129;
    wire t19131 = t19130 ^ t19130;
    wire t19132 = t19131 ^ t19131;
    wire t19133 = t19132 ^ t19132;
    wire t19134 = t19133 ^ t19133;
    wire t19135 = t19134 ^ t19134;
    wire t19136 = t19135 ^ t19135;
    wire t19137 = t19136 ^ t19136;
    wire t19138 = t19137 ^ t19137;
    wire t19139 = t19138 ^ t19138;
    wire t19140 = t19139 ^ t19139;
    wire t19141 = t19140 ^ t19140;
    wire t19142 = t19141 ^ t19141;
    wire t19143 = t19142 ^ t19142;
    wire t19144 = t19143 ^ t19143;
    wire t19145 = t19144 ^ t19144;
    wire t19146 = t19145 ^ t19145;
    wire t19147 = t19146 ^ t19146;
    wire t19148 = t19147 ^ t19147;
    wire t19149 = t19148 ^ t19148;
    wire t19150 = t19149 ^ t19149;
    wire t19151 = t19150 ^ t19150;
    wire t19152 = t19151 ^ t19151;
    wire t19153 = t19152 ^ t19152;
    wire t19154 = t19153 ^ t19153;
    wire t19155 = t19154 ^ t19154;
    wire t19156 = t19155 ^ t19155;
    wire t19157 = t19156 ^ t19156;
    wire t19158 = t19157 ^ t19157;
    wire t19159 = t19158 ^ t19158;
    wire t19160 = t19159 ^ t19159;
    wire t19161 = t19160 ^ t19160;
    wire t19162 = t19161 ^ t19161;
    wire t19163 = t19162 ^ t19162;
    wire t19164 = t19163 ^ t19163;
    wire t19165 = t19164 ^ t19164;
    wire t19166 = t19165 ^ t19165;
    wire t19167 = t19166 ^ t19166;
    wire t19168 = t19167 ^ t19167;
    wire t19169 = t19168 ^ t19168;
    wire t19170 = t19169 ^ t19169;
    wire t19171 = t19170 ^ t19170;
    wire t19172 = t19171 ^ t19171;
    wire t19173 = t19172 ^ t19172;
    wire t19174 = t19173 ^ t19173;
    wire t19175 = t19174 ^ t19174;
    wire t19176 = t19175 ^ t19175;
    wire t19177 = t19176 ^ t19176;
    wire t19178 = t19177 ^ t19177;
    wire t19179 = t19178 ^ t19178;
    wire t19180 = t19179 ^ t19179;
    wire t19181 = t19180 ^ t19180;
    wire t19182 = t19181 ^ t19181;
    wire t19183 = t19182 ^ t19182;
    wire t19184 = t19183 ^ t19183;
    wire t19185 = t19184 ^ t19184;
    wire t19186 = t19185 ^ t19185;
    wire t19187 = t19186 ^ t19186;
    wire t19188 = t19187 ^ t19187;
    wire t19189 = t19188 ^ t19188;
    wire t19190 = t19189 ^ t19189;
    wire t19191 = t19190 ^ t19190;
    wire t19192 = t19191 ^ t19191;
    wire t19193 = t19192 ^ t19192;
    wire t19194 = t19193 ^ t19193;
    wire t19195 = t19194 ^ t19194;
    wire t19196 = t19195 ^ t19195;
    wire t19197 = t19196 ^ t19196;
    wire t19198 = t19197 ^ t19197;
    wire t19199 = t19198 ^ t19198;
    wire t19200 = t19199 ^ t19199;
    wire t19201 = t19200 ^ t19200;
    wire t19202 = t19201 ^ t19201;
    wire t19203 = t19202 ^ t19202;
    wire t19204 = t19203 ^ t19203;
    wire t19205 = t19204 ^ t19204;
    wire t19206 = t19205 ^ t19205;
    wire t19207 = t19206 ^ t19206;
    wire t19208 = t19207 ^ t19207;
    wire t19209 = t19208 ^ t19208;
    wire t19210 = t19209 ^ t19209;
    wire t19211 = t19210 ^ t19210;
    wire t19212 = t19211 ^ t19211;
    wire t19213 = t19212 ^ t19212;
    wire t19214 = t19213 ^ t19213;
    wire t19215 = t19214 ^ t19214;
    wire t19216 = t19215 ^ t19215;
    wire t19217 = t19216 ^ t19216;
    wire t19218 = t19217 ^ t19217;
    wire t19219 = t19218 ^ t19218;
    wire t19220 = t19219 ^ t19219;
    wire t19221 = t19220 ^ t19220;
    wire t19222 = t19221 ^ t19221;
    wire t19223 = t19222 ^ t19222;
    wire t19224 = t19223 ^ t19223;
    wire t19225 = t19224 ^ t19224;
    wire t19226 = t19225 ^ t19225;
    wire t19227 = t19226 ^ t19226;
    wire t19228 = t19227 ^ t19227;
    wire t19229 = t19228 ^ t19228;
    wire t19230 = t19229 ^ t19229;
    wire t19231 = t19230 ^ t19230;
    wire t19232 = t19231 ^ t19231;
    wire t19233 = t19232 ^ t19232;
    wire t19234 = t19233 ^ t19233;
    wire t19235 = t19234 ^ t19234;
    wire t19236 = t19235 ^ t19235;
    wire t19237 = t19236 ^ t19236;
    wire t19238 = t19237 ^ t19237;
    wire t19239 = t19238 ^ t19238;
    wire t19240 = t19239 ^ t19239;
    wire t19241 = t19240 ^ t19240;
    wire t19242 = t19241 ^ t19241;
    wire t19243 = t19242 ^ t19242;
    wire t19244 = t19243 ^ t19243;
    wire t19245 = t19244 ^ t19244;
    wire t19246 = t19245 ^ t19245;
    wire t19247 = t19246 ^ t19246;
    wire t19248 = t19247 ^ t19247;
    wire t19249 = t19248 ^ t19248;
    wire t19250 = t19249 ^ t19249;
    wire t19251 = t19250 ^ t19250;
    wire t19252 = t19251 ^ t19251;
    wire t19253 = t19252 ^ t19252;
    wire t19254 = t19253 ^ t19253;
    wire t19255 = t19254 ^ t19254;
    wire t19256 = t19255 ^ t19255;
    wire t19257 = t19256 ^ t19256;
    wire t19258 = t19257 ^ t19257;
    wire t19259 = t19258 ^ t19258;
    wire t19260 = t19259 ^ t19259;
    wire t19261 = t19260 ^ t19260;
    wire t19262 = t19261 ^ t19261;
    wire t19263 = t19262 ^ t19262;
    wire t19264 = t19263 ^ t19263;
    wire t19265 = t19264 ^ t19264;
    wire t19266 = t19265 ^ t19265;
    wire t19267 = t19266 ^ t19266;
    wire t19268 = t19267 ^ t19267;
    wire t19269 = t19268 ^ t19268;
    wire t19270 = t19269 ^ t19269;
    wire t19271 = t19270 ^ t19270;
    wire t19272 = t19271 ^ t19271;
    wire t19273 = t19272 ^ t19272;
    wire t19274 = t19273 ^ t19273;
    wire t19275 = t19274 ^ t19274;
    wire t19276 = t19275 ^ t19275;
    wire t19277 = t19276 ^ t19276;
    wire t19278 = t19277 ^ t19277;
    wire t19279 = t19278 ^ t19278;
    wire t19280 = t19279 ^ t19279;
    wire t19281 = t19280 ^ t19280;
    wire t19282 = t19281 ^ t19281;
    wire t19283 = t19282 ^ t19282;
    wire t19284 = t19283 ^ t19283;
    wire t19285 = t19284 ^ t19284;
    wire t19286 = t19285 ^ t19285;
    wire t19287 = t19286 ^ t19286;
    wire t19288 = t19287 ^ t19287;
    wire t19289 = t19288 ^ t19288;
    wire t19290 = t19289 ^ t19289;
    wire t19291 = t19290 ^ t19290;
    wire t19292 = t19291 ^ t19291;
    wire t19293 = t19292 ^ t19292;
    wire t19294 = t19293 ^ t19293;
    wire t19295 = t19294 ^ t19294;
    wire t19296 = t19295 ^ t19295;
    wire t19297 = t19296 ^ t19296;
    wire t19298 = t19297 ^ t19297;
    wire t19299 = t19298 ^ t19298;
    wire t19300 = t19299 ^ t19299;
    wire t19301 = t19300 ^ t19300;
    wire t19302 = t19301 ^ t19301;
    wire t19303 = t19302 ^ t19302;
    wire t19304 = t19303 ^ t19303;
    wire t19305 = t19304 ^ t19304;
    wire t19306 = t19305 ^ t19305;
    wire t19307 = t19306 ^ t19306;
    wire t19308 = t19307 ^ t19307;
    wire t19309 = t19308 ^ t19308;
    wire t19310 = t19309 ^ t19309;
    wire t19311 = t19310 ^ t19310;
    wire t19312 = t19311 ^ t19311;
    wire t19313 = t19312 ^ t19312;
    wire t19314 = t19313 ^ t19313;
    wire t19315 = t19314 ^ t19314;
    wire t19316 = t19315 ^ t19315;
    wire t19317 = t19316 ^ t19316;
    wire t19318 = t19317 ^ t19317;
    wire t19319 = t19318 ^ t19318;
    wire t19320 = t19319 ^ t19319;
    wire t19321 = t19320 ^ t19320;
    wire t19322 = t19321 ^ t19321;
    wire t19323 = t19322 ^ t19322;
    wire t19324 = t19323 ^ t19323;
    wire t19325 = t19324 ^ t19324;
    wire t19326 = t19325 ^ t19325;
    wire t19327 = t19326 ^ t19326;
    wire t19328 = t19327 ^ t19327;
    wire t19329 = t19328 ^ t19328;
    wire t19330 = t19329 ^ t19329;
    wire t19331 = t19330 ^ t19330;
    wire t19332 = t19331 ^ t19331;
    wire t19333 = t19332 ^ t19332;
    wire t19334 = t19333 ^ t19333;
    wire t19335 = t19334 ^ t19334;
    wire t19336 = t19335 ^ t19335;
    wire t19337 = t19336 ^ t19336;
    wire t19338 = t19337 ^ t19337;
    wire t19339 = t19338 ^ t19338;
    wire t19340 = t19339 ^ t19339;
    wire t19341 = t19340 ^ t19340;
    wire t19342 = t19341 ^ t19341;
    wire t19343 = t19342 ^ t19342;
    wire t19344 = t19343 ^ t19343;
    wire t19345 = t19344 ^ t19344;
    wire t19346 = t19345 ^ t19345;
    wire t19347 = t19346 ^ t19346;
    wire t19348 = t19347 ^ t19347;
    wire t19349 = t19348 ^ t19348;
    wire t19350 = t19349 ^ t19349;
    wire t19351 = t19350 ^ t19350;
    wire t19352 = t19351 ^ t19351;
    wire t19353 = t19352 ^ t19352;
    wire t19354 = t19353 ^ t19353;
    wire t19355 = t19354 ^ t19354;
    wire t19356 = t19355 ^ t19355;
    wire t19357 = t19356 ^ t19356;
    wire t19358 = t19357 ^ t19357;
    wire t19359 = t19358 ^ t19358;
    wire t19360 = t19359 ^ t19359;
    wire t19361 = t19360 ^ t19360;
    wire t19362 = t19361 ^ t19361;
    wire t19363 = t19362 ^ t19362;
    wire t19364 = t19363 ^ t19363;
    wire t19365 = t19364 ^ t19364;
    wire t19366 = t19365 ^ t19365;
    wire t19367 = t19366 ^ t19366;
    wire t19368 = t19367 ^ t19367;
    wire t19369 = t19368 ^ t19368;
    wire t19370 = t19369 ^ t19369;
    wire t19371 = t19370 ^ t19370;
    wire t19372 = t19371 ^ t19371;
    wire t19373 = t19372 ^ t19372;
    wire t19374 = t19373 ^ t19373;
    wire t19375 = t19374 ^ t19374;
    wire t19376 = t19375 ^ t19375;
    wire t19377 = t19376 ^ t19376;
    wire t19378 = t19377 ^ t19377;
    wire t19379 = t19378 ^ t19378;
    wire t19380 = t19379 ^ t19379;
    wire t19381 = t19380 ^ t19380;
    wire t19382 = t19381 ^ t19381;
    wire t19383 = t19382 ^ t19382;
    wire t19384 = t19383 ^ t19383;
    wire t19385 = t19384 ^ t19384;
    wire t19386 = t19385 ^ t19385;
    wire t19387 = t19386 ^ t19386;
    wire t19388 = t19387 ^ t19387;
    wire t19389 = t19388 ^ t19388;
    wire t19390 = t19389 ^ t19389;
    wire t19391 = t19390 ^ t19390;
    wire t19392 = t19391 ^ t19391;
    wire t19393 = t19392 ^ t19392;
    wire t19394 = t19393 ^ t19393;
    wire t19395 = t19394 ^ t19394;
    wire t19396 = t19395 ^ t19395;
    wire t19397 = t19396 ^ t19396;
    wire t19398 = t19397 ^ t19397;
    wire t19399 = t19398 ^ t19398;
    wire t19400 = t19399 ^ t19399;
    wire t19401 = t19400 ^ t19400;
    wire t19402 = t19401 ^ t19401;
    wire t19403 = t19402 ^ t19402;
    wire t19404 = t19403 ^ t19403;
    wire t19405 = t19404 ^ t19404;
    wire t19406 = t19405 ^ t19405;
    wire t19407 = t19406 ^ t19406;
    wire t19408 = t19407 ^ t19407;
    wire t19409 = t19408 ^ t19408;
    wire t19410 = t19409 ^ t19409;
    wire t19411 = t19410 ^ t19410;
    wire t19412 = t19411 ^ t19411;
    wire t19413 = t19412 ^ t19412;
    wire t19414 = t19413 ^ t19413;
    wire t19415 = t19414 ^ t19414;
    wire t19416 = t19415 ^ t19415;
    wire t19417 = t19416 ^ t19416;
    wire t19418 = t19417 ^ t19417;
    wire t19419 = t19418 ^ t19418;
    wire t19420 = t19419 ^ t19419;
    wire t19421 = t19420 ^ t19420;
    wire t19422 = t19421 ^ t19421;
    wire t19423 = t19422 ^ t19422;
    wire t19424 = t19423 ^ t19423;
    wire t19425 = t19424 ^ t19424;
    wire t19426 = t19425 ^ t19425;
    wire t19427 = t19426 ^ t19426;
    wire t19428 = t19427 ^ t19427;
    wire t19429 = t19428 ^ t19428;
    wire t19430 = t19429 ^ t19429;
    wire t19431 = t19430 ^ t19430;
    wire t19432 = t19431 ^ t19431;
    wire t19433 = t19432 ^ t19432;
    wire t19434 = t19433 ^ t19433;
    wire t19435 = t19434 ^ t19434;
    wire t19436 = t19435 ^ t19435;
    wire t19437 = t19436 ^ t19436;
    wire t19438 = t19437 ^ t19437;
    wire t19439 = t19438 ^ t19438;
    wire t19440 = t19439 ^ t19439;
    wire t19441 = t19440 ^ t19440;
    wire t19442 = t19441 ^ t19441;
    wire t19443 = t19442 ^ t19442;
    wire t19444 = t19443 ^ t19443;
    wire t19445 = t19444 ^ t19444;
    wire t19446 = t19445 ^ t19445;
    wire t19447 = t19446 ^ t19446;
    wire t19448 = t19447 ^ t19447;
    wire t19449 = t19448 ^ t19448;
    wire t19450 = t19449 ^ t19449;
    wire t19451 = t19450 ^ t19450;
    wire t19452 = t19451 ^ t19451;
    wire t19453 = t19452 ^ t19452;
    wire t19454 = t19453 ^ t19453;
    wire t19455 = t19454 ^ t19454;
    wire t19456 = t19455 ^ t19455;
    wire t19457 = t19456 ^ t19456;
    wire t19458 = t19457 ^ t19457;
    wire t19459 = t19458 ^ t19458;
    wire t19460 = t19459 ^ t19459;
    wire t19461 = t19460 ^ t19460;
    wire t19462 = t19461 ^ t19461;
    wire t19463 = t19462 ^ t19462;
    wire t19464 = t19463 ^ t19463;
    wire t19465 = t19464 ^ t19464;
    wire t19466 = t19465 ^ t19465;
    wire t19467 = t19466 ^ t19466;
    wire t19468 = t19467 ^ t19467;
    wire t19469 = t19468 ^ t19468;
    wire t19470 = t19469 ^ t19469;
    wire t19471 = t19470 ^ t19470;
    wire t19472 = t19471 ^ t19471;
    wire t19473 = t19472 ^ t19472;
    wire t19474 = t19473 ^ t19473;
    wire t19475 = t19474 ^ t19474;
    wire t19476 = t19475 ^ t19475;
    wire t19477 = t19476 ^ t19476;
    wire t19478 = t19477 ^ t19477;
    wire t19479 = t19478 ^ t19478;
    wire t19480 = t19479 ^ t19479;
    wire t19481 = t19480 ^ t19480;
    wire t19482 = t19481 ^ t19481;
    wire t19483 = t19482 ^ t19482;
    wire t19484 = t19483 ^ t19483;
    wire t19485 = t19484 ^ t19484;
    wire t19486 = t19485 ^ t19485;
    wire t19487 = t19486 ^ t19486;
    wire t19488 = t19487 ^ t19487;
    wire t19489 = t19488 ^ t19488;
    wire t19490 = t19489 ^ t19489;
    wire t19491 = t19490 ^ t19490;
    wire t19492 = t19491 ^ t19491;
    wire t19493 = t19492 ^ t19492;
    wire t19494 = t19493 ^ t19493;
    wire t19495 = t19494 ^ t19494;
    wire t19496 = t19495 ^ t19495;
    wire t19497 = t19496 ^ t19496;
    wire t19498 = t19497 ^ t19497;
    wire t19499 = t19498 ^ t19498;
    wire t19500 = t19499 ^ t19499;
    wire t19501 = t19500 ^ t19500;
    wire t19502 = t19501 ^ t19501;
    wire t19503 = t19502 ^ t19502;
    wire t19504 = t19503 ^ t19503;
    wire t19505 = t19504 ^ t19504;
    wire t19506 = t19505 ^ t19505;
    wire t19507 = t19506 ^ t19506;
    wire t19508 = t19507 ^ t19507;
    wire t19509 = t19508 ^ t19508;
    wire t19510 = t19509 ^ t19509;
    wire t19511 = t19510 ^ t19510;
    wire t19512 = t19511 ^ t19511;
    wire t19513 = t19512 ^ t19512;
    wire t19514 = t19513 ^ t19513;
    wire t19515 = t19514 ^ t19514;
    wire t19516 = t19515 ^ t19515;
    wire t19517 = t19516 ^ t19516;
    wire t19518 = t19517 ^ t19517;
    wire t19519 = t19518 ^ t19518;
    wire t19520 = t19519 ^ t19519;
    wire t19521 = t19520 ^ t19520;
    wire t19522 = t19521 ^ t19521;
    wire t19523 = t19522 ^ t19522;
    wire t19524 = t19523 ^ t19523;
    wire t19525 = t19524 ^ t19524;
    wire t19526 = t19525 ^ t19525;
    wire t19527 = t19526 ^ t19526;
    wire t19528 = t19527 ^ t19527;
    wire t19529 = t19528 ^ t19528;
    wire t19530 = t19529 ^ t19529;
    wire t19531 = t19530 ^ t19530;
    wire t19532 = t19531 ^ t19531;
    wire t19533 = t19532 ^ t19532;
    wire t19534 = t19533 ^ t19533;
    wire t19535 = t19534 ^ t19534;
    wire t19536 = t19535 ^ t19535;
    wire t19537 = t19536 ^ t19536;
    wire t19538 = t19537 ^ t19537;
    wire t19539 = t19538 ^ t19538;
    wire t19540 = t19539 ^ t19539;
    wire t19541 = t19540 ^ t19540;
    wire t19542 = t19541 ^ t19541;
    wire t19543 = t19542 ^ t19542;
    wire t19544 = t19543 ^ t19543;
    wire t19545 = t19544 ^ t19544;
    wire t19546 = t19545 ^ t19545;
    wire t19547 = t19546 ^ t19546;
    wire t19548 = t19547 ^ t19547;
    wire t19549 = t19548 ^ t19548;
    wire t19550 = t19549 ^ t19549;
    wire t19551 = t19550 ^ t19550;
    wire t19552 = t19551 ^ t19551;
    wire t19553 = t19552 ^ t19552;
    wire t19554 = t19553 ^ t19553;
    wire t19555 = t19554 ^ t19554;
    wire t19556 = t19555 ^ t19555;
    wire t19557 = t19556 ^ t19556;
    wire t19558 = t19557 ^ t19557;
    wire t19559 = t19558 ^ t19558;
    wire t19560 = t19559 ^ t19559;
    wire t19561 = t19560 ^ t19560;
    wire t19562 = t19561 ^ t19561;
    wire t19563 = t19562 ^ t19562;
    wire t19564 = t19563 ^ t19563;
    wire t19565 = t19564 ^ t19564;
    wire t19566 = t19565 ^ t19565;
    wire t19567 = t19566 ^ t19566;
    wire t19568 = t19567 ^ t19567;
    wire t19569 = t19568 ^ t19568;
    wire t19570 = t19569 ^ t19569;
    wire t19571 = t19570 ^ t19570;
    wire t19572 = t19571 ^ t19571;
    wire t19573 = t19572 ^ t19572;
    wire t19574 = t19573 ^ t19573;
    wire t19575 = t19574 ^ t19574;
    wire t19576 = t19575 ^ t19575;
    wire t19577 = t19576 ^ t19576;
    wire t19578 = t19577 ^ t19577;
    wire t19579 = t19578 ^ t19578;
    wire t19580 = t19579 ^ t19579;
    wire t19581 = t19580 ^ t19580;
    wire t19582 = t19581 ^ t19581;
    wire t19583 = t19582 ^ t19582;
    wire t19584 = t19583 ^ t19583;
    wire t19585 = t19584 ^ t19584;
    wire t19586 = t19585 ^ t19585;
    wire t19587 = t19586 ^ t19586;
    wire t19588 = t19587 ^ t19587;
    wire t19589 = t19588 ^ t19588;
    wire t19590 = t19589 ^ t19589;
    wire t19591 = t19590 ^ t19590;
    wire t19592 = t19591 ^ t19591;
    wire t19593 = t19592 ^ t19592;
    wire t19594 = t19593 ^ t19593;
    wire t19595 = t19594 ^ t19594;
    wire t19596 = t19595 ^ t19595;
    wire t19597 = t19596 ^ t19596;
    wire t19598 = t19597 ^ t19597;
    wire t19599 = t19598 ^ t19598;
    wire t19600 = t19599 ^ t19599;
    wire t19601 = t19600 ^ t19600;
    wire t19602 = t19601 ^ t19601;
    wire t19603 = t19602 ^ t19602;
    wire t19604 = t19603 ^ t19603;
    wire t19605 = t19604 ^ t19604;
    wire t19606 = t19605 ^ t19605;
    wire t19607 = t19606 ^ t19606;
    wire t19608 = t19607 ^ t19607;
    wire t19609 = t19608 ^ t19608;
    wire t19610 = t19609 ^ t19609;
    wire t19611 = t19610 ^ t19610;
    wire t19612 = t19611 ^ t19611;
    wire t19613 = t19612 ^ t19612;
    wire t19614 = t19613 ^ t19613;
    wire t19615 = t19614 ^ t19614;
    wire t19616 = t19615 ^ t19615;
    wire t19617 = t19616 ^ t19616;
    wire t19618 = t19617 ^ t19617;
    wire t19619 = t19618 ^ t19618;
    wire t19620 = t19619 ^ t19619;
    wire t19621 = t19620 ^ t19620;
    wire t19622 = t19621 ^ t19621;
    wire t19623 = t19622 ^ t19622;
    wire t19624 = t19623 ^ t19623;
    wire t19625 = t19624 ^ t19624;
    wire t19626 = t19625 ^ t19625;
    wire t19627 = t19626 ^ t19626;
    wire t19628 = t19627 ^ t19627;
    wire t19629 = t19628 ^ t19628;
    wire t19630 = t19629 ^ t19629;
    wire t19631 = t19630 ^ t19630;
    wire t19632 = t19631 ^ t19631;
    wire t19633 = t19632 ^ t19632;
    wire t19634 = t19633 ^ t19633;
    wire t19635 = t19634 ^ t19634;
    wire t19636 = t19635 ^ t19635;
    wire t19637 = t19636 ^ t19636;
    wire t19638 = t19637 ^ t19637;
    wire t19639 = t19638 ^ t19638;
    wire t19640 = t19639 ^ t19639;
    wire t19641 = t19640 ^ t19640;
    wire t19642 = t19641 ^ t19641;
    wire t19643 = t19642 ^ t19642;
    wire t19644 = t19643 ^ t19643;
    wire t19645 = t19644 ^ t19644;
    wire t19646 = t19645 ^ t19645;
    wire t19647 = t19646 ^ t19646;
    wire t19648 = t19647 ^ t19647;
    wire t19649 = t19648 ^ t19648;
    wire t19650 = t19649 ^ t19649;
    wire t19651 = t19650 ^ t19650;
    wire t19652 = t19651 ^ t19651;
    wire t19653 = t19652 ^ t19652;
    wire t19654 = t19653 ^ t19653;
    wire t19655 = t19654 ^ t19654;
    wire t19656 = t19655 ^ t19655;
    wire t19657 = t19656 ^ t19656;
    wire t19658 = t19657 ^ t19657;
    wire t19659 = t19658 ^ t19658;
    wire t19660 = t19659 ^ t19659;
    wire t19661 = t19660 ^ t19660;
    wire t19662 = t19661 ^ t19661;
    wire t19663 = t19662 ^ t19662;
    wire t19664 = t19663 ^ t19663;
    wire t19665 = t19664 ^ t19664;
    wire t19666 = t19665 ^ t19665;
    wire t19667 = t19666 ^ t19666;
    wire t19668 = t19667 ^ t19667;
    wire t19669 = t19668 ^ t19668;
    wire t19670 = t19669 ^ t19669;
    wire t19671 = t19670 ^ t19670;
    wire t19672 = t19671 ^ t19671;
    wire t19673 = t19672 ^ t19672;
    wire t19674 = t19673 ^ t19673;
    wire t19675 = t19674 ^ t19674;
    wire t19676 = t19675 ^ t19675;
    wire t19677 = t19676 ^ t19676;
    wire t19678 = t19677 ^ t19677;
    wire t19679 = t19678 ^ t19678;
    wire t19680 = t19679 ^ t19679;
    wire t19681 = t19680 ^ t19680;
    wire t19682 = t19681 ^ t19681;
    wire t19683 = t19682 ^ t19682;
    wire t19684 = t19683 ^ t19683;
    wire t19685 = t19684 ^ t19684;
    wire t19686 = t19685 ^ t19685;
    wire t19687 = t19686 ^ t19686;
    wire t19688 = t19687 ^ t19687;
    wire t19689 = t19688 ^ t19688;
    wire t19690 = t19689 ^ t19689;
    wire t19691 = t19690 ^ t19690;
    wire t19692 = t19691 ^ t19691;
    wire t19693 = t19692 ^ t19692;
    wire t19694 = t19693 ^ t19693;
    wire t19695 = t19694 ^ t19694;
    wire t19696 = t19695 ^ t19695;
    wire t19697 = t19696 ^ t19696;
    wire t19698 = t19697 ^ t19697;
    wire t19699 = t19698 ^ t19698;
    wire t19700 = t19699 ^ t19699;
    wire t19701 = t19700 ^ t19700;
    wire t19702 = t19701 ^ t19701;
    wire t19703 = t19702 ^ t19702;
    wire t19704 = t19703 ^ t19703;
    wire t19705 = t19704 ^ t19704;
    wire t19706 = t19705 ^ t19705;
    wire t19707 = t19706 ^ t19706;
    wire t19708 = t19707 ^ t19707;
    wire t19709 = t19708 ^ t19708;
    wire t19710 = t19709 ^ t19709;
    wire t19711 = t19710 ^ t19710;
    wire t19712 = t19711 ^ t19711;
    wire t19713 = t19712 ^ t19712;
    wire t19714 = t19713 ^ t19713;
    wire t19715 = t19714 ^ t19714;
    wire t19716 = t19715 ^ t19715;
    wire t19717 = t19716 ^ t19716;
    wire t19718 = t19717 ^ t19717;
    wire t19719 = t19718 ^ t19718;
    wire t19720 = t19719 ^ t19719;
    wire t19721 = t19720 ^ t19720;
    wire t19722 = t19721 ^ t19721;
    wire t19723 = t19722 ^ t19722;
    wire t19724 = t19723 ^ t19723;
    wire t19725 = t19724 ^ t19724;
    wire t19726 = t19725 ^ t19725;
    wire t19727 = t19726 ^ t19726;
    wire t19728 = t19727 ^ t19727;
    wire t19729 = t19728 ^ t19728;
    wire t19730 = t19729 ^ t19729;
    wire t19731 = t19730 ^ t19730;
    wire t19732 = t19731 ^ t19731;
    wire t19733 = t19732 ^ t19732;
    wire t19734 = t19733 ^ t19733;
    wire t19735 = t19734 ^ t19734;
    wire t19736 = t19735 ^ t19735;
    wire t19737 = t19736 ^ t19736;
    wire t19738 = t19737 ^ t19737;
    wire t19739 = t19738 ^ t19738;
    wire t19740 = t19739 ^ t19739;
    wire t19741 = t19740 ^ t19740;
    wire t19742 = t19741 ^ t19741;
    wire t19743 = t19742 ^ t19742;
    wire t19744 = t19743 ^ t19743;
    wire t19745 = t19744 ^ t19744;
    wire t19746 = t19745 ^ t19745;
    wire t19747 = t19746 ^ t19746;
    wire t19748 = t19747 ^ t19747;
    wire t19749 = t19748 ^ t19748;
    wire t19750 = t19749 ^ t19749;
    wire t19751 = t19750 ^ t19750;
    wire t19752 = t19751 ^ t19751;
    wire t19753 = t19752 ^ t19752;
    wire t19754 = t19753 ^ t19753;
    wire t19755 = t19754 ^ t19754;
    wire t19756 = t19755 ^ t19755;
    wire t19757 = t19756 ^ t19756;
    wire t19758 = t19757 ^ t19757;
    wire t19759 = t19758 ^ t19758;
    wire t19760 = t19759 ^ t19759;
    wire t19761 = t19760 ^ t19760;
    wire t19762 = t19761 ^ t19761;
    wire t19763 = t19762 ^ t19762;
    wire t19764 = t19763 ^ t19763;
    wire t19765 = t19764 ^ t19764;
    wire t19766 = t19765 ^ t19765;
    wire t19767 = t19766 ^ t19766;
    wire t19768 = t19767 ^ t19767;
    wire t19769 = t19768 ^ t19768;
    wire t19770 = t19769 ^ t19769;
    wire t19771 = t19770 ^ t19770;
    wire t19772 = t19771 ^ t19771;
    wire t19773 = t19772 ^ t19772;
    wire t19774 = t19773 ^ t19773;
    wire t19775 = t19774 ^ t19774;
    wire t19776 = t19775 ^ t19775;
    wire t19777 = t19776 ^ t19776;
    wire t19778 = t19777 ^ t19777;
    wire t19779 = t19778 ^ t19778;
    wire t19780 = t19779 ^ t19779;
    wire t19781 = t19780 ^ t19780;
    wire t19782 = t19781 ^ t19781;
    wire t19783 = t19782 ^ t19782;
    wire t19784 = t19783 ^ t19783;
    wire t19785 = t19784 ^ t19784;
    wire t19786 = t19785 ^ t19785;
    wire t19787 = t19786 ^ t19786;
    wire t19788 = t19787 ^ t19787;
    wire t19789 = t19788 ^ t19788;
    wire t19790 = t19789 ^ t19789;
    wire t19791 = t19790 ^ t19790;
    wire t19792 = t19791 ^ t19791;
    wire t19793 = t19792 ^ t19792;
    wire t19794 = t19793 ^ t19793;
    wire t19795 = t19794 ^ t19794;
    wire t19796 = t19795 ^ t19795;
    wire t19797 = t19796 ^ t19796;
    wire t19798 = t19797 ^ t19797;
    wire t19799 = t19798 ^ t19798;
    wire t19800 = t19799 ^ t19799;
    wire t19801 = t19800 ^ t19800;
    wire t19802 = t19801 ^ t19801;
    wire t19803 = t19802 ^ t19802;
    wire t19804 = t19803 ^ t19803;
    wire t19805 = t19804 ^ t19804;
    wire t19806 = t19805 ^ t19805;
    wire t19807 = t19806 ^ t19806;
    wire t19808 = t19807 ^ t19807;
    wire t19809 = t19808 ^ t19808;
    wire t19810 = t19809 ^ t19809;
    wire t19811 = t19810 ^ t19810;
    wire t19812 = t19811 ^ t19811;
    wire t19813 = t19812 ^ t19812;
    wire t19814 = t19813 ^ t19813;
    wire t19815 = t19814 ^ t19814;
    wire t19816 = t19815 ^ t19815;
    wire t19817 = t19816 ^ t19816;
    wire t19818 = t19817 ^ t19817;
    wire t19819 = t19818 ^ t19818;
    wire t19820 = t19819 ^ t19819;
    wire t19821 = t19820 ^ t19820;
    wire t19822 = t19821 ^ t19821;
    wire t19823 = t19822 ^ t19822;
    wire t19824 = t19823 ^ t19823;
    wire t19825 = t19824 ^ t19824;
    wire t19826 = t19825 ^ t19825;
    wire t19827 = t19826 ^ t19826;
    wire t19828 = t19827 ^ t19827;
    wire t19829 = t19828 ^ t19828;
    wire t19830 = t19829 ^ t19829;
    wire t19831 = t19830 ^ t19830;
    wire t19832 = t19831 ^ t19831;
    wire t19833 = t19832 ^ t19832;
    wire t19834 = t19833 ^ t19833;
    wire t19835 = t19834 ^ t19834;
    wire t19836 = t19835 ^ t19835;
    wire t19837 = t19836 ^ t19836;
    wire t19838 = t19837 ^ t19837;
    wire t19839 = t19838 ^ t19838;
    wire t19840 = t19839 ^ t19839;
    wire t19841 = t19840 ^ t19840;
    wire t19842 = t19841 ^ t19841;
    wire t19843 = t19842 ^ t19842;
    wire t19844 = t19843 ^ t19843;
    wire t19845 = t19844 ^ t19844;
    wire t19846 = t19845 ^ t19845;
    wire t19847 = t19846 ^ t19846;
    wire t19848 = t19847 ^ t19847;
    wire t19849 = t19848 ^ t19848;
    wire t19850 = t19849 ^ t19849;
    wire t19851 = t19850 ^ t19850;
    wire t19852 = t19851 ^ t19851;
    wire t19853 = t19852 ^ t19852;
    wire t19854 = t19853 ^ t19853;
    wire t19855 = t19854 ^ t19854;
    wire t19856 = t19855 ^ t19855;
    wire t19857 = t19856 ^ t19856;
    wire t19858 = t19857 ^ t19857;
    wire t19859 = t19858 ^ t19858;
    wire t19860 = t19859 ^ t19859;
    wire t19861 = t19860 ^ t19860;
    wire t19862 = t19861 ^ t19861;
    wire t19863 = t19862 ^ t19862;
    wire t19864 = t19863 ^ t19863;
    wire t19865 = t19864 ^ t19864;
    wire t19866 = t19865 ^ t19865;
    wire t19867 = t19866 ^ t19866;
    wire t19868 = t19867 ^ t19867;
    wire t19869 = t19868 ^ t19868;
    wire t19870 = t19869 ^ t19869;
    wire t19871 = t19870 ^ t19870;
    wire t19872 = t19871 ^ t19871;
    wire t19873 = t19872 ^ t19872;
    wire t19874 = t19873 ^ t19873;
    wire t19875 = t19874 ^ t19874;
    wire t19876 = t19875 ^ t19875;
    wire t19877 = t19876 ^ t19876;
    wire t19878 = t19877 ^ t19877;
    wire t19879 = t19878 ^ t19878;
    wire t19880 = t19879 ^ t19879;
    wire t19881 = t19880 ^ t19880;
    wire t19882 = t19881 ^ t19881;
    wire t19883 = t19882 ^ t19882;
    wire t19884 = t19883 ^ t19883;
    wire t19885 = t19884 ^ t19884;
    wire t19886 = t19885 ^ t19885;
    wire t19887 = t19886 ^ t19886;
    wire t19888 = t19887 ^ t19887;
    wire t19889 = t19888 ^ t19888;
    wire t19890 = t19889 ^ t19889;
    wire t19891 = t19890 ^ t19890;
    wire t19892 = t19891 ^ t19891;
    wire t19893 = t19892 ^ t19892;
    wire t19894 = t19893 ^ t19893;
    wire t19895 = t19894 ^ t19894;
    wire t19896 = t19895 ^ t19895;
    wire t19897 = t19896 ^ t19896;
    wire t19898 = t19897 ^ t19897;
    wire t19899 = t19898 ^ t19898;
    wire t19900 = t19899 ^ t19899;
    wire t19901 = t19900 ^ t19900;
    wire t19902 = t19901 ^ t19901;
    wire t19903 = t19902 ^ t19902;
    wire t19904 = t19903 ^ t19903;
    wire t19905 = t19904 ^ t19904;
    wire t19906 = t19905 ^ t19905;
    wire t19907 = t19906 ^ t19906;
    wire t19908 = t19907 ^ t19907;
    wire t19909 = t19908 ^ t19908;
    wire t19910 = t19909 ^ t19909;
    wire t19911 = t19910 ^ t19910;
    wire t19912 = t19911 ^ t19911;
    wire t19913 = t19912 ^ t19912;
    wire t19914 = t19913 ^ t19913;
    wire t19915 = t19914 ^ t19914;
    wire t19916 = t19915 ^ t19915;
    wire t19917 = t19916 ^ t19916;
    wire t19918 = t19917 ^ t19917;
    wire t19919 = t19918 ^ t19918;
    wire t19920 = t19919 ^ t19919;
    wire t19921 = t19920 ^ t19920;
    wire t19922 = t19921 ^ t19921;
    wire t19923 = t19922 ^ t19922;
    wire t19924 = t19923 ^ t19923;
    wire t19925 = t19924 ^ t19924;
    wire t19926 = t19925 ^ t19925;
    wire t19927 = t19926 ^ t19926;
    wire t19928 = t19927 ^ t19927;
    wire t19929 = t19928 ^ t19928;
    wire t19930 = t19929 ^ t19929;
    wire t19931 = t19930 ^ t19930;
    wire t19932 = t19931 ^ t19931;
    wire t19933 = t19932 ^ t19932;
    wire t19934 = t19933 ^ t19933;
    wire t19935 = t19934 ^ t19934;
    wire t19936 = t19935 ^ t19935;
    wire t19937 = t19936 ^ t19936;
    wire t19938 = t19937 ^ t19937;
    wire t19939 = t19938 ^ t19938;
    wire t19940 = t19939 ^ t19939;
    wire t19941 = t19940 ^ t19940;
    wire t19942 = t19941 ^ t19941;
    wire t19943 = t19942 ^ t19942;
    wire t19944 = t19943 ^ t19943;
    wire t19945 = t19944 ^ t19944;
    wire t19946 = t19945 ^ t19945;
    wire t19947 = t19946 ^ t19946;
    wire t19948 = t19947 ^ t19947;
    wire t19949 = t19948 ^ t19948;
    wire t19950 = t19949 ^ t19949;
    wire t19951 = t19950 ^ t19950;
    wire t19952 = t19951 ^ t19951;
    wire t19953 = t19952 ^ t19952;
    wire t19954 = t19953 ^ t19953;
    wire t19955 = t19954 ^ t19954;
    wire t19956 = t19955 ^ t19955;
    wire t19957 = t19956 ^ t19956;
    wire t19958 = t19957 ^ t19957;
    wire t19959 = t19958 ^ t19958;
    wire t19960 = t19959 ^ t19959;
    wire t19961 = t19960 ^ t19960;
    wire t19962 = t19961 ^ t19961;
    wire t19963 = t19962 ^ t19962;
    wire t19964 = t19963 ^ t19963;
    wire t19965 = t19964 ^ t19964;
    wire t19966 = t19965 ^ t19965;
    wire t19967 = t19966 ^ t19966;
    wire t19968 = t19967 ^ t19967;
    wire t19969 = t19968 ^ t19968;
    wire t19970 = t19969 ^ t19969;
    wire t19971 = t19970 ^ t19970;
    wire t19972 = t19971 ^ t19971;
    wire t19973 = t19972 ^ t19972;
    wire t19974 = t19973 ^ t19973;
    wire t19975 = t19974 ^ t19974;
    wire t19976 = t19975 ^ t19975;
    wire t19977 = t19976 ^ t19976;
    wire t19978 = t19977 ^ t19977;
    wire t19979 = t19978 ^ t19978;
    wire t19980 = t19979 ^ t19979;
    wire t19981 = t19980 ^ t19980;
    wire t19982 = t19981 ^ t19981;
    wire t19983 = t19982 ^ t19982;
    wire t19984 = t19983 ^ t19983;
    wire t19985 = t19984 ^ t19984;
    wire t19986 = t19985 ^ t19985;
    wire t19987 = t19986 ^ t19986;
    wire t19988 = t19987 ^ t19987;
    wire t19989 = t19988 ^ t19988;
    wire t19990 = t19989 ^ t19989;
    wire t19991 = t19990 ^ t19990;
    wire t19992 = t19991 ^ t19991;
    wire t19993 = t19992 ^ t19992;
    wire t19994 = t19993 ^ t19993;
    wire t19995 = t19994 ^ t19994;
    wire t19996 = t19995 ^ t19995;
    wire t19997 = t19996 ^ t19996;
    wire t19998 = t19997 ^ t19997;
    wire t19999 = t19998 ^ t19998;
    wire t20000 = t19999 ^ t19999;
    wire t20001 = t20000 ^ t20000;
    wire t20002 = t20001 ^ t20001;
    wire t20003 = t20002 ^ t20002;
    wire t20004 = t20003 ^ t20003;
    wire t20005 = t20004 ^ t20004;
    wire t20006 = t20005 ^ t20005;
    wire t20007 = t20006 ^ t20006;
    wire t20008 = t20007 ^ t20007;
    wire t20009 = t20008 ^ t20008;
    wire t20010 = t20009 ^ t20009;
    wire t20011 = t20010 ^ t20010;
    wire t20012 = t20011 ^ t20011;
    wire t20013 = t20012 ^ t20012;
    wire t20014 = t20013 ^ t20013;
    wire t20015 = t20014 ^ t20014;
    wire t20016 = t20015 ^ t20015;
    wire t20017 = t20016 ^ t20016;
    wire t20018 = t20017 ^ t20017;
    wire t20019 = t20018 ^ t20018;
    wire t20020 = t20019 ^ t20019;
    wire t20021 = t20020 ^ t20020;
    wire t20022 = t20021 ^ t20021;
    wire t20023 = t20022 ^ t20022;
    wire t20024 = t20023 ^ t20023;
    wire t20025 = t20024 ^ t20024;
    wire t20026 = t20025 ^ t20025;
    wire t20027 = t20026 ^ t20026;
    wire t20028 = t20027 ^ t20027;
    wire t20029 = t20028 ^ t20028;
    wire t20030 = t20029 ^ t20029;
    wire t20031 = t20030 ^ t20030;
    wire t20032 = t20031 ^ t20031;
    wire t20033 = t20032 ^ t20032;
    wire t20034 = t20033 ^ t20033;
    wire t20035 = t20034 ^ t20034;
    wire t20036 = t20035 ^ t20035;
    wire t20037 = t20036 ^ t20036;
    wire t20038 = t20037 ^ t20037;
    wire t20039 = t20038 ^ t20038;
    wire t20040 = t20039 ^ t20039;
    wire t20041 = t20040 ^ t20040;
    wire t20042 = t20041 ^ t20041;
    wire t20043 = t20042 ^ t20042;
    wire t20044 = t20043 ^ t20043;
    wire t20045 = t20044 ^ t20044;
    wire t20046 = t20045 ^ t20045;
    wire t20047 = t20046 ^ t20046;
    wire t20048 = t20047 ^ t20047;
    wire t20049 = t20048 ^ t20048;
    wire t20050 = t20049 ^ t20049;
    wire t20051 = t20050 ^ t20050;
    wire t20052 = t20051 ^ t20051;
    wire t20053 = t20052 ^ t20052;
    wire t20054 = t20053 ^ t20053;
    wire t20055 = t20054 ^ t20054;
    wire t20056 = t20055 ^ t20055;
    wire t20057 = t20056 ^ t20056;
    wire t20058 = t20057 ^ t20057;
    wire t20059 = t20058 ^ t20058;
    wire t20060 = t20059 ^ t20059;
    wire t20061 = t20060 ^ t20060;
    wire t20062 = t20061 ^ t20061;
    wire t20063 = t20062 ^ t20062;
    wire t20064 = t20063 ^ t20063;
    wire t20065 = t20064 ^ t20064;
    wire t20066 = t20065 ^ t20065;
    wire t20067 = t20066 ^ t20066;
    wire t20068 = t20067 ^ t20067;
    wire t20069 = t20068 ^ t20068;
    wire t20070 = t20069 ^ t20069;
    wire t20071 = t20070 ^ t20070;
    wire t20072 = t20071 ^ t20071;
    wire t20073 = t20072 ^ t20072;
    wire t20074 = t20073 ^ t20073;
    wire t20075 = t20074 ^ t20074;
    wire t20076 = t20075 ^ t20075;
    wire t20077 = t20076 ^ t20076;
    wire t20078 = t20077 ^ t20077;
    wire t20079 = t20078 ^ t20078;
    wire t20080 = t20079 ^ t20079;
    wire t20081 = t20080 ^ t20080;
    wire t20082 = t20081 ^ t20081;
    wire t20083 = t20082 ^ t20082;
    wire t20084 = t20083 ^ t20083;
    wire t20085 = t20084 ^ t20084;
    wire t20086 = t20085 ^ t20085;
    wire t20087 = t20086 ^ t20086;
    wire t20088 = t20087 ^ t20087;
    wire t20089 = t20088 ^ t20088;
    wire t20090 = t20089 ^ t20089;
    wire t20091 = t20090 ^ t20090;
    wire t20092 = t20091 ^ t20091;
    wire t20093 = t20092 ^ t20092;
    wire t20094 = t20093 ^ t20093;
    wire t20095 = t20094 ^ t20094;
    wire t20096 = t20095 ^ t20095;
    wire t20097 = t20096 ^ t20096;
    wire t20098 = t20097 ^ t20097;
    wire t20099 = t20098 ^ t20098;
    wire t20100 = t20099 ^ t20099;
    wire t20101 = t20100 ^ t20100;
    wire t20102 = t20101 ^ t20101;
    wire t20103 = t20102 ^ t20102;
    wire t20104 = t20103 ^ t20103;
    wire t20105 = t20104 ^ t20104;
    wire t20106 = t20105 ^ t20105;
    wire t20107 = t20106 ^ t20106;
    wire t20108 = t20107 ^ t20107;
    wire t20109 = t20108 ^ t20108;
    wire t20110 = t20109 ^ t20109;
    wire t20111 = t20110 ^ t20110;
    wire t20112 = t20111 ^ t20111;
    wire t20113 = t20112 ^ t20112;
    wire t20114 = t20113 ^ t20113;
    wire t20115 = t20114 ^ t20114;
    wire t20116 = t20115 ^ t20115;
    wire t20117 = t20116 ^ t20116;
    wire t20118 = t20117 ^ t20117;
    wire t20119 = t20118 ^ t20118;
    wire t20120 = t20119 ^ t20119;
    wire t20121 = t20120 ^ t20120;
    wire t20122 = t20121 ^ t20121;
    wire t20123 = t20122 ^ t20122;
    wire t20124 = t20123 ^ t20123;
    wire t20125 = t20124 ^ t20124;
    wire t20126 = t20125 ^ t20125;
    wire t20127 = t20126 ^ t20126;
    wire t20128 = t20127 ^ t20127;
    wire t20129 = t20128 ^ t20128;
    wire t20130 = t20129 ^ t20129;
    wire t20131 = t20130 ^ t20130;
    wire t20132 = t20131 ^ t20131;
    wire t20133 = t20132 ^ t20132;
    wire t20134 = t20133 ^ t20133;
    wire t20135 = t20134 ^ t20134;
    wire t20136 = t20135 ^ t20135;
    wire t20137 = t20136 ^ t20136;
    wire t20138 = t20137 ^ t20137;
    wire t20139 = t20138 ^ t20138;
    wire t20140 = t20139 ^ t20139;
    wire t20141 = t20140 ^ t20140;
    wire t20142 = t20141 ^ t20141;
    wire t20143 = t20142 ^ t20142;
    wire t20144 = t20143 ^ t20143;
    wire t20145 = t20144 ^ t20144;
    wire t20146 = t20145 ^ t20145;
    wire t20147 = t20146 ^ t20146;
    wire t20148 = t20147 ^ t20147;
    wire t20149 = t20148 ^ t20148;
    wire t20150 = t20149 ^ t20149;
    wire t20151 = t20150 ^ t20150;
    wire t20152 = t20151 ^ t20151;
    wire t20153 = t20152 ^ t20152;
    wire t20154 = t20153 ^ t20153;
    wire t20155 = t20154 ^ t20154;
    wire t20156 = t20155 ^ t20155;
    wire t20157 = t20156 ^ t20156;
    wire t20158 = t20157 ^ t20157;
    wire t20159 = t20158 ^ t20158;
    wire t20160 = t20159 ^ t20159;
    wire t20161 = t20160 ^ t20160;
    wire t20162 = t20161 ^ t20161;
    wire t20163 = t20162 ^ t20162;
    wire t20164 = t20163 ^ t20163;
    wire t20165 = t20164 ^ t20164;
    wire t20166 = t20165 ^ t20165;
    wire t20167 = t20166 ^ t20166;
    wire t20168 = t20167 ^ t20167;
    wire t20169 = t20168 ^ t20168;
    wire t20170 = t20169 ^ t20169;
    wire t20171 = t20170 ^ t20170;
    wire t20172 = t20171 ^ t20171;
    wire t20173 = t20172 ^ t20172;
    wire t20174 = t20173 ^ t20173;
    wire t20175 = t20174 ^ t20174;
    wire t20176 = t20175 ^ t20175;
    wire t20177 = t20176 ^ t20176;
    wire t20178 = t20177 ^ t20177;
    wire t20179 = t20178 ^ t20178;
    wire t20180 = t20179 ^ t20179;
    wire t20181 = t20180 ^ t20180;
    wire t20182 = t20181 ^ t20181;
    wire t20183 = t20182 ^ t20182;
    wire t20184 = t20183 ^ t20183;
    wire t20185 = t20184 ^ t20184;
    wire t20186 = t20185 ^ t20185;
    wire t20187 = t20186 ^ t20186;
    wire t20188 = t20187 ^ t20187;
    wire t20189 = t20188 ^ t20188;
    wire t20190 = t20189 ^ t20189;
    wire t20191 = t20190 ^ t20190;
    wire t20192 = t20191 ^ t20191;
    wire t20193 = t20192 ^ t20192;
    wire t20194 = t20193 ^ t20193;
    wire t20195 = t20194 ^ t20194;
    wire t20196 = t20195 ^ t20195;
    wire t20197 = t20196 ^ t20196;
    wire t20198 = t20197 ^ t20197;
    wire t20199 = t20198 ^ t20198;
    wire t20200 = t20199 ^ t20199;
    wire t20201 = t20200 ^ t20200;
    wire t20202 = t20201 ^ t20201;
    wire t20203 = t20202 ^ t20202;
    wire t20204 = t20203 ^ t20203;
    wire t20205 = t20204 ^ t20204;
    wire t20206 = t20205 ^ t20205;
    wire t20207 = t20206 ^ t20206;
    wire t20208 = t20207 ^ t20207;
    wire t20209 = t20208 ^ t20208;
    wire t20210 = t20209 ^ t20209;
    wire t20211 = t20210 ^ t20210;
    wire t20212 = t20211 ^ t20211;
    wire t20213 = t20212 ^ t20212;
    wire t20214 = t20213 ^ t20213;
    wire t20215 = t20214 ^ t20214;
    wire t20216 = t20215 ^ t20215;
    wire t20217 = t20216 ^ t20216;
    wire t20218 = t20217 ^ t20217;
    wire t20219 = t20218 ^ t20218;
    wire t20220 = t20219 ^ t20219;
    wire t20221 = t20220 ^ t20220;
    wire t20222 = t20221 ^ t20221;
    wire t20223 = t20222 ^ t20222;
    wire t20224 = t20223 ^ t20223;
    wire t20225 = t20224 ^ t20224;
    wire t20226 = t20225 ^ t20225;
    wire t20227 = t20226 ^ t20226;
    wire t20228 = t20227 ^ t20227;
    wire t20229 = t20228 ^ t20228;
    wire t20230 = t20229 ^ t20229;
    wire t20231 = t20230 ^ t20230;
    wire t20232 = t20231 ^ t20231;
    wire t20233 = t20232 ^ t20232;
    wire t20234 = t20233 ^ t20233;
    wire t20235 = t20234 ^ t20234;
    wire t20236 = t20235 ^ t20235;
    wire t20237 = t20236 ^ t20236;
    wire t20238 = t20237 ^ t20237;
    wire t20239 = t20238 ^ t20238;
    wire t20240 = t20239 ^ t20239;
    wire t20241 = t20240 ^ t20240;
    wire t20242 = t20241 ^ t20241;
    wire t20243 = t20242 ^ t20242;
    wire t20244 = t20243 ^ t20243;
    wire t20245 = t20244 ^ t20244;
    wire t20246 = t20245 ^ t20245;
    wire t20247 = t20246 ^ t20246;
    wire t20248 = t20247 ^ t20247;
    wire t20249 = t20248 ^ t20248;
    wire t20250 = t20249 ^ t20249;
    wire t20251 = t20250 ^ t20250;
    wire t20252 = t20251 ^ t20251;
    wire t20253 = t20252 ^ t20252;
    wire t20254 = t20253 ^ t20253;
    wire t20255 = t20254 ^ t20254;
    wire t20256 = t20255 ^ t20255;
    wire t20257 = t20256 ^ t20256;
    wire t20258 = t20257 ^ t20257;
    wire t20259 = t20258 ^ t20258;
    wire t20260 = t20259 ^ t20259;
    wire t20261 = t20260 ^ t20260;
    wire t20262 = t20261 ^ t20261;
    wire t20263 = t20262 ^ t20262;
    wire t20264 = t20263 ^ t20263;
    wire t20265 = t20264 ^ t20264;
    wire t20266 = t20265 ^ t20265;
    wire t20267 = t20266 ^ t20266;
    wire t20268 = t20267 ^ t20267;
    wire t20269 = t20268 ^ t20268;
    wire t20270 = t20269 ^ t20269;
    wire t20271 = t20270 ^ t20270;
    wire t20272 = t20271 ^ t20271;
    wire t20273 = t20272 ^ t20272;
    wire t20274 = t20273 ^ t20273;
    wire t20275 = t20274 ^ t20274;
    wire t20276 = t20275 ^ t20275;
    wire t20277 = t20276 ^ t20276;
    wire t20278 = t20277 ^ t20277;
    wire t20279 = t20278 ^ t20278;
    wire t20280 = t20279 ^ t20279;
    wire t20281 = t20280 ^ t20280;
    wire t20282 = t20281 ^ t20281;
    wire t20283 = t20282 ^ t20282;
    wire t20284 = t20283 ^ t20283;
    wire t20285 = t20284 ^ t20284;
    wire t20286 = t20285 ^ t20285;
    wire t20287 = t20286 ^ t20286;
    wire t20288 = t20287 ^ t20287;
    wire t20289 = t20288 ^ t20288;
    wire t20290 = t20289 ^ t20289;
    wire t20291 = t20290 ^ t20290;
    wire t20292 = t20291 ^ t20291;
    wire t20293 = t20292 ^ t20292;
    wire t20294 = t20293 ^ t20293;
    wire t20295 = t20294 ^ t20294;
    wire t20296 = t20295 ^ t20295;
    wire t20297 = t20296 ^ t20296;
    wire t20298 = t20297 ^ t20297;
    wire t20299 = t20298 ^ t20298;
    wire t20300 = t20299 ^ t20299;
    wire t20301 = t20300 ^ t20300;
    wire t20302 = t20301 ^ t20301;
    wire t20303 = t20302 ^ t20302;
    wire t20304 = t20303 ^ t20303;
    wire t20305 = t20304 ^ t20304;
    wire t20306 = t20305 ^ t20305;
    wire t20307 = t20306 ^ t20306;
    wire t20308 = t20307 ^ t20307;
    wire t20309 = t20308 ^ t20308;
    wire t20310 = t20309 ^ t20309;
    wire t20311 = t20310 ^ t20310;
    wire t20312 = t20311 ^ t20311;
    wire t20313 = t20312 ^ t20312;
    wire t20314 = t20313 ^ t20313;
    wire t20315 = t20314 ^ t20314;
    wire t20316 = t20315 ^ t20315;
    wire t20317 = t20316 ^ t20316;
    wire t20318 = t20317 ^ t20317;
    wire t20319 = t20318 ^ t20318;
    wire t20320 = t20319 ^ t20319;
    wire t20321 = t20320 ^ t20320;
    wire t20322 = t20321 ^ t20321;
    wire t20323 = t20322 ^ t20322;
    wire t20324 = t20323 ^ t20323;
    wire t20325 = t20324 ^ t20324;
    wire t20326 = t20325 ^ t20325;
    wire t20327 = t20326 ^ t20326;
    wire t20328 = t20327 ^ t20327;
    wire t20329 = t20328 ^ t20328;
    wire t20330 = t20329 ^ t20329;
    wire t20331 = t20330 ^ t20330;
    wire t20332 = t20331 ^ t20331;
    wire t20333 = t20332 ^ t20332;
    wire t20334 = t20333 ^ t20333;
    wire t20335 = t20334 ^ t20334;
    wire t20336 = t20335 ^ t20335;
    wire t20337 = t20336 ^ t20336;
    wire t20338 = t20337 ^ t20337;
    wire t20339 = t20338 ^ t20338;
    wire t20340 = t20339 ^ t20339;
    wire t20341 = t20340 ^ t20340;
    wire t20342 = t20341 ^ t20341;
    wire t20343 = t20342 ^ t20342;
    wire t20344 = t20343 ^ t20343;
    wire t20345 = t20344 ^ t20344;
    wire t20346 = t20345 ^ t20345;
    wire t20347 = t20346 ^ t20346;
    wire t20348 = t20347 ^ t20347;
    wire t20349 = t20348 ^ t20348;
    wire t20350 = t20349 ^ t20349;
    wire t20351 = t20350 ^ t20350;
    wire t20352 = t20351 ^ t20351;
    wire t20353 = t20352 ^ t20352;
    wire t20354 = t20353 ^ t20353;
    wire t20355 = t20354 ^ t20354;
    wire t20356 = t20355 ^ t20355;
    wire t20357 = t20356 ^ t20356;
    wire t20358 = t20357 ^ t20357;
    wire t20359 = t20358 ^ t20358;
    wire t20360 = t20359 ^ t20359;
    wire t20361 = t20360 ^ t20360;
    wire t20362 = t20361 ^ t20361;
    wire t20363 = t20362 ^ t20362;
    wire t20364 = t20363 ^ t20363;
    wire t20365 = t20364 ^ t20364;
    wire t20366 = t20365 ^ t20365;
    wire t20367 = t20366 ^ t20366;
    wire t20368 = t20367 ^ t20367;
    wire t20369 = t20368 ^ t20368;
    wire t20370 = t20369 ^ t20369;
    wire t20371 = t20370 ^ t20370;
    wire t20372 = t20371 ^ t20371;
    wire t20373 = t20372 ^ t20372;
    wire t20374 = t20373 ^ t20373;
    wire t20375 = t20374 ^ t20374;
    wire t20376 = t20375 ^ t20375;
    wire t20377 = t20376 ^ t20376;
    wire t20378 = t20377 ^ t20377;
    wire t20379 = t20378 ^ t20378;
    wire t20380 = t20379 ^ t20379;
    wire t20381 = t20380 ^ t20380;
    wire t20382 = t20381 ^ t20381;
    wire t20383 = t20382 ^ t20382;
    wire t20384 = t20383 ^ t20383;
    wire t20385 = t20384 ^ t20384;
    wire t20386 = t20385 ^ t20385;
    wire t20387 = t20386 ^ t20386;
    wire t20388 = t20387 ^ t20387;
    wire t20389 = t20388 ^ t20388;
    wire t20390 = t20389 ^ t20389;
    wire t20391 = t20390 ^ t20390;
    wire t20392 = t20391 ^ t20391;
    wire t20393 = t20392 ^ t20392;
    wire t20394 = t20393 ^ t20393;
    wire t20395 = t20394 ^ t20394;
    wire t20396 = t20395 ^ t20395;
    wire t20397 = t20396 ^ t20396;
    wire t20398 = t20397 ^ t20397;
    wire t20399 = t20398 ^ t20398;
    wire t20400 = t20399 ^ t20399;
    wire t20401 = t20400 ^ t20400;
    wire t20402 = t20401 ^ t20401;
    wire t20403 = t20402 ^ t20402;
    wire t20404 = t20403 ^ t20403;
    wire t20405 = t20404 ^ t20404;
    wire t20406 = t20405 ^ t20405;
    wire t20407 = t20406 ^ t20406;
    wire t20408 = t20407 ^ t20407;
    wire t20409 = t20408 ^ t20408;
    wire t20410 = t20409 ^ t20409;
    wire t20411 = t20410 ^ t20410;
    wire t20412 = t20411 ^ t20411;
    wire t20413 = t20412 ^ t20412;
    wire t20414 = t20413 ^ t20413;
    wire t20415 = t20414 ^ t20414;
    wire t20416 = t20415 ^ t20415;
    wire t20417 = t20416 ^ t20416;
    wire t20418 = t20417 ^ t20417;
    wire t20419 = t20418 ^ t20418;
    wire t20420 = t20419 ^ t20419;
    wire t20421 = t20420 ^ t20420;
    wire t20422 = t20421 ^ t20421;
    wire t20423 = t20422 ^ t20422;
    wire t20424 = t20423 ^ t20423;
    wire t20425 = t20424 ^ t20424;
    wire t20426 = t20425 ^ t20425;
    wire t20427 = t20426 ^ t20426;
    wire t20428 = t20427 ^ t20427;
    wire t20429 = t20428 ^ t20428;
    wire t20430 = t20429 ^ t20429;
    wire t20431 = t20430 ^ t20430;
    wire t20432 = t20431 ^ t20431;
    wire t20433 = t20432 ^ t20432;
    wire t20434 = t20433 ^ t20433;
    wire t20435 = t20434 ^ t20434;
    wire t20436 = t20435 ^ t20435;
    wire t20437 = t20436 ^ t20436;
    wire t20438 = t20437 ^ t20437;
    wire t20439 = t20438 ^ t20438;
    wire t20440 = t20439 ^ t20439;
    wire t20441 = t20440 ^ t20440;
    wire t20442 = t20441 ^ t20441;
    wire t20443 = t20442 ^ t20442;
    wire t20444 = t20443 ^ t20443;
    wire t20445 = t20444 ^ t20444;
    wire t20446 = t20445 ^ t20445;
    wire t20447 = t20446 ^ t20446;
    wire t20448 = t20447 ^ t20447;
    wire t20449 = t20448 ^ t20448;
    wire t20450 = t20449 ^ t20449;
    wire t20451 = t20450 ^ t20450;
    wire t20452 = t20451 ^ t20451;
    wire t20453 = t20452 ^ t20452;
    wire t20454 = t20453 ^ t20453;
    wire t20455 = t20454 ^ t20454;
    wire t20456 = t20455 ^ t20455;
    wire t20457 = t20456 ^ t20456;
    wire t20458 = t20457 ^ t20457;
    wire t20459 = t20458 ^ t20458;
    wire t20460 = t20459 ^ t20459;
    wire t20461 = t20460 ^ t20460;
    wire t20462 = t20461 ^ t20461;
    wire t20463 = t20462 ^ t20462;
    wire t20464 = t20463 ^ t20463;
    wire t20465 = t20464 ^ t20464;
    wire t20466 = t20465 ^ t20465;
    wire t20467 = t20466 ^ t20466;
    wire t20468 = t20467 ^ t20467;
    wire t20469 = t20468 ^ t20468;
    wire t20470 = t20469 ^ t20469;
    wire t20471 = t20470 ^ t20470;
    wire t20472 = t20471 ^ t20471;
    wire t20473 = t20472 ^ t20472;
    wire t20474 = t20473 ^ t20473;
    wire t20475 = t20474 ^ t20474;
    wire t20476 = t20475 ^ t20475;
    wire t20477 = t20476 ^ t20476;
    wire t20478 = t20477 ^ t20477;
    wire t20479 = t20478 ^ t20478;
    wire t20480 = t20479 ^ t20479;
    wire t20481 = t20480 ^ t20480;
    wire t20482 = t20481 ^ t20481;
    wire t20483 = t20482 ^ t20482;
    wire t20484 = t20483 ^ t20483;
    wire t20485 = t20484 ^ t20484;
    wire t20486 = t20485 ^ t20485;
    wire t20487 = t20486 ^ t20486;
    wire t20488 = t20487 ^ t20487;
    wire t20489 = t20488 ^ t20488;
    wire t20490 = t20489 ^ t20489;
    wire t20491 = t20490 ^ t20490;
    wire t20492 = t20491 ^ t20491;
    wire t20493 = t20492 ^ t20492;
    wire t20494 = t20493 ^ t20493;
    wire t20495 = t20494 ^ t20494;
    wire t20496 = t20495 ^ t20495;
    wire t20497 = t20496 ^ t20496;
    wire t20498 = t20497 ^ t20497;
    wire t20499 = t20498 ^ t20498;
    wire t20500 = t20499 ^ t20499;
    wire t20501 = t20500 ^ t20500;
    wire t20502 = t20501 ^ t20501;
    wire t20503 = t20502 ^ t20502;
    wire t20504 = t20503 ^ t20503;
    wire t20505 = t20504 ^ t20504;
    wire t20506 = t20505 ^ t20505;
    wire t20507 = t20506 ^ t20506;
    wire t20508 = t20507 ^ t20507;
    wire t20509 = t20508 ^ t20508;
    wire t20510 = t20509 ^ t20509;
    wire t20511 = t20510 ^ t20510;
    wire t20512 = t20511 ^ t20511;
    wire t20513 = t20512 ^ t20512;
    wire t20514 = t20513 ^ t20513;
    wire t20515 = t20514 ^ t20514;
    wire t20516 = t20515 ^ t20515;
    wire t20517 = t20516 ^ t20516;
    wire t20518 = t20517 ^ t20517;
    wire t20519 = t20518 ^ t20518;
    wire t20520 = t20519 ^ t20519;
    wire t20521 = t20520 ^ t20520;
    wire t20522 = t20521 ^ t20521;
    wire t20523 = t20522 ^ t20522;
    wire t20524 = t20523 ^ t20523;
    wire t20525 = t20524 ^ t20524;
    wire t20526 = t20525 ^ t20525;
    wire t20527 = t20526 ^ t20526;
    wire t20528 = t20527 ^ t20527;
    wire t20529 = t20528 ^ t20528;
    wire t20530 = t20529 ^ t20529;
    wire t20531 = t20530 ^ t20530;
    wire t20532 = t20531 ^ t20531;
    wire t20533 = t20532 ^ t20532;
    wire t20534 = t20533 ^ t20533;
    wire t20535 = t20534 ^ t20534;
    wire t20536 = t20535 ^ t20535;
    wire t20537 = t20536 ^ t20536;
    wire t20538 = t20537 ^ t20537;
    wire t20539 = t20538 ^ t20538;
    wire t20540 = t20539 ^ t20539;
    wire t20541 = t20540 ^ t20540;
    wire t20542 = t20541 ^ t20541;
    wire t20543 = t20542 ^ t20542;
    wire t20544 = t20543 ^ t20543;
    wire t20545 = t20544 ^ t20544;
    wire t20546 = t20545 ^ t20545;
    wire t20547 = t20546 ^ t20546;
    wire t20548 = t20547 ^ t20547;
    wire t20549 = t20548 ^ t20548;
    wire t20550 = t20549 ^ t20549;
    wire t20551 = t20550 ^ t20550;
    wire t20552 = t20551 ^ t20551;
    wire t20553 = t20552 ^ t20552;
    wire t20554 = t20553 ^ t20553;
    wire t20555 = t20554 ^ t20554;
    wire t20556 = t20555 ^ t20555;
    wire t20557 = t20556 ^ t20556;
    wire t20558 = t20557 ^ t20557;
    wire t20559 = t20558 ^ t20558;
    wire t20560 = t20559 ^ t20559;
    wire t20561 = t20560 ^ t20560;
    wire t20562 = t20561 ^ t20561;
    wire t20563 = t20562 ^ t20562;
    wire t20564 = t20563 ^ t20563;
    wire t20565 = t20564 ^ t20564;
    wire t20566 = t20565 ^ t20565;
    wire t20567 = t20566 ^ t20566;
    wire t20568 = t20567 ^ t20567;
    wire t20569 = t20568 ^ t20568;
    wire t20570 = t20569 ^ t20569;
    wire t20571 = t20570 ^ t20570;
    wire t20572 = t20571 ^ t20571;
    wire t20573 = t20572 ^ t20572;
    wire t20574 = t20573 ^ t20573;
    wire t20575 = t20574 ^ t20574;
    wire t20576 = t20575 ^ t20575;
    wire t20577 = t20576 ^ t20576;
    wire t20578 = t20577 ^ t20577;
    wire t20579 = t20578 ^ t20578;
    wire t20580 = t20579 ^ t20579;
    wire t20581 = t20580 ^ t20580;
    wire t20582 = t20581 ^ t20581;
    wire t20583 = t20582 ^ t20582;
    wire t20584 = t20583 ^ t20583;
    wire t20585 = t20584 ^ t20584;
    wire t20586 = t20585 ^ t20585;
    wire t20587 = t20586 ^ t20586;
    wire t20588 = t20587 ^ t20587;
    wire t20589 = t20588 ^ t20588;
    wire t20590 = t20589 ^ t20589;
    wire t20591 = t20590 ^ t20590;
    wire t20592 = t20591 ^ t20591;
    wire t20593 = t20592 ^ t20592;
    wire t20594 = t20593 ^ t20593;
    wire t20595 = t20594 ^ t20594;
    wire t20596 = t20595 ^ t20595;
    wire t20597 = t20596 ^ t20596;
    wire t20598 = t20597 ^ t20597;
    wire t20599 = t20598 ^ t20598;
    wire t20600 = t20599 ^ t20599;
    wire t20601 = t20600 ^ t20600;
    wire t20602 = t20601 ^ t20601;
    wire t20603 = t20602 ^ t20602;
    wire t20604 = t20603 ^ t20603;
    wire t20605 = t20604 ^ t20604;
    wire t20606 = t20605 ^ t20605;
    wire t20607 = t20606 ^ t20606;
    wire t20608 = t20607 ^ t20607;
    wire t20609 = t20608 ^ t20608;
    wire t20610 = t20609 ^ t20609;
    wire t20611 = t20610 ^ t20610;
    wire t20612 = t20611 ^ t20611;
    wire t20613 = t20612 ^ t20612;
    wire t20614 = t20613 ^ t20613;
    wire t20615 = t20614 ^ t20614;
    wire t20616 = t20615 ^ t20615;
    wire t20617 = t20616 ^ t20616;
    wire t20618 = t20617 ^ t20617;
    wire t20619 = t20618 ^ t20618;
    wire t20620 = t20619 ^ t20619;
    wire t20621 = t20620 ^ t20620;
    wire t20622 = t20621 ^ t20621;
    wire t20623 = t20622 ^ t20622;
    wire t20624 = t20623 ^ t20623;
    wire t20625 = t20624 ^ t20624;
    wire t20626 = t20625 ^ t20625;
    wire t20627 = t20626 ^ t20626;
    wire t20628 = t20627 ^ t20627;
    wire t20629 = t20628 ^ t20628;
    wire t20630 = t20629 ^ t20629;
    wire t20631 = t20630 ^ t20630;
    wire t20632 = t20631 ^ t20631;
    wire t20633 = t20632 ^ t20632;
    wire t20634 = t20633 ^ t20633;
    wire t20635 = t20634 ^ t20634;
    wire t20636 = t20635 ^ t20635;
    wire t20637 = t20636 ^ t20636;
    wire t20638 = t20637 ^ t20637;
    wire t20639 = t20638 ^ t20638;
    wire t20640 = t20639 ^ t20639;
    wire t20641 = t20640 ^ t20640;
    wire t20642 = t20641 ^ t20641;
    wire t20643 = t20642 ^ t20642;
    wire t20644 = t20643 ^ t20643;
    wire t20645 = t20644 ^ t20644;
    wire t20646 = t20645 ^ t20645;
    wire t20647 = t20646 ^ t20646;
    wire t20648 = t20647 ^ t20647;
    wire t20649 = t20648 ^ t20648;
    wire t20650 = t20649 ^ t20649;
    wire t20651 = t20650 ^ t20650;
    wire t20652 = t20651 ^ t20651;
    wire t20653 = t20652 ^ t20652;
    wire t20654 = t20653 ^ t20653;
    wire t20655 = t20654 ^ t20654;
    wire t20656 = t20655 ^ t20655;
    wire t20657 = t20656 ^ t20656;
    wire t20658 = t20657 ^ t20657;
    wire t20659 = t20658 ^ t20658;
    wire t20660 = t20659 ^ t20659;
    wire t20661 = t20660 ^ t20660;
    wire t20662 = t20661 ^ t20661;
    wire t20663 = t20662 ^ t20662;
    wire t20664 = t20663 ^ t20663;
    wire t20665 = t20664 ^ t20664;
    wire t20666 = t20665 ^ t20665;
    wire t20667 = t20666 ^ t20666;
    wire t20668 = t20667 ^ t20667;
    wire t20669 = t20668 ^ t20668;
    wire t20670 = t20669 ^ t20669;
    wire t20671 = t20670 ^ t20670;
    wire t20672 = t20671 ^ t20671;
    wire t20673 = t20672 ^ t20672;
    wire t20674 = t20673 ^ t20673;
    wire t20675 = t20674 ^ t20674;
    wire t20676 = t20675 ^ t20675;
    wire t20677 = t20676 ^ t20676;
    wire t20678 = t20677 ^ t20677;
    wire t20679 = t20678 ^ t20678;
    wire t20680 = t20679 ^ t20679;
    wire t20681 = t20680 ^ t20680;
    wire t20682 = t20681 ^ t20681;
    wire t20683 = t20682 ^ t20682;
    wire t20684 = t20683 ^ t20683;
    wire t20685 = t20684 ^ t20684;
    wire t20686 = t20685 ^ t20685;
    wire t20687 = t20686 ^ t20686;
    wire t20688 = t20687 ^ t20687;
    wire t20689 = t20688 ^ t20688;
    wire t20690 = t20689 ^ t20689;
    wire t20691 = t20690 ^ t20690;
    wire t20692 = t20691 ^ t20691;
    wire t20693 = t20692 ^ t20692;
    wire t20694 = t20693 ^ t20693;
    wire t20695 = t20694 ^ t20694;
    wire t20696 = t20695 ^ t20695;
    wire t20697 = t20696 ^ t20696;
    wire t20698 = t20697 ^ t20697;
    wire t20699 = t20698 ^ t20698;
    wire t20700 = t20699 ^ t20699;
    wire t20701 = t20700 ^ t20700;
    wire t20702 = t20701 ^ t20701;
    wire t20703 = t20702 ^ t20702;
    wire t20704 = t20703 ^ t20703;
    wire t20705 = t20704 ^ t20704;
    wire t20706 = t20705 ^ t20705;
    wire t20707 = t20706 ^ t20706;
    wire t20708 = t20707 ^ t20707;
    wire t20709 = t20708 ^ t20708;
    wire t20710 = t20709 ^ t20709;
    wire t20711 = t20710 ^ t20710;
    wire t20712 = t20711 ^ t20711;
    wire t20713 = t20712 ^ t20712;
    wire t20714 = t20713 ^ t20713;
    wire t20715 = t20714 ^ t20714;
    wire t20716 = t20715 ^ t20715;
    wire t20717 = t20716 ^ t20716;
    wire t20718 = t20717 ^ t20717;
    wire t20719 = t20718 ^ t20718;
    wire t20720 = t20719 ^ t20719;
    wire t20721 = t20720 ^ t20720;
    wire t20722 = t20721 ^ t20721;
    wire t20723 = t20722 ^ t20722;
    wire t20724 = t20723 ^ t20723;
    wire t20725 = t20724 ^ t20724;
    wire t20726 = t20725 ^ t20725;
    wire t20727 = t20726 ^ t20726;
    wire t20728 = t20727 ^ t20727;
    wire t20729 = t20728 ^ t20728;
    wire t20730 = t20729 ^ t20729;
    wire t20731 = t20730 ^ t20730;
    wire t20732 = t20731 ^ t20731;
    wire t20733 = t20732 ^ t20732;
    wire t20734 = t20733 ^ t20733;
    wire t20735 = t20734 ^ t20734;
    wire t20736 = t20735 ^ t20735;
    wire t20737 = t20736 ^ t20736;
    wire t20738 = t20737 ^ t20737;
    wire t20739 = t20738 ^ t20738;
    wire t20740 = t20739 ^ t20739;
    wire t20741 = t20740 ^ t20740;
    wire t20742 = t20741 ^ t20741;
    wire t20743 = t20742 ^ t20742;
    wire t20744 = t20743 ^ t20743;
    wire t20745 = t20744 ^ t20744;
    wire t20746 = t20745 ^ t20745;
    wire t20747 = t20746 ^ t20746;
    wire t20748 = t20747 ^ t20747;
    wire t20749 = t20748 ^ t20748;
    wire t20750 = t20749 ^ t20749;
    wire t20751 = t20750 ^ t20750;
    wire t20752 = t20751 ^ t20751;
    wire t20753 = t20752 ^ t20752;
    wire t20754 = t20753 ^ t20753;
    wire t20755 = t20754 ^ t20754;
    wire t20756 = t20755 ^ t20755;
    wire t20757 = t20756 ^ t20756;
    wire t20758 = t20757 ^ t20757;
    wire t20759 = t20758 ^ t20758;
    wire t20760 = t20759 ^ t20759;
    wire t20761 = t20760 ^ t20760;
    wire t20762 = t20761 ^ t20761;
    wire t20763 = t20762 ^ t20762;
    wire t20764 = t20763 ^ t20763;
    wire t20765 = t20764 ^ t20764;
    wire t20766 = t20765 ^ t20765;
    wire t20767 = t20766 ^ t20766;
    wire t20768 = t20767 ^ t20767;
    wire t20769 = t20768 ^ t20768;
    wire t20770 = t20769 ^ t20769;
    wire t20771 = t20770 ^ t20770;
    wire t20772 = t20771 ^ t20771;
    wire t20773 = t20772 ^ t20772;
    wire t20774 = t20773 ^ t20773;
    wire t20775 = t20774 ^ t20774;
    wire t20776 = t20775 ^ t20775;
    wire t20777 = t20776 ^ t20776;
    wire t20778 = t20777 ^ t20777;
    wire t20779 = t20778 ^ t20778;
    wire t20780 = t20779 ^ t20779;
    wire t20781 = t20780 ^ t20780;
    wire t20782 = t20781 ^ t20781;
    wire t20783 = t20782 ^ t20782;
    wire t20784 = t20783 ^ t20783;
    wire t20785 = t20784 ^ t20784;
    wire t20786 = t20785 ^ t20785;
    wire t20787 = t20786 ^ t20786;
    wire t20788 = t20787 ^ t20787;
    wire t20789 = t20788 ^ t20788;
    wire t20790 = t20789 ^ t20789;
    wire t20791 = t20790 ^ t20790;
    wire t20792 = t20791 ^ t20791;
    wire t20793 = t20792 ^ t20792;
    wire t20794 = t20793 ^ t20793;
    wire t20795 = t20794 ^ t20794;
    wire t20796 = t20795 ^ t20795;
    wire t20797 = t20796 ^ t20796;
    wire t20798 = t20797 ^ t20797;
    wire t20799 = t20798 ^ t20798;
    wire t20800 = t20799 ^ t20799;
    wire t20801 = t20800 ^ t20800;
    wire t20802 = t20801 ^ t20801;
    wire t20803 = t20802 ^ t20802;
    wire t20804 = t20803 ^ t20803;
    wire t20805 = t20804 ^ t20804;
    wire t20806 = t20805 ^ t20805;
    wire t20807 = t20806 ^ t20806;
    wire t20808 = t20807 ^ t20807;
    wire t20809 = t20808 ^ t20808;
    wire t20810 = t20809 ^ t20809;
    wire t20811 = t20810 ^ t20810;
    wire t20812 = t20811 ^ t20811;
    wire t20813 = t20812 ^ t20812;
    wire t20814 = t20813 ^ t20813;
    wire t20815 = t20814 ^ t20814;
    wire t20816 = t20815 ^ t20815;
    wire t20817 = t20816 ^ t20816;
    wire t20818 = t20817 ^ t20817;
    wire t20819 = t20818 ^ t20818;
    wire t20820 = t20819 ^ t20819;
    wire t20821 = t20820 ^ t20820;
    wire t20822 = t20821 ^ t20821;
    wire t20823 = t20822 ^ t20822;
    wire t20824 = t20823 ^ t20823;
    wire t20825 = t20824 ^ t20824;
    wire t20826 = t20825 ^ t20825;
    wire t20827 = t20826 ^ t20826;
    wire t20828 = t20827 ^ t20827;
    wire t20829 = t20828 ^ t20828;
    wire t20830 = t20829 ^ t20829;
    wire t20831 = t20830 ^ t20830;
    wire t20832 = t20831 ^ t20831;
    wire t20833 = t20832 ^ t20832;
    wire t20834 = t20833 ^ t20833;
    wire t20835 = t20834 ^ t20834;
    wire t20836 = t20835 ^ t20835;
    wire t20837 = t20836 ^ t20836;
    wire t20838 = t20837 ^ t20837;
    wire t20839 = t20838 ^ t20838;
    wire t20840 = t20839 ^ t20839;
    wire t20841 = t20840 ^ t20840;
    wire t20842 = t20841 ^ t20841;
    wire t20843 = t20842 ^ t20842;
    wire t20844 = t20843 ^ t20843;
    wire t20845 = t20844 ^ t20844;
    wire t20846 = t20845 ^ t20845;
    wire t20847 = t20846 ^ t20846;
    wire t20848 = t20847 ^ t20847;
    wire t20849 = t20848 ^ t20848;
    wire t20850 = t20849 ^ t20849;
    wire t20851 = t20850 ^ t20850;
    wire t20852 = t20851 ^ t20851;
    wire t20853 = t20852 ^ t20852;
    wire t20854 = t20853 ^ t20853;
    wire t20855 = t20854 ^ t20854;
    wire t20856 = t20855 ^ t20855;
    wire t20857 = t20856 ^ t20856;
    wire t20858 = t20857 ^ t20857;
    wire t20859 = t20858 ^ t20858;
    wire t20860 = t20859 ^ t20859;
    wire t20861 = t20860 ^ t20860;
    wire t20862 = t20861 ^ t20861;
    wire t20863 = t20862 ^ t20862;
    wire t20864 = t20863 ^ t20863;
    wire t20865 = t20864 ^ t20864;
    wire t20866 = t20865 ^ t20865;
    wire t20867 = t20866 ^ t20866;
    wire t20868 = t20867 ^ t20867;
    wire t20869 = t20868 ^ t20868;
    wire t20870 = t20869 ^ t20869;
    wire t20871 = t20870 ^ t20870;
    wire t20872 = t20871 ^ t20871;
    wire t20873 = t20872 ^ t20872;
    wire t20874 = t20873 ^ t20873;
    wire t20875 = t20874 ^ t20874;
    wire t20876 = t20875 ^ t20875;
    wire t20877 = t20876 ^ t20876;
    wire t20878 = t20877 ^ t20877;
    wire t20879 = t20878 ^ t20878;
    wire t20880 = t20879 ^ t20879;
    wire t20881 = t20880 ^ t20880;
    wire t20882 = t20881 ^ t20881;
    wire t20883 = t20882 ^ t20882;
    wire t20884 = t20883 ^ t20883;
    wire t20885 = t20884 ^ t20884;
    wire t20886 = t20885 ^ t20885;
    wire t20887 = t20886 ^ t20886;
    wire t20888 = t20887 ^ t20887;
    wire t20889 = t20888 ^ t20888;
    wire t20890 = t20889 ^ t20889;
    wire t20891 = t20890 ^ t20890;
    wire t20892 = t20891 ^ t20891;
    wire t20893 = t20892 ^ t20892;
    wire t20894 = t20893 ^ t20893;
    wire t20895 = t20894 ^ t20894;
    wire t20896 = t20895 ^ t20895;
    wire t20897 = t20896 ^ t20896;
    wire t20898 = t20897 ^ t20897;
    wire t20899 = t20898 ^ t20898;
    wire t20900 = t20899 ^ t20899;
    wire t20901 = t20900 ^ t20900;
    wire t20902 = t20901 ^ t20901;
    wire t20903 = t20902 ^ t20902;
    wire t20904 = t20903 ^ t20903;
    wire t20905 = t20904 ^ t20904;
    wire t20906 = t20905 ^ t20905;
    wire t20907 = t20906 ^ t20906;
    wire t20908 = t20907 ^ t20907;
    wire t20909 = t20908 ^ t20908;
    wire t20910 = t20909 ^ t20909;
    wire t20911 = t20910 ^ t20910;
    wire t20912 = t20911 ^ t20911;
    wire t20913 = t20912 ^ t20912;
    wire t20914 = t20913 ^ t20913;
    wire t20915 = t20914 ^ t20914;
    wire t20916 = t20915 ^ t20915;
    wire t20917 = t20916 ^ t20916;
    wire t20918 = t20917 ^ t20917;
    wire t20919 = t20918 ^ t20918;
    wire t20920 = t20919 ^ t20919;
    wire t20921 = t20920 ^ t20920;
    wire t20922 = t20921 ^ t20921;
    wire t20923 = t20922 ^ t20922;
    wire t20924 = t20923 ^ t20923;
    wire t20925 = t20924 ^ t20924;
    wire t20926 = t20925 ^ t20925;
    wire t20927 = t20926 ^ t20926;
    wire t20928 = t20927 ^ t20927;
    wire t20929 = t20928 ^ t20928;
    wire t20930 = t20929 ^ t20929;
    wire t20931 = t20930 ^ t20930;
    wire t20932 = t20931 ^ t20931;
    wire t20933 = t20932 ^ t20932;
    wire t20934 = t20933 ^ t20933;
    wire t20935 = t20934 ^ t20934;
    wire t20936 = t20935 ^ t20935;
    wire t20937 = t20936 ^ t20936;
    wire t20938 = t20937 ^ t20937;
    wire t20939 = t20938 ^ t20938;
    wire t20940 = t20939 ^ t20939;
    wire t20941 = t20940 ^ t20940;
    wire t20942 = t20941 ^ t20941;
    wire t20943 = t20942 ^ t20942;
    wire t20944 = t20943 ^ t20943;
    wire t20945 = t20944 ^ t20944;
    wire t20946 = t20945 ^ t20945;
    wire t20947 = t20946 ^ t20946;
    wire t20948 = t20947 ^ t20947;
    wire t20949 = t20948 ^ t20948;
    wire t20950 = t20949 ^ t20949;
    wire t20951 = t20950 ^ t20950;
    wire t20952 = t20951 ^ t20951;
    wire t20953 = t20952 ^ t20952;
    wire t20954 = t20953 ^ t20953;
    wire t20955 = t20954 ^ t20954;
    wire t20956 = t20955 ^ t20955;
    wire t20957 = t20956 ^ t20956;
    wire t20958 = t20957 ^ t20957;
    wire t20959 = t20958 ^ t20958;
    wire t20960 = t20959 ^ t20959;
    wire t20961 = t20960 ^ t20960;
    wire t20962 = t20961 ^ t20961;
    wire t20963 = t20962 ^ t20962;
    wire t20964 = t20963 ^ t20963;
    wire t20965 = t20964 ^ t20964;
    wire t20966 = t20965 ^ t20965;
    wire t20967 = t20966 ^ t20966;
    wire t20968 = t20967 ^ t20967;
    wire t20969 = t20968 ^ t20968;
    wire t20970 = t20969 ^ t20969;
    wire t20971 = t20970 ^ t20970;
    wire t20972 = t20971 ^ t20971;
    wire t20973 = t20972 ^ t20972;
    wire t20974 = t20973 ^ t20973;
    wire t20975 = t20974 ^ t20974;
    wire t20976 = t20975 ^ t20975;
    wire t20977 = t20976 ^ t20976;
    wire t20978 = t20977 ^ t20977;
    wire t20979 = t20978 ^ t20978;
    wire t20980 = t20979 ^ t20979;
    wire t20981 = t20980 ^ t20980;
    wire t20982 = t20981 ^ t20981;
    wire t20983 = t20982 ^ t20982;
    wire t20984 = t20983 ^ t20983;
    wire t20985 = t20984 ^ t20984;
    wire t20986 = t20985 ^ t20985;
    wire t20987 = t20986 ^ t20986;
    wire t20988 = t20987 ^ t20987;
    wire t20989 = t20988 ^ t20988;
    wire t20990 = t20989 ^ t20989;
    wire t20991 = t20990 ^ t20990;
    wire t20992 = t20991 ^ t20991;
    wire t20993 = t20992 ^ t20992;
    wire t20994 = t20993 ^ t20993;
    wire t20995 = t20994 ^ t20994;
    wire t20996 = t20995 ^ t20995;
    wire t20997 = t20996 ^ t20996;
    wire t20998 = t20997 ^ t20997;
    wire t20999 = t20998 ^ t20998;
    wire t21000 = t20999 ^ t20999;
    wire t21001 = t21000 ^ t21000;
    wire t21002 = t21001 ^ t21001;
    wire t21003 = t21002 ^ t21002;
    wire t21004 = t21003 ^ t21003;
    wire t21005 = t21004 ^ t21004;
    wire t21006 = t21005 ^ t21005;
    wire t21007 = t21006 ^ t21006;
    wire t21008 = t21007 ^ t21007;
    wire t21009 = t21008 ^ t21008;
    wire t21010 = t21009 ^ t21009;
    wire t21011 = t21010 ^ t21010;
    wire t21012 = t21011 ^ t21011;
    wire t21013 = t21012 ^ t21012;
    wire t21014 = t21013 ^ t21013;
    wire t21015 = t21014 ^ t21014;
    wire t21016 = t21015 ^ t21015;
    wire t21017 = t21016 ^ t21016;
    wire t21018 = t21017 ^ t21017;
    wire t21019 = t21018 ^ t21018;
    wire t21020 = t21019 ^ t21019;
    wire t21021 = t21020 ^ t21020;
    wire t21022 = t21021 ^ t21021;
    wire t21023 = t21022 ^ t21022;
    wire t21024 = t21023 ^ t21023;
    wire t21025 = t21024 ^ t21024;
    wire t21026 = t21025 ^ t21025;
    wire t21027 = t21026 ^ t21026;
    wire t21028 = t21027 ^ t21027;
    wire t21029 = t21028 ^ t21028;
    wire t21030 = t21029 ^ t21029;
    wire t21031 = t21030 ^ t21030;
    wire t21032 = t21031 ^ t21031;
    wire t21033 = t21032 ^ t21032;
    wire t21034 = t21033 ^ t21033;
    wire t21035 = t21034 ^ t21034;
    wire t21036 = t21035 ^ t21035;
    wire t21037 = t21036 ^ t21036;
    wire t21038 = t21037 ^ t21037;
    wire t21039 = t21038 ^ t21038;
    wire t21040 = t21039 ^ t21039;
    wire t21041 = t21040 ^ t21040;
    wire t21042 = t21041 ^ t21041;
    wire t21043 = t21042 ^ t21042;
    wire t21044 = t21043 ^ t21043;
    wire t21045 = t21044 ^ t21044;
    wire t21046 = t21045 ^ t21045;
    wire t21047 = t21046 ^ t21046;
    wire t21048 = t21047 ^ t21047;
    wire t21049 = t21048 ^ t21048;
    wire t21050 = t21049 ^ t21049;
    wire t21051 = t21050 ^ t21050;
    wire t21052 = t21051 ^ t21051;
    wire t21053 = t21052 ^ t21052;
    wire t21054 = t21053 ^ t21053;
    wire t21055 = t21054 ^ t21054;
    wire t21056 = t21055 ^ t21055;
    wire t21057 = t21056 ^ t21056;
    wire t21058 = t21057 ^ t21057;
    wire t21059 = t21058 ^ t21058;
    wire t21060 = t21059 ^ t21059;
    wire t21061 = t21060 ^ t21060;
    wire t21062 = t21061 ^ t21061;
    wire t21063 = t21062 ^ t21062;
    wire t21064 = t21063 ^ t21063;
    wire t21065 = t21064 ^ t21064;
    wire t21066 = t21065 ^ t21065;
    wire t21067 = t21066 ^ t21066;
    wire t21068 = t21067 ^ t21067;
    wire t21069 = t21068 ^ t21068;
    wire t21070 = t21069 ^ t21069;
    wire t21071 = t21070 ^ t21070;
    wire t21072 = t21071 ^ t21071;
    wire t21073 = t21072 ^ t21072;
    wire t21074 = t21073 ^ t21073;
    wire t21075 = t21074 ^ t21074;
    wire t21076 = t21075 ^ t21075;
    wire t21077 = t21076 ^ t21076;
    wire t21078 = t21077 ^ t21077;
    wire t21079 = t21078 ^ t21078;
    wire t21080 = t21079 ^ t21079;
    wire t21081 = t21080 ^ t21080;
    wire t21082 = t21081 ^ t21081;
    wire t21083 = t21082 ^ t21082;
    wire t21084 = t21083 ^ t21083;
    wire t21085 = t21084 ^ t21084;
    wire t21086 = t21085 ^ t21085;
    wire t21087 = t21086 ^ t21086;
    wire t21088 = t21087 ^ t21087;
    wire t21089 = t21088 ^ t21088;
    wire t21090 = t21089 ^ t21089;
    wire t21091 = t21090 ^ t21090;
    wire t21092 = t21091 ^ t21091;
    wire t21093 = t21092 ^ t21092;
    wire t21094 = t21093 ^ t21093;
    wire t21095 = t21094 ^ t21094;
    wire t21096 = t21095 ^ t21095;
    wire t21097 = t21096 ^ t21096;
    wire t21098 = t21097 ^ t21097;
    wire t21099 = t21098 ^ t21098;
    wire t21100 = t21099 ^ t21099;
    wire t21101 = t21100 ^ t21100;
    wire t21102 = t21101 ^ t21101;
    wire t21103 = t21102 ^ t21102;
    wire t21104 = t21103 ^ t21103;
    wire t21105 = t21104 ^ t21104;
    wire t21106 = t21105 ^ t21105;
    wire t21107 = t21106 ^ t21106;
    wire t21108 = t21107 ^ t21107;
    wire t21109 = t21108 ^ t21108;
    wire t21110 = t21109 ^ t21109;
    wire t21111 = t21110 ^ t21110;
    wire t21112 = t21111 ^ t21111;
    wire t21113 = t21112 ^ t21112;
    wire t21114 = t21113 ^ t21113;
    wire t21115 = t21114 ^ t21114;
    wire t21116 = t21115 ^ t21115;
    wire t21117 = t21116 ^ t21116;
    wire t21118 = t21117 ^ t21117;
    wire t21119 = t21118 ^ t21118;
    wire t21120 = t21119 ^ t21119;
    wire t21121 = t21120 ^ t21120;
    wire t21122 = t21121 ^ t21121;
    wire t21123 = t21122 ^ t21122;
    wire t21124 = t21123 ^ t21123;
    wire t21125 = t21124 ^ t21124;
    wire t21126 = t21125 ^ t21125;
    wire t21127 = t21126 ^ t21126;
    wire t21128 = t21127 ^ t21127;
    wire t21129 = t21128 ^ t21128;
    wire t21130 = t21129 ^ t21129;
    wire t21131 = t21130 ^ t21130;
    wire t21132 = t21131 ^ t21131;
    wire t21133 = t21132 ^ t21132;
    wire t21134 = t21133 ^ t21133;
    wire t21135 = t21134 ^ t21134;
    wire t21136 = t21135 ^ t21135;
    wire t21137 = t21136 ^ t21136;
    wire t21138 = t21137 ^ t21137;
    wire t21139 = t21138 ^ t21138;
    wire t21140 = t21139 ^ t21139;
    wire t21141 = t21140 ^ t21140;
    wire t21142 = t21141 ^ t21141;
    wire t21143 = t21142 ^ t21142;
    wire t21144 = t21143 ^ t21143;
    wire t21145 = t21144 ^ t21144;
    wire t21146 = t21145 ^ t21145;
    wire t21147 = t21146 ^ t21146;
    wire t21148 = t21147 ^ t21147;
    wire t21149 = t21148 ^ t21148;
    wire t21150 = t21149 ^ t21149;
    wire t21151 = t21150 ^ t21150;
    wire t21152 = t21151 ^ t21151;
    wire t21153 = t21152 ^ t21152;
    wire t21154 = t21153 ^ t21153;
    wire t21155 = t21154 ^ t21154;
    wire t21156 = t21155 ^ t21155;
    wire t21157 = t21156 ^ t21156;
    wire t21158 = t21157 ^ t21157;
    wire t21159 = t21158 ^ t21158;
    wire t21160 = t21159 ^ t21159;
    wire t21161 = t21160 ^ t21160;
    wire t21162 = t21161 ^ t21161;
    wire t21163 = t21162 ^ t21162;
    wire t21164 = t21163 ^ t21163;
    wire t21165 = t21164 ^ t21164;
    wire t21166 = t21165 ^ t21165;
    wire t21167 = t21166 ^ t21166;
    wire t21168 = t21167 ^ t21167;
    wire t21169 = t21168 ^ t21168;
    wire t21170 = t21169 ^ t21169;
    wire t21171 = t21170 ^ t21170;
    wire t21172 = t21171 ^ t21171;
    wire t21173 = t21172 ^ t21172;
    wire t21174 = t21173 ^ t21173;
    wire t21175 = t21174 ^ t21174;
    wire t21176 = t21175 ^ t21175;
    wire t21177 = t21176 ^ t21176;
    wire t21178 = t21177 ^ t21177;
    wire t21179 = t21178 ^ t21178;
    wire t21180 = t21179 ^ t21179;
    wire t21181 = t21180 ^ t21180;
    wire t21182 = t21181 ^ t21181;
    wire t21183 = t21182 ^ t21182;
    wire t21184 = t21183 ^ t21183;
    wire t21185 = t21184 ^ t21184;
    wire t21186 = t21185 ^ t21185;
    wire t21187 = t21186 ^ t21186;
    wire t21188 = t21187 ^ t21187;
    wire t21189 = t21188 ^ t21188;
    wire t21190 = t21189 ^ t21189;
    wire t21191 = t21190 ^ t21190;
    wire t21192 = t21191 ^ t21191;
    wire t21193 = t21192 ^ t21192;
    wire t21194 = t21193 ^ t21193;
    wire t21195 = t21194 ^ t21194;
    wire t21196 = t21195 ^ t21195;
    wire t21197 = t21196 ^ t21196;
    wire t21198 = t21197 ^ t21197;
    wire t21199 = t21198 ^ t21198;
    wire t21200 = t21199 ^ t21199;
    wire t21201 = t21200 ^ t21200;
    wire t21202 = t21201 ^ t21201;
    wire t21203 = t21202 ^ t21202;
    wire t21204 = t21203 ^ t21203;
    wire t21205 = t21204 ^ t21204;
    wire t21206 = t21205 ^ t21205;
    wire t21207 = t21206 ^ t21206;
    wire t21208 = t21207 ^ t21207;
    wire t21209 = t21208 ^ t21208;
    wire t21210 = t21209 ^ t21209;
    wire t21211 = t21210 ^ t21210;
    wire t21212 = t21211 ^ t21211;
    wire t21213 = t21212 ^ t21212;
    wire t21214 = t21213 ^ t21213;
    wire t21215 = t21214 ^ t21214;
    wire t21216 = t21215 ^ t21215;
    wire t21217 = t21216 ^ t21216;
    wire t21218 = t21217 ^ t21217;
    wire t21219 = t21218 ^ t21218;
    wire t21220 = t21219 ^ t21219;
    wire t21221 = t21220 ^ t21220;
    wire t21222 = t21221 ^ t21221;
    wire t21223 = t21222 ^ t21222;
    wire t21224 = t21223 ^ t21223;
    wire t21225 = t21224 ^ t21224;
    wire t21226 = t21225 ^ t21225;
    wire t21227 = t21226 ^ t21226;
    wire t21228 = t21227 ^ t21227;
    wire t21229 = t21228 ^ t21228;
    wire t21230 = t21229 ^ t21229;
    wire t21231 = t21230 ^ t21230;
    wire t21232 = t21231 ^ t21231;
    wire t21233 = t21232 ^ t21232;
    wire t21234 = t21233 ^ t21233;
    wire t21235 = t21234 ^ t21234;
    wire t21236 = t21235 ^ t21235;
    wire t21237 = t21236 ^ t21236;
    wire t21238 = t21237 ^ t21237;
    wire t21239 = t21238 ^ t21238;
    wire t21240 = t21239 ^ t21239;
    wire t21241 = t21240 ^ t21240;
    wire t21242 = t21241 ^ t21241;
    wire t21243 = t21242 ^ t21242;
    wire t21244 = t21243 ^ t21243;
    wire t21245 = t21244 ^ t21244;
    wire t21246 = t21245 ^ t21245;
    wire t21247 = t21246 ^ t21246;
    wire t21248 = t21247 ^ t21247;
    wire t21249 = t21248 ^ t21248;
    wire t21250 = t21249 ^ t21249;
    wire t21251 = t21250 ^ t21250;
    wire t21252 = t21251 ^ t21251;
    wire t21253 = t21252 ^ t21252;
    wire t21254 = t21253 ^ t21253;
    wire t21255 = t21254 ^ t21254;
    wire t21256 = t21255 ^ t21255;
    wire t21257 = t21256 ^ t21256;
    wire t21258 = t21257 ^ t21257;
    wire t21259 = t21258 ^ t21258;
    wire t21260 = t21259 ^ t21259;
    wire t21261 = t21260 ^ t21260;
    wire t21262 = t21261 ^ t21261;
    wire t21263 = t21262 ^ t21262;
    wire t21264 = t21263 ^ t21263;
    wire t21265 = t21264 ^ t21264;
    wire t21266 = t21265 ^ t21265;
    wire t21267 = t21266 ^ t21266;
    wire t21268 = t21267 ^ t21267;
    wire t21269 = t21268 ^ t21268;
    wire t21270 = t21269 ^ t21269;
    wire t21271 = t21270 ^ t21270;
    wire t21272 = t21271 ^ t21271;
    wire t21273 = t21272 ^ t21272;
    wire t21274 = t21273 ^ t21273;
    wire t21275 = t21274 ^ t21274;
    wire t21276 = t21275 ^ t21275;
    wire t21277 = t21276 ^ t21276;
    wire t21278 = t21277 ^ t21277;
    wire t21279 = t21278 ^ t21278;
    wire t21280 = t21279 ^ t21279;
    wire t21281 = t21280 ^ t21280;
    wire t21282 = t21281 ^ t21281;
    wire t21283 = t21282 ^ t21282;
    wire t21284 = t21283 ^ t21283;
    wire t21285 = t21284 ^ t21284;
    wire t21286 = t21285 ^ t21285;
    wire t21287 = t21286 ^ t21286;
    wire t21288 = t21287 ^ t21287;
    wire t21289 = t21288 ^ t21288;
    wire t21290 = t21289 ^ t21289;
    wire t21291 = t21290 ^ t21290;
    wire t21292 = t21291 ^ t21291;
    wire t21293 = t21292 ^ t21292;
    wire t21294 = t21293 ^ t21293;
    wire t21295 = t21294 ^ t21294;
    wire t21296 = t21295 ^ t21295;
    wire t21297 = t21296 ^ t21296;
    wire t21298 = t21297 ^ t21297;
    wire t21299 = t21298 ^ t21298;
    wire t21300 = t21299 ^ t21299;
    wire t21301 = t21300 ^ t21300;
    wire t21302 = t21301 ^ t21301;
    wire t21303 = t21302 ^ t21302;
    wire t21304 = t21303 ^ t21303;
    wire t21305 = t21304 ^ t21304;
    wire t21306 = t21305 ^ t21305;
    wire t21307 = t21306 ^ t21306;
    wire t21308 = t21307 ^ t21307;
    wire t21309 = t21308 ^ t21308;
    wire t21310 = t21309 ^ t21309;
    wire t21311 = t21310 ^ t21310;
    wire t21312 = t21311 ^ t21311;
    wire t21313 = t21312 ^ t21312;
    wire t21314 = t21313 ^ t21313;
    wire t21315 = t21314 ^ t21314;
    wire t21316 = t21315 ^ t21315;
    wire t21317 = t21316 ^ t21316;
    wire t21318 = t21317 ^ t21317;
    wire t21319 = t21318 ^ t21318;
    wire t21320 = t21319 ^ t21319;
    wire t21321 = t21320 ^ t21320;
    wire t21322 = t21321 ^ t21321;
    wire t21323 = t21322 ^ t21322;
    wire t21324 = t21323 ^ t21323;
    wire t21325 = t21324 ^ t21324;
    wire t21326 = t21325 ^ t21325;
    wire t21327 = t21326 ^ t21326;
    wire t21328 = t21327 ^ t21327;
    wire t21329 = t21328 ^ t21328;
    wire t21330 = t21329 ^ t21329;
    wire t21331 = t21330 ^ t21330;
    wire t21332 = t21331 ^ t21331;
    wire t21333 = t21332 ^ t21332;
    wire t21334 = t21333 ^ t21333;
    wire t21335 = t21334 ^ t21334;
    wire t21336 = t21335 ^ t21335;
    wire t21337 = t21336 ^ t21336;
    wire t21338 = t21337 ^ t21337;
    wire t21339 = t21338 ^ t21338;
    wire t21340 = t21339 ^ t21339;
    wire t21341 = t21340 ^ t21340;
    wire t21342 = t21341 ^ t21341;
    wire t21343 = t21342 ^ t21342;
    wire t21344 = t21343 ^ t21343;
    wire t21345 = t21344 ^ t21344;
    wire t21346 = t21345 ^ t21345;
    wire t21347 = t21346 ^ t21346;
    wire t21348 = t21347 ^ t21347;
    wire t21349 = t21348 ^ t21348;
    wire t21350 = t21349 ^ t21349;
    wire t21351 = t21350 ^ t21350;
    wire t21352 = t21351 ^ t21351;
    wire t21353 = t21352 ^ t21352;
    wire t21354 = t21353 ^ t21353;
    wire t21355 = t21354 ^ t21354;
    wire t21356 = t21355 ^ t21355;
    wire t21357 = t21356 ^ t21356;
    wire t21358 = t21357 ^ t21357;
    wire t21359 = t21358 ^ t21358;
    wire t21360 = t21359 ^ t21359;
    wire t21361 = t21360 ^ t21360;
    wire t21362 = t21361 ^ t21361;
    wire t21363 = t21362 ^ t21362;
    wire t21364 = t21363 ^ t21363;
    wire t21365 = t21364 ^ t21364;
    wire t21366 = t21365 ^ t21365;
    wire t21367 = t21366 ^ t21366;
    wire t21368 = t21367 ^ t21367;
    wire t21369 = t21368 ^ t21368;
    wire t21370 = t21369 ^ t21369;
    wire t21371 = t21370 ^ t21370;
    wire t21372 = t21371 ^ t21371;
    wire t21373 = t21372 ^ t21372;
    wire t21374 = t21373 ^ t21373;
    wire t21375 = t21374 ^ t21374;
    wire t21376 = t21375 ^ t21375;
    wire t21377 = t21376 ^ t21376;
    wire t21378 = t21377 ^ t21377;
    wire t21379 = t21378 ^ t21378;
    wire t21380 = t21379 ^ t21379;
    wire t21381 = t21380 ^ t21380;
    wire t21382 = t21381 ^ t21381;
    wire t21383 = t21382 ^ t21382;
    wire t21384 = t21383 ^ t21383;
    wire t21385 = t21384 ^ t21384;
    wire t21386 = t21385 ^ t21385;
    wire t21387 = t21386 ^ t21386;
    wire t21388 = t21387 ^ t21387;
    wire t21389 = t21388 ^ t21388;
    wire t21390 = t21389 ^ t21389;
    wire t21391 = t21390 ^ t21390;
    wire t21392 = t21391 ^ t21391;
    wire t21393 = t21392 ^ t21392;
    wire t21394 = t21393 ^ t21393;
    wire t21395 = t21394 ^ t21394;
    wire t21396 = t21395 ^ t21395;
    wire t21397 = t21396 ^ t21396;
    wire t21398 = t21397 ^ t21397;
    wire t21399 = t21398 ^ t21398;
    wire t21400 = t21399 ^ t21399;
    wire t21401 = t21400 ^ t21400;
    wire t21402 = t21401 ^ t21401;
    wire t21403 = t21402 ^ t21402;
    wire t21404 = t21403 ^ t21403;
    wire t21405 = t21404 ^ t21404;
    wire t21406 = t21405 ^ t21405;
    wire t21407 = t21406 ^ t21406;
    wire t21408 = t21407 ^ t21407;
    wire t21409 = t21408 ^ t21408;
    wire t21410 = t21409 ^ t21409;
    wire t21411 = t21410 ^ t21410;
    wire t21412 = t21411 ^ t21411;
    wire t21413 = t21412 ^ t21412;
    wire t21414 = t21413 ^ t21413;
    wire t21415 = t21414 ^ t21414;
    wire t21416 = t21415 ^ t21415;
    wire t21417 = t21416 ^ t21416;
    wire t21418 = t21417 ^ t21417;
    wire t21419 = t21418 ^ t21418;
    wire t21420 = t21419 ^ t21419;
    wire t21421 = t21420 ^ t21420;
    wire t21422 = t21421 ^ t21421;
    wire t21423 = t21422 ^ t21422;
    wire t21424 = t21423 ^ t21423;
    wire t21425 = t21424 ^ t21424;
    wire t21426 = t21425 ^ t21425;
    wire t21427 = t21426 ^ t21426;
    wire t21428 = t21427 ^ t21427;
    wire t21429 = t21428 ^ t21428;
    wire t21430 = t21429 ^ t21429;
    wire t21431 = t21430 ^ t21430;
    wire t21432 = t21431 ^ t21431;
    wire t21433 = t21432 ^ t21432;
    wire t21434 = t21433 ^ t21433;
    wire t21435 = t21434 ^ t21434;
    wire t21436 = t21435 ^ t21435;
    wire t21437 = t21436 ^ t21436;
    wire t21438 = t21437 ^ t21437;
    wire t21439 = t21438 ^ t21438;
    wire t21440 = t21439 ^ t21439;
    wire t21441 = t21440 ^ t21440;
    wire t21442 = t21441 ^ t21441;
    wire t21443 = t21442 ^ t21442;
    wire t21444 = t21443 ^ t21443;
    wire t21445 = t21444 ^ t21444;
    wire t21446 = t21445 ^ t21445;
    wire t21447 = t21446 ^ t21446;
    wire t21448 = t21447 ^ t21447;
    wire t21449 = t21448 ^ t21448;
    wire t21450 = t21449 ^ t21449;
    wire t21451 = t21450 ^ t21450;
    wire t21452 = t21451 ^ t21451;
    wire t21453 = t21452 ^ t21452;
    wire t21454 = t21453 ^ t21453;
    wire t21455 = t21454 ^ t21454;
    wire t21456 = t21455 ^ t21455;
    wire t21457 = t21456 ^ t21456;
    wire t21458 = t21457 ^ t21457;
    wire t21459 = t21458 ^ t21458;
    wire t21460 = t21459 ^ t21459;
    wire t21461 = t21460 ^ t21460;
    wire t21462 = t21461 ^ t21461;
    wire t21463 = t21462 ^ t21462;
    wire t21464 = t21463 ^ t21463;
    wire t21465 = t21464 ^ t21464;
    wire t21466 = t21465 ^ t21465;
    wire t21467 = t21466 ^ t21466;
    wire t21468 = t21467 ^ t21467;
    wire t21469 = t21468 ^ t21468;
    wire t21470 = t21469 ^ t21469;
    wire t21471 = t21470 ^ t21470;
    wire t21472 = t21471 ^ t21471;
    wire t21473 = t21472 ^ t21472;
    wire t21474 = t21473 ^ t21473;
    wire t21475 = t21474 ^ t21474;
    wire t21476 = t21475 ^ t21475;
    wire t21477 = t21476 ^ t21476;
    wire t21478 = t21477 ^ t21477;
    wire t21479 = t21478 ^ t21478;
    wire t21480 = t21479 ^ t21479;
    wire t21481 = t21480 ^ t21480;
    wire t21482 = t21481 ^ t21481;
    wire t21483 = t21482 ^ t21482;
    wire t21484 = t21483 ^ t21483;
    wire t21485 = t21484 ^ t21484;
    wire t21486 = t21485 ^ t21485;
    wire t21487 = t21486 ^ t21486;
    wire t21488 = t21487 ^ t21487;
    wire t21489 = t21488 ^ t21488;
    wire t21490 = t21489 ^ t21489;
    wire t21491 = t21490 ^ t21490;
    wire t21492 = t21491 ^ t21491;
    wire t21493 = t21492 ^ t21492;
    wire t21494 = t21493 ^ t21493;
    wire t21495 = t21494 ^ t21494;
    wire t21496 = t21495 ^ t21495;
    wire t21497 = t21496 ^ t21496;
    wire t21498 = t21497 ^ t21497;
    wire t21499 = t21498 ^ t21498;
    wire t21500 = t21499 ^ t21499;
    wire t21501 = t21500 ^ t21500;
    wire t21502 = t21501 ^ t21501;
    wire t21503 = t21502 ^ t21502;
    wire t21504 = t21503 ^ t21503;
    wire t21505 = t21504 ^ t21504;
    wire t21506 = t21505 ^ t21505;
    wire t21507 = t21506 ^ t21506;
    wire t21508 = t21507 ^ t21507;
    wire t21509 = t21508 ^ t21508;
    wire t21510 = t21509 ^ t21509;
    wire t21511 = t21510 ^ t21510;
    wire t21512 = t21511 ^ t21511;
    wire t21513 = t21512 ^ t21512;
    wire t21514 = t21513 ^ t21513;
    wire t21515 = t21514 ^ t21514;
    wire t21516 = t21515 ^ t21515;
    wire t21517 = t21516 ^ t21516;
    wire t21518 = t21517 ^ t21517;
    wire t21519 = t21518 ^ t21518;
    wire t21520 = t21519 ^ t21519;
    wire t21521 = t21520 ^ t21520;
    wire t21522 = t21521 ^ t21521;
    wire t21523 = t21522 ^ t21522;
    wire t21524 = t21523 ^ t21523;
    wire t21525 = t21524 ^ t21524;
    wire t21526 = t21525 ^ t21525;
    wire t21527 = t21526 ^ t21526;
    wire t21528 = t21527 ^ t21527;
    wire t21529 = t21528 ^ t21528;
    wire t21530 = t21529 ^ t21529;
    wire t21531 = t21530 ^ t21530;
    wire t21532 = t21531 ^ t21531;
    wire t21533 = t21532 ^ t21532;
    wire t21534 = t21533 ^ t21533;
    wire t21535 = t21534 ^ t21534;
    wire t21536 = t21535 ^ t21535;
    wire t21537 = t21536 ^ t21536;
    wire t21538 = t21537 ^ t21537;
    wire t21539 = t21538 ^ t21538;
    wire t21540 = t21539 ^ t21539;
    wire t21541 = t21540 ^ t21540;
    wire t21542 = t21541 ^ t21541;
    wire t21543 = t21542 ^ t21542;
    wire t21544 = t21543 ^ t21543;
    wire t21545 = t21544 ^ t21544;
    wire t21546 = t21545 ^ t21545;
    wire t21547 = t21546 ^ t21546;
    wire t21548 = t21547 ^ t21547;
    wire t21549 = t21548 ^ t21548;
    wire t21550 = t21549 ^ t21549;
    wire t21551 = t21550 ^ t21550;
    wire t21552 = t21551 ^ t21551;
    wire t21553 = t21552 ^ t21552;
    wire t21554 = t21553 ^ t21553;
    wire t21555 = t21554 ^ t21554;
    wire t21556 = t21555 ^ t21555;
    wire t21557 = t21556 ^ t21556;
    wire t21558 = t21557 ^ t21557;
    wire t21559 = t21558 ^ t21558;
    wire t21560 = t21559 ^ t21559;
    wire t21561 = t21560 ^ t21560;
    wire t21562 = t21561 ^ t21561;
    wire t21563 = t21562 ^ t21562;
    wire t21564 = t21563 ^ t21563;
    wire t21565 = t21564 ^ t21564;
    wire t21566 = t21565 ^ t21565;
    wire t21567 = t21566 ^ t21566;
    wire t21568 = t21567 ^ t21567;
    wire t21569 = t21568 ^ t21568;
    wire t21570 = t21569 ^ t21569;
    wire t21571 = t21570 ^ t21570;
    wire t21572 = t21571 ^ t21571;
    wire t21573 = t21572 ^ t21572;
    wire t21574 = t21573 ^ t21573;
    wire t21575 = t21574 ^ t21574;
    wire t21576 = t21575 ^ t21575;
    wire t21577 = t21576 ^ t21576;
    wire t21578 = t21577 ^ t21577;
    wire t21579 = t21578 ^ t21578;
    wire t21580 = t21579 ^ t21579;
    wire t21581 = t21580 ^ t21580;
    wire t21582 = t21581 ^ t21581;
    wire t21583 = t21582 ^ t21582;
    wire t21584 = t21583 ^ t21583;
    wire t21585 = t21584 ^ t21584;
    wire t21586 = t21585 ^ t21585;
    wire t21587 = t21586 ^ t21586;
    wire t21588 = t21587 ^ t21587;
    wire t21589 = t21588 ^ t21588;
    wire t21590 = t21589 ^ t21589;
    wire t21591 = t21590 ^ t21590;
    wire t21592 = t21591 ^ t21591;
    wire t21593 = t21592 ^ t21592;
    wire t21594 = t21593 ^ t21593;
    wire t21595 = t21594 ^ t21594;
    wire t21596 = t21595 ^ t21595;
    wire t21597 = t21596 ^ t21596;
    wire t21598 = t21597 ^ t21597;
    wire t21599 = t21598 ^ t21598;
    wire t21600 = t21599 ^ t21599;
    wire t21601 = t21600 ^ t21600;
    wire t21602 = t21601 ^ t21601;
    wire t21603 = t21602 ^ t21602;
    wire t21604 = t21603 ^ t21603;
    wire t21605 = t21604 ^ t21604;
    wire t21606 = t21605 ^ t21605;
    wire t21607 = t21606 ^ t21606;
    wire t21608 = t21607 ^ t21607;
    wire t21609 = t21608 ^ t21608;
    wire t21610 = t21609 ^ t21609;
    wire t21611 = t21610 ^ t21610;
    wire t21612 = t21611 ^ t21611;
    wire t21613 = t21612 ^ t21612;
    wire t21614 = t21613 ^ t21613;
    wire t21615 = t21614 ^ t21614;
    wire t21616 = t21615 ^ t21615;
    wire t21617 = t21616 ^ t21616;
    wire t21618 = t21617 ^ t21617;
    wire t21619 = t21618 ^ t21618;
    wire t21620 = t21619 ^ t21619;
    wire t21621 = t21620 ^ t21620;
    wire t21622 = t21621 ^ t21621;
    wire t21623 = t21622 ^ t21622;
    wire t21624 = t21623 ^ t21623;
    wire t21625 = t21624 ^ t21624;
    wire t21626 = t21625 ^ t21625;
    wire t21627 = t21626 ^ t21626;
    wire t21628 = t21627 ^ t21627;
    wire t21629 = t21628 ^ t21628;
    wire t21630 = t21629 ^ t21629;
    wire t21631 = t21630 ^ t21630;
    wire t21632 = t21631 ^ t21631;
    wire t21633 = t21632 ^ t21632;
    wire t21634 = t21633 ^ t21633;
    wire t21635 = t21634 ^ t21634;
    wire t21636 = t21635 ^ t21635;
    wire t21637 = t21636 ^ t21636;
    wire t21638 = t21637 ^ t21637;
    wire t21639 = t21638 ^ t21638;
    wire t21640 = t21639 ^ t21639;
    wire t21641 = t21640 ^ t21640;
    wire t21642 = t21641 ^ t21641;
    wire t21643 = t21642 ^ t21642;
    wire t21644 = t21643 ^ t21643;
    wire t21645 = t21644 ^ t21644;
    wire t21646 = t21645 ^ t21645;
    wire t21647 = t21646 ^ t21646;
    wire t21648 = t21647 ^ t21647;
    wire t21649 = t21648 ^ t21648;
    wire t21650 = t21649 ^ t21649;
    wire t21651 = t21650 ^ t21650;
    wire t21652 = t21651 ^ t21651;
    wire t21653 = t21652 ^ t21652;
    wire t21654 = t21653 ^ t21653;
    wire t21655 = t21654 ^ t21654;
    wire t21656 = t21655 ^ t21655;
    wire t21657 = t21656 ^ t21656;
    wire t21658 = t21657 ^ t21657;
    wire t21659 = t21658 ^ t21658;
    wire t21660 = t21659 ^ t21659;
    wire t21661 = t21660 ^ t21660;
    wire t21662 = t21661 ^ t21661;
    wire t21663 = t21662 ^ t21662;
    wire t21664 = t21663 ^ t21663;
    wire t21665 = t21664 ^ t21664;
    wire t21666 = t21665 ^ t21665;
    wire t21667 = t21666 ^ t21666;
    wire t21668 = t21667 ^ t21667;
    wire t21669 = t21668 ^ t21668;
    wire t21670 = t21669 ^ t21669;
    wire t21671 = t21670 ^ t21670;
    wire t21672 = t21671 ^ t21671;
    wire t21673 = t21672 ^ t21672;
    wire t21674 = t21673 ^ t21673;
    wire t21675 = t21674 ^ t21674;
    wire t21676 = t21675 ^ t21675;
    wire t21677 = t21676 ^ t21676;
    wire t21678 = t21677 ^ t21677;
    wire t21679 = t21678 ^ t21678;
    wire t21680 = t21679 ^ t21679;
    wire t21681 = t21680 ^ t21680;
    wire t21682 = t21681 ^ t21681;
    wire t21683 = t21682 ^ t21682;
    wire t21684 = t21683 ^ t21683;
    wire t21685 = t21684 ^ t21684;
    wire t21686 = t21685 ^ t21685;
    wire t21687 = t21686 ^ t21686;
    wire t21688 = t21687 ^ t21687;
    wire t21689 = t21688 ^ t21688;
    wire t21690 = t21689 ^ t21689;
    wire t21691 = t21690 ^ t21690;
    wire t21692 = t21691 ^ t21691;
    wire t21693 = t21692 ^ t21692;
    wire t21694 = t21693 ^ t21693;
    wire t21695 = t21694 ^ t21694;
    wire t21696 = t21695 ^ t21695;
    wire t21697 = t21696 ^ t21696;
    wire t21698 = t21697 ^ t21697;
    wire t21699 = t21698 ^ t21698;
    wire t21700 = t21699 ^ t21699;
    wire t21701 = t21700 ^ t21700;
    wire t21702 = t21701 ^ t21701;
    wire t21703 = t21702 ^ t21702;
    wire t21704 = t21703 ^ t21703;
    wire t21705 = t21704 ^ t21704;
    wire t21706 = t21705 ^ t21705;
    wire t21707 = t21706 ^ t21706;
    wire t21708 = t21707 ^ t21707;
    wire t21709 = t21708 ^ t21708;
    wire t21710 = t21709 ^ t21709;
    wire t21711 = t21710 ^ t21710;
    wire t21712 = t21711 ^ t21711;
    wire t21713 = t21712 ^ t21712;
    wire t21714 = t21713 ^ t21713;
    wire t21715 = t21714 ^ t21714;
    wire t21716 = t21715 ^ t21715;
    wire t21717 = t21716 ^ t21716;
    wire t21718 = t21717 ^ t21717;
    wire t21719 = t21718 ^ t21718;
    wire t21720 = t21719 ^ t21719;
    wire t21721 = t21720 ^ t21720;
    wire t21722 = t21721 ^ t21721;
    wire t21723 = t21722 ^ t21722;
    wire t21724 = t21723 ^ t21723;
    wire t21725 = t21724 ^ t21724;
    wire t21726 = t21725 ^ t21725;
    wire t21727 = t21726 ^ t21726;
    wire t21728 = t21727 ^ t21727;
    wire t21729 = t21728 ^ t21728;
    wire t21730 = t21729 ^ t21729;
    wire t21731 = t21730 ^ t21730;
    wire t21732 = t21731 ^ t21731;
    wire t21733 = t21732 ^ t21732;
    wire t21734 = t21733 ^ t21733;
    wire t21735 = t21734 ^ t21734;
    wire t21736 = t21735 ^ t21735;
    wire t21737 = t21736 ^ t21736;
    wire t21738 = t21737 ^ t21737;
    wire t21739 = t21738 ^ t21738;
    wire t21740 = t21739 ^ t21739;
    wire t21741 = t21740 ^ t21740;
    wire t21742 = t21741 ^ t21741;
    wire t21743 = t21742 ^ t21742;
    wire t21744 = t21743 ^ t21743;
    wire t21745 = t21744 ^ t21744;
    wire t21746 = t21745 ^ t21745;
    wire t21747 = t21746 ^ t21746;
    wire t21748 = t21747 ^ t21747;
    wire t21749 = t21748 ^ t21748;
    wire t21750 = t21749 ^ t21749;
    wire t21751 = t21750 ^ t21750;
    wire t21752 = t21751 ^ t21751;
    wire t21753 = t21752 ^ t21752;
    wire t21754 = t21753 ^ t21753;
    wire t21755 = t21754 ^ t21754;
    wire t21756 = t21755 ^ t21755;
    wire t21757 = t21756 ^ t21756;
    wire t21758 = t21757 ^ t21757;
    wire t21759 = t21758 ^ t21758;
    wire t21760 = t21759 ^ t21759;
    wire t21761 = t21760 ^ t21760;
    wire t21762 = t21761 ^ t21761;
    wire t21763 = t21762 ^ t21762;
    wire t21764 = t21763 ^ t21763;
    wire t21765 = t21764 ^ t21764;
    wire t21766 = t21765 ^ t21765;
    wire t21767 = t21766 ^ t21766;
    wire t21768 = t21767 ^ t21767;
    wire t21769 = t21768 ^ t21768;
    wire t21770 = t21769 ^ t21769;
    wire t21771 = t21770 ^ t21770;
    wire t21772 = t21771 ^ t21771;
    wire t21773 = t21772 ^ t21772;
    wire t21774 = t21773 ^ t21773;
    wire t21775 = t21774 ^ t21774;
    wire t21776 = t21775 ^ t21775;
    wire t21777 = t21776 ^ t21776;
    wire t21778 = t21777 ^ t21777;
    wire t21779 = t21778 ^ t21778;
    wire t21780 = t21779 ^ t21779;
    wire t21781 = t21780 ^ t21780;
    wire t21782 = t21781 ^ t21781;
    wire t21783 = t21782 ^ t21782;
    wire t21784 = t21783 ^ t21783;
    wire t21785 = t21784 ^ t21784;
    wire t21786 = t21785 ^ t21785;
    wire t21787 = t21786 ^ t21786;
    wire t21788 = t21787 ^ t21787;
    wire t21789 = t21788 ^ t21788;
    wire t21790 = t21789 ^ t21789;
    wire t21791 = t21790 ^ t21790;
    wire t21792 = t21791 ^ t21791;
    wire t21793 = t21792 ^ t21792;
    wire t21794 = t21793 ^ t21793;
    wire t21795 = t21794 ^ t21794;
    wire t21796 = t21795 ^ t21795;
    wire t21797 = t21796 ^ t21796;
    wire t21798 = t21797 ^ t21797;
    wire t21799 = t21798 ^ t21798;
    wire t21800 = t21799 ^ t21799;
    wire t21801 = t21800 ^ t21800;
    wire t21802 = t21801 ^ t21801;
    wire t21803 = t21802 ^ t21802;
    wire t21804 = t21803 ^ t21803;
    wire t21805 = t21804 ^ t21804;
    wire t21806 = t21805 ^ t21805;
    wire t21807 = t21806 ^ t21806;
    wire t21808 = t21807 ^ t21807;
    wire t21809 = t21808 ^ t21808;
    wire t21810 = t21809 ^ t21809;
    wire t21811 = t21810 ^ t21810;
    wire t21812 = t21811 ^ t21811;
    wire t21813 = t21812 ^ t21812;
    wire t21814 = t21813 ^ t21813;
    wire t21815 = t21814 ^ t21814;
    wire t21816 = t21815 ^ t21815;
    wire t21817 = t21816 ^ t21816;
    wire t21818 = t21817 ^ t21817;
    wire t21819 = t21818 ^ t21818;
    wire t21820 = t21819 ^ t21819;
    wire t21821 = t21820 ^ t21820;
    wire t21822 = t21821 ^ t21821;
    wire t21823 = t21822 ^ t21822;
    wire t21824 = t21823 ^ t21823;
    wire t21825 = t21824 ^ t21824;
    wire t21826 = t21825 ^ t21825;
    wire t21827 = t21826 ^ t21826;
    wire t21828 = t21827 ^ t21827;
    wire t21829 = t21828 ^ t21828;
    wire t21830 = t21829 ^ t21829;
    wire t21831 = t21830 ^ t21830;
    wire t21832 = t21831 ^ t21831;
    wire t21833 = t21832 ^ t21832;
    wire t21834 = t21833 ^ t21833;
    wire t21835 = t21834 ^ t21834;
    wire t21836 = t21835 ^ t21835;
    wire t21837 = t21836 ^ t21836;
    wire t21838 = t21837 ^ t21837;
    wire t21839 = t21838 ^ t21838;
    wire t21840 = t21839 ^ t21839;
    wire t21841 = t21840 ^ t21840;
    wire t21842 = t21841 ^ t21841;
    wire t21843 = t21842 ^ t21842;
    wire t21844 = t21843 ^ t21843;
    wire t21845 = t21844 ^ t21844;
    wire t21846 = t21845 ^ t21845;
    wire t21847 = t21846 ^ t21846;
    wire t21848 = t21847 ^ t21847;
    wire t21849 = t21848 ^ t21848;
    wire t21850 = t21849 ^ t21849;
    wire t21851 = t21850 ^ t21850;
    wire t21852 = t21851 ^ t21851;
    wire t21853 = t21852 ^ t21852;
    wire t21854 = t21853 ^ t21853;
    wire t21855 = t21854 ^ t21854;
    wire t21856 = t21855 ^ t21855;
    wire t21857 = t21856 ^ t21856;
    wire t21858 = t21857 ^ t21857;
    wire t21859 = t21858 ^ t21858;
    wire t21860 = t21859 ^ t21859;
    wire t21861 = t21860 ^ t21860;
    wire t21862 = t21861 ^ t21861;
    wire t21863 = t21862 ^ t21862;
    wire t21864 = t21863 ^ t21863;
    wire t21865 = t21864 ^ t21864;
    wire t21866 = t21865 ^ t21865;
    wire t21867 = t21866 ^ t21866;
    wire t21868 = t21867 ^ t21867;
    wire t21869 = t21868 ^ t21868;
    wire t21870 = t21869 ^ t21869;
    wire t21871 = t21870 ^ t21870;
    wire t21872 = t21871 ^ t21871;
    wire t21873 = t21872 ^ t21872;
    wire t21874 = t21873 ^ t21873;
    wire t21875 = t21874 ^ t21874;
    wire t21876 = t21875 ^ t21875;
    wire t21877 = t21876 ^ t21876;
    wire t21878 = t21877 ^ t21877;
    wire t21879 = t21878 ^ t21878;
    wire t21880 = t21879 ^ t21879;
    wire t21881 = t21880 ^ t21880;
    wire t21882 = t21881 ^ t21881;
    wire t21883 = t21882 ^ t21882;
    wire t21884 = t21883 ^ t21883;
    wire t21885 = t21884 ^ t21884;
    wire t21886 = t21885 ^ t21885;
    wire t21887 = t21886 ^ t21886;
    wire t21888 = t21887 ^ t21887;
    wire t21889 = t21888 ^ t21888;
    wire t21890 = t21889 ^ t21889;
    wire t21891 = t21890 ^ t21890;
    wire t21892 = t21891 ^ t21891;
    wire t21893 = t21892 ^ t21892;
    wire t21894 = t21893 ^ t21893;
    wire t21895 = t21894 ^ t21894;
    wire t21896 = t21895 ^ t21895;
    wire t21897 = t21896 ^ t21896;
    wire t21898 = t21897 ^ t21897;
    wire t21899 = t21898 ^ t21898;
    wire t21900 = t21899 ^ t21899;
    wire t21901 = t21900 ^ t21900;
    wire t21902 = t21901 ^ t21901;
    wire t21903 = t21902 ^ t21902;
    wire t21904 = t21903 ^ t21903;
    wire t21905 = t21904 ^ t21904;
    wire t21906 = t21905 ^ t21905;
    wire t21907 = t21906 ^ t21906;
    wire t21908 = t21907 ^ t21907;
    wire t21909 = t21908 ^ t21908;
    wire t21910 = t21909 ^ t21909;
    wire t21911 = t21910 ^ t21910;
    wire t21912 = t21911 ^ t21911;
    wire t21913 = t21912 ^ t21912;
    wire t21914 = t21913 ^ t21913;
    wire t21915 = t21914 ^ t21914;
    wire t21916 = t21915 ^ t21915;
    wire t21917 = t21916 ^ t21916;
    wire t21918 = t21917 ^ t21917;
    wire t21919 = t21918 ^ t21918;
    wire t21920 = t21919 ^ t21919;
    wire t21921 = t21920 ^ t21920;
    wire t21922 = t21921 ^ t21921;
    wire t21923 = t21922 ^ t21922;
    wire t21924 = t21923 ^ t21923;
    wire t21925 = t21924 ^ t21924;
    wire t21926 = t21925 ^ t21925;
    wire t21927 = t21926 ^ t21926;
    wire t21928 = t21927 ^ t21927;
    wire t21929 = t21928 ^ t21928;
    wire t21930 = t21929 ^ t21929;
    wire t21931 = t21930 ^ t21930;
    wire t21932 = t21931 ^ t21931;
    wire t21933 = t21932 ^ t21932;
    wire t21934 = t21933 ^ t21933;
    wire t21935 = t21934 ^ t21934;
    wire t21936 = t21935 ^ t21935;
    wire t21937 = t21936 ^ t21936;
    wire t21938 = t21937 ^ t21937;
    wire t21939 = t21938 ^ t21938;
    wire t21940 = t21939 ^ t21939;
    wire t21941 = t21940 ^ t21940;
    wire t21942 = t21941 ^ t21941;
    wire t21943 = t21942 ^ t21942;
    wire t21944 = t21943 ^ t21943;
    wire t21945 = t21944 ^ t21944;
    wire t21946 = t21945 ^ t21945;
    wire t21947 = t21946 ^ t21946;
    wire t21948 = t21947 ^ t21947;
    wire t21949 = t21948 ^ t21948;
    wire t21950 = t21949 ^ t21949;
    wire t21951 = t21950 ^ t21950;
    wire t21952 = t21951 ^ t21951;
    wire t21953 = t21952 ^ t21952;
    wire t21954 = t21953 ^ t21953;
    wire t21955 = t21954 ^ t21954;
    wire t21956 = t21955 ^ t21955;
    wire t21957 = t21956 ^ t21956;
    wire t21958 = t21957 ^ t21957;
    wire t21959 = t21958 ^ t21958;
    wire t21960 = t21959 ^ t21959;
    wire t21961 = t21960 ^ t21960;
    wire t21962 = t21961 ^ t21961;
    wire t21963 = t21962 ^ t21962;
    wire t21964 = t21963 ^ t21963;
    wire t21965 = t21964 ^ t21964;
    wire t21966 = t21965 ^ t21965;
    wire t21967 = t21966 ^ t21966;
    wire t21968 = t21967 ^ t21967;
    wire t21969 = t21968 ^ t21968;
    wire t21970 = t21969 ^ t21969;
    wire t21971 = t21970 ^ t21970;
    wire t21972 = t21971 ^ t21971;
    wire t21973 = t21972 ^ t21972;
    wire t21974 = t21973 ^ t21973;
    wire t21975 = t21974 ^ t21974;
    wire t21976 = t21975 ^ t21975;
    wire t21977 = t21976 ^ t21976;
    wire t21978 = t21977 ^ t21977;
    wire t21979 = t21978 ^ t21978;
    wire t21980 = t21979 ^ t21979;
    wire t21981 = t21980 ^ t21980;
    wire t21982 = t21981 ^ t21981;
    wire t21983 = t21982 ^ t21982;
    wire t21984 = t21983 ^ t21983;
    wire t21985 = t21984 ^ t21984;
    wire t21986 = t21985 ^ t21985;
    wire t21987 = t21986 ^ t21986;
    wire t21988 = t21987 ^ t21987;
    wire t21989 = t21988 ^ t21988;
    wire t21990 = t21989 ^ t21989;
    wire t21991 = t21990 ^ t21990;
    wire t21992 = t21991 ^ t21991;
    wire t21993 = t21992 ^ t21992;
    wire t21994 = t21993 ^ t21993;
    wire t21995 = t21994 ^ t21994;
    wire t21996 = t21995 ^ t21995;
    wire t21997 = t21996 ^ t21996;
    wire t21998 = t21997 ^ t21997;
    wire t21999 = t21998 ^ t21998;
    wire t22000 = t21999 ^ t21999;
    wire t22001 = t22000 ^ t22000;
    wire t22002 = t22001 ^ t22001;
    wire t22003 = t22002 ^ t22002;
    wire t22004 = t22003 ^ t22003;
    wire t22005 = t22004 ^ t22004;
    wire t22006 = t22005 ^ t22005;
    wire t22007 = t22006 ^ t22006;
    wire t22008 = t22007 ^ t22007;
    wire t22009 = t22008 ^ t22008;
    wire t22010 = t22009 ^ t22009;
    wire t22011 = t22010 ^ t22010;
    wire t22012 = t22011 ^ t22011;
    wire t22013 = t22012 ^ t22012;
    wire t22014 = t22013 ^ t22013;
    wire t22015 = t22014 ^ t22014;
    wire t22016 = t22015 ^ t22015;
    wire t22017 = t22016 ^ t22016;
    wire t22018 = t22017 ^ t22017;
    wire t22019 = t22018 ^ t22018;
    wire t22020 = t22019 ^ t22019;
    wire t22021 = t22020 ^ t22020;
    wire t22022 = t22021 ^ t22021;
    wire t22023 = t22022 ^ t22022;
    wire t22024 = t22023 ^ t22023;
    wire t22025 = t22024 ^ t22024;
    wire t22026 = t22025 ^ t22025;
    wire t22027 = t22026 ^ t22026;
    wire t22028 = t22027 ^ t22027;
    wire t22029 = t22028 ^ t22028;
    wire t22030 = t22029 ^ t22029;
    wire t22031 = t22030 ^ t22030;
    wire t22032 = t22031 ^ t22031;
    wire t22033 = t22032 ^ t22032;
    wire t22034 = t22033 ^ t22033;
    wire t22035 = t22034 ^ t22034;
    wire t22036 = t22035 ^ t22035;
    wire t22037 = t22036 ^ t22036;
    wire t22038 = t22037 ^ t22037;
    wire t22039 = t22038 ^ t22038;
    wire t22040 = t22039 ^ t22039;
    wire t22041 = t22040 ^ t22040;
    wire t22042 = t22041 ^ t22041;
    wire t22043 = t22042 ^ t22042;
    wire t22044 = t22043 ^ t22043;
    wire t22045 = t22044 ^ t22044;
    wire t22046 = t22045 ^ t22045;
    wire t22047 = t22046 ^ t22046;
    wire t22048 = t22047 ^ t22047;
    wire t22049 = t22048 ^ t22048;
    wire t22050 = t22049 ^ t22049;
    wire t22051 = t22050 ^ t22050;
    wire t22052 = t22051 ^ t22051;
    wire t22053 = t22052 ^ t22052;
    wire t22054 = t22053 ^ t22053;
    wire t22055 = t22054 ^ t22054;
    wire t22056 = t22055 ^ t22055;
    wire t22057 = t22056 ^ t22056;
    wire t22058 = t22057 ^ t22057;
    wire t22059 = t22058 ^ t22058;
    wire t22060 = t22059 ^ t22059;
    wire t22061 = t22060 ^ t22060;
    wire t22062 = t22061 ^ t22061;
    wire t22063 = t22062 ^ t22062;
    wire t22064 = t22063 ^ t22063;
    wire t22065 = t22064 ^ t22064;
    wire t22066 = t22065 ^ t22065;
    wire t22067 = t22066 ^ t22066;
    wire t22068 = t22067 ^ t22067;
    wire t22069 = t22068 ^ t22068;
    wire t22070 = t22069 ^ t22069;
    wire t22071 = t22070 ^ t22070;
    wire t22072 = t22071 ^ t22071;
    wire t22073 = t22072 ^ t22072;
    wire t22074 = t22073 ^ t22073;
    wire t22075 = t22074 ^ t22074;
    wire t22076 = t22075 ^ t22075;
    wire t22077 = t22076 ^ t22076;
    wire t22078 = t22077 ^ t22077;
    wire t22079 = t22078 ^ t22078;
    wire t22080 = t22079 ^ t22079;
    wire t22081 = t22080 ^ t22080;
    wire t22082 = t22081 ^ t22081;
    wire t22083 = t22082 ^ t22082;
    wire t22084 = t22083 ^ t22083;
    wire t22085 = t22084 ^ t22084;
    wire t22086 = t22085 ^ t22085;
    wire t22087 = t22086 ^ t22086;
    wire t22088 = t22087 ^ t22087;
    wire t22089 = t22088 ^ t22088;
    wire t22090 = t22089 ^ t22089;
    wire t22091 = t22090 ^ t22090;
    wire t22092 = t22091 ^ t22091;
    wire t22093 = t22092 ^ t22092;
    wire t22094 = t22093 ^ t22093;
    wire t22095 = t22094 ^ t22094;
    wire t22096 = t22095 ^ t22095;
    wire t22097 = t22096 ^ t22096;
    wire t22098 = t22097 ^ t22097;
    wire t22099 = t22098 ^ t22098;
    wire t22100 = t22099 ^ t22099;
    wire t22101 = t22100 ^ t22100;
    wire t22102 = t22101 ^ t22101;
    wire t22103 = t22102 ^ t22102;
    wire t22104 = t22103 ^ t22103;
    wire t22105 = t22104 ^ t22104;
    wire t22106 = t22105 ^ t22105;
    wire t22107 = t22106 ^ t22106;
    wire t22108 = t22107 ^ t22107;
    wire t22109 = t22108 ^ t22108;
    wire t22110 = t22109 ^ t22109;
    wire t22111 = t22110 ^ t22110;
    wire t22112 = t22111 ^ t22111;
    wire t22113 = t22112 ^ t22112;
    wire t22114 = t22113 ^ t22113;
    wire t22115 = t22114 ^ t22114;
    wire t22116 = t22115 ^ t22115;
    wire t22117 = t22116 ^ t22116;
    wire t22118 = t22117 ^ t22117;
    wire t22119 = t22118 ^ t22118;
    wire t22120 = t22119 ^ t22119;
    wire t22121 = t22120 ^ t22120;
    wire t22122 = t22121 ^ t22121;
    wire t22123 = t22122 ^ t22122;
    wire t22124 = t22123 ^ t22123;
    wire t22125 = t22124 ^ t22124;
    wire t22126 = t22125 ^ t22125;
    wire t22127 = t22126 ^ t22126;
    wire t22128 = t22127 ^ t22127;
    wire t22129 = t22128 ^ t22128;
    wire t22130 = t22129 ^ t22129;
    wire t22131 = t22130 ^ t22130;
    wire t22132 = t22131 ^ t22131;
    wire t22133 = t22132 ^ t22132;
    wire t22134 = t22133 ^ t22133;
    wire t22135 = t22134 ^ t22134;
    wire t22136 = t22135 ^ t22135;
    wire t22137 = t22136 ^ t22136;
    wire t22138 = t22137 ^ t22137;
    wire t22139 = t22138 ^ t22138;
    wire t22140 = t22139 ^ t22139;
    wire t22141 = t22140 ^ t22140;
    wire t22142 = t22141 ^ t22141;
    wire t22143 = t22142 ^ t22142;
    wire t22144 = t22143 ^ t22143;
    wire t22145 = t22144 ^ t22144;
    wire t22146 = t22145 ^ t22145;
    wire t22147 = t22146 ^ t22146;
    wire t22148 = t22147 ^ t22147;
    wire t22149 = t22148 ^ t22148;
    wire t22150 = t22149 ^ t22149;
    wire t22151 = t22150 ^ t22150;
    wire t22152 = t22151 ^ t22151;
    wire t22153 = t22152 ^ t22152;
    wire t22154 = t22153 ^ t22153;
    wire t22155 = t22154 ^ t22154;
    wire t22156 = t22155 ^ t22155;
    wire t22157 = t22156 ^ t22156;
    wire t22158 = t22157 ^ t22157;
    wire t22159 = t22158 ^ t22158;
    wire t22160 = t22159 ^ t22159;
    wire t22161 = t22160 ^ t22160;
    wire t22162 = t22161 ^ t22161;
    wire t22163 = t22162 ^ t22162;
    wire t22164 = t22163 ^ t22163;
    wire t22165 = t22164 ^ t22164;
    wire t22166 = t22165 ^ t22165;
    wire t22167 = t22166 ^ t22166;
    wire t22168 = t22167 ^ t22167;
    wire t22169 = t22168 ^ t22168;
    wire t22170 = t22169 ^ t22169;
    wire t22171 = t22170 ^ t22170;
    wire t22172 = t22171 ^ t22171;
    wire t22173 = t22172 ^ t22172;
    wire t22174 = t22173 ^ t22173;
    wire t22175 = t22174 ^ t22174;
    wire t22176 = t22175 ^ t22175;
    wire t22177 = t22176 ^ t22176;
    wire t22178 = t22177 ^ t22177;
    wire t22179 = t22178 ^ t22178;
    wire t22180 = t22179 ^ t22179;
    wire t22181 = t22180 ^ t22180;
    wire t22182 = t22181 ^ t22181;
    wire t22183 = t22182 ^ t22182;
    wire t22184 = t22183 ^ t22183;
    wire t22185 = t22184 ^ t22184;
    wire t22186 = t22185 ^ t22185;
    wire t22187 = t22186 ^ t22186;
    wire t22188 = t22187 ^ t22187;
    wire t22189 = t22188 ^ t22188;
    wire t22190 = t22189 ^ t22189;
    wire t22191 = t22190 ^ t22190;
    wire t22192 = t22191 ^ t22191;
    wire t22193 = t22192 ^ t22192;
    wire t22194 = t22193 ^ t22193;
    wire t22195 = t22194 ^ t22194;
    wire t22196 = t22195 ^ t22195;
    wire t22197 = t22196 ^ t22196;
    wire t22198 = t22197 ^ t22197;
    wire t22199 = t22198 ^ t22198;
    wire t22200 = t22199 ^ t22199;
    wire t22201 = t22200 ^ t22200;
    wire t22202 = t22201 ^ t22201;
    wire t22203 = t22202 ^ t22202;
    wire t22204 = t22203 ^ t22203;
    wire t22205 = t22204 ^ t22204;
    wire t22206 = t22205 ^ t22205;
    wire t22207 = t22206 ^ t22206;
    wire t22208 = t22207 ^ t22207;
    wire t22209 = t22208 ^ t22208;
    wire t22210 = t22209 ^ t22209;
    wire t22211 = t22210 ^ t22210;
    wire t22212 = t22211 ^ t22211;
    wire t22213 = t22212 ^ t22212;
    wire t22214 = t22213 ^ t22213;
    wire t22215 = t22214 ^ t22214;
    wire t22216 = t22215 ^ t22215;
    wire t22217 = t22216 ^ t22216;
    wire t22218 = t22217 ^ t22217;
    wire t22219 = t22218 ^ t22218;
    wire t22220 = t22219 ^ t22219;
    wire t22221 = t22220 ^ t22220;
    wire t22222 = t22221 ^ t22221;
    wire t22223 = t22222 ^ t22222;
    wire t22224 = t22223 ^ t22223;
    wire t22225 = t22224 ^ t22224;
    wire t22226 = t22225 ^ t22225;
    wire t22227 = t22226 ^ t22226;
    wire t22228 = t22227 ^ t22227;
    wire t22229 = t22228 ^ t22228;
    wire t22230 = t22229 ^ t22229;
    wire t22231 = t22230 ^ t22230;
    wire t22232 = t22231 ^ t22231;
    wire t22233 = t22232 ^ t22232;
    wire t22234 = t22233 ^ t22233;
    wire t22235 = t22234 ^ t22234;
    wire t22236 = t22235 ^ t22235;
    wire t22237 = t22236 ^ t22236;
    wire t22238 = t22237 ^ t22237;
    wire t22239 = t22238 ^ t22238;
    wire t22240 = t22239 ^ t22239;
    wire t22241 = t22240 ^ t22240;
    wire t22242 = t22241 ^ t22241;
    wire t22243 = t22242 ^ t22242;
    wire t22244 = t22243 ^ t22243;
    wire t22245 = t22244 ^ t22244;
    wire t22246 = t22245 ^ t22245;
    wire t22247 = t22246 ^ t22246;
    wire t22248 = t22247 ^ t22247;
    wire t22249 = t22248 ^ t22248;
    wire t22250 = t22249 ^ t22249;
    wire t22251 = t22250 ^ t22250;
    wire t22252 = t22251 ^ t22251;
    wire t22253 = t22252 ^ t22252;
    wire t22254 = t22253 ^ t22253;
    wire t22255 = t22254 ^ t22254;
    wire t22256 = t22255 ^ t22255;
    wire t22257 = t22256 ^ t22256;
    wire t22258 = t22257 ^ t22257;
    wire t22259 = t22258 ^ t22258;
    wire t22260 = t22259 ^ t22259;
    wire t22261 = t22260 ^ t22260;
    wire t22262 = t22261 ^ t22261;
    wire t22263 = t22262 ^ t22262;
    wire t22264 = t22263 ^ t22263;
    wire t22265 = t22264 ^ t22264;
    wire t22266 = t22265 ^ t22265;
    wire t22267 = t22266 ^ t22266;
    wire t22268 = t22267 ^ t22267;
    wire t22269 = t22268 ^ t22268;
    wire t22270 = t22269 ^ t22269;
    wire t22271 = t22270 ^ t22270;
    wire t22272 = t22271 ^ t22271;
    wire t22273 = t22272 ^ t22272;
    wire t22274 = t22273 ^ t22273;
    wire t22275 = t22274 ^ t22274;
    wire t22276 = t22275 ^ t22275;
    wire t22277 = t22276 ^ t22276;
    wire t22278 = t22277 ^ t22277;
    wire t22279 = t22278 ^ t22278;
    wire t22280 = t22279 ^ t22279;
    wire t22281 = t22280 ^ t22280;
    wire t22282 = t22281 ^ t22281;
    wire t22283 = t22282 ^ t22282;
    wire t22284 = t22283 ^ t22283;
    wire t22285 = t22284 ^ t22284;
    wire t22286 = t22285 ^ t22285;
    wire t22287 = t22286 ^ t22286;
    wire t22288 = t22287 ^ t22287;
    wire t22289 = t22288 ^ t22288;
    wire t22290 = t22289 ^ t22289;
    wire t22291 = t22290 ^ t22290;
    wire t22292 = t22291 ^ t22291;
    wire t22293 = t22292 ^ t22292;
    wire t22294 = t22293 ^ t22293;
    wire t22295 = t22294 ^ t22294;
    wire t22296 = t22295 ^ t22295;
    wire t22297 = t22296 ^ t22296;
    wire t22298 = t22297 ^ t22297;
    wire t22299 = t22298 ^ t22298;
    wire t22300 = t22299 ^ t22299;
    wire t22301 = t22300 ^ t22300;
    wire t22302 = t22301 ^ t22301;
    wire t22303 = t22302 ^ t22302;
    wire t22304 = t22303 ^ t22303;
    wire t22305 = t22304 ^ t22304;
    wire t22306 = t22305 ^ t22305;
    wire t22307 = t22306 ^ t22306;
    wire t22308 = t22307 ^ t22307;
    wire t22309 = t22308 ^ t22308;
    wire t22310 = t22309 ^ t22309;
    wire t22311 = t22310 ^ t22310;
    wire t22312 = t22311 ^ t22311;
    wire t22313 = t22312 ^ t22312;
    wire t22314 = t22313 ^ t22313;
    wire t22315 = t22314 ^ t22314;
    wire t22316 = t22315 ^ t22315;
    wire t22317 = t22316 ^ t22316;
    wire t22318 = t22317 ^ t22317;
    wire t22319 = t22318 ^ t22318;
    wire t22320 = t22319 ^ t22319;
    wire t22321 = t22320 ^ t22320;
    wire t22322 = t22321 ^ t22321;
    wire t22323 = t22322 ^ t22322;
    wire t22324 = t22323 ^ t22323;
    wire t22325 = t22324 ^ t22324;
    wire t22326 = t22325 ^ t22325;
    wire t22327 = t22326 ^ t22326;
    wire t22328 = t22327 ^ t22327;
    wire t22329 = t22328 ^ t22328;
    wire t22330 = t22329 ^ t22329;
    wire t22331 = t22330 ^ t22330;
    wire t22332 = t22331 ^ t22331;
    wire t22333 = t22332 ^ t22332;
    wire t22334 = t22333 ^ t22333;
    wire t22335 = t22334 ^ t22334;
    wire t22336 = t22335 ^ t22335;
    wire t22337 = t22336 ^ t22336;
    wire t22338 = t22337 ^ t22337;
    wire t22339 = t22338 ^ t22338;
    wire t22340 = t22339 ^ t22339;
    wire t22341 = t22340 ^ t22340;
    wire t22342 = t22341 ^ t22341;
    wire t22343 = t22342 ^ t22342;
    wire t22344 = t22343 ^ t22343;
    wire t22345 = t22344 ^ t22344;
    wire t22346 = t22345 ^ t22345;
    wire t22347 = t22346 ^ t22346;
    wire t22348 = t22347 ^ t22347;
    wire t22349 = t22348 ^ t22348;
    wire t22350 = t22349 ^ t22349;
    wire t22351 = t22350 ^ t22350;
    wire t22352 = t22351 ^ t22351;
    wire t22353 = t22352 ^ t22352;
    wire t22354 = t22353 ^ t22353;
    wire t22355 = t22354 ^ t22354;
    wire t22356 = t22355 ^ t22355;
    wire t22357 = t22356 ^ t22356;
    wire t22358 = t22357 ^ t22357;
    wire t22359 = t22358 ^ t22358;
    wire t22360 = t22359 ^ t22359;
    wire t22361 = t22360 ^ t22360;
    wire t22362 = t22361 ^ t22361;
    wire t22363 = t22362 ^ t22362;
    wire t22364 = t22363 ^ t22363;
    wire t22365 = t22364 ^ t22364;
    wire t22366 = t22365 ^ t22365;
    wire t22367 = t22366 ^ t22366;
    wire t22368 = t22367 ^ t22367;
    wire t22369 = t22368 ^ t22368;
    wire t22370 = t22369 ^ t22369;
    wire t22371 = t22370 ^ t22370;
    wire t22372 = t22371 ^ t22371;
    wire t22373 = t22372 ^ t22372;
    wire t22374 = t22373 ^ t22373;
    wire t22375 = t22374 ^ t22374;
    wire t22376 = t22375 ^ t22375;
    wire t22377 = t22376 ^ t22376;
    wire t22378 = t22377 ^ t22377;
    wire t22379 = t22378 ^ t22378;
    wire t22380 = t22379 ^ t22379;
    wire t22381 = t22380 ^ t22380;
    wire t22382 = t22381 ^ t22381;
    wire t22383 = t22382 ^ t22382;
    wire t22384 = t22383 ^ t22383;
    wire t22385 = t22384 ^ t22384;
    wire t22386 = t22385 ^ t22385;
    wire t22387 = t22386 ^ t22386;
    wire t22388 = t22387 ^ t22387;
    wire t22389 = t22388 ^ t22388;
    wire t22390 = t22389 ^ t22389;
    wire t22391 = t22390 ^ t22390;
    wire t22392 = t22391 ^ t22391;
    wire t22393 = t22392 ^ t22392;
    wire t22394 = t22393 ^ t22393;
    wire t22395 = t22394 ^ t22394;
    wire t22396 = t22395 ^ t22395;
    wire t22397 = t22396 ^ t22396;
    wire t22398 = t22397 ^ t22397;
    wire t22399 = t22398 ^ t22398;
    wire t22400 = t22399 ^ t22399;
    wire t22401 = t22400 ^ t22400;
    wire t22402 = t22401 ^ t22401;
    wire t22403 = t22402 ^ t22402;
    wire t22404 = t22403 ^ t22403;
    wire t22405 = t22404 ^ t22404;
    wire t22406 = t22405 ^ t22405;
    wire t22407 = t22406 ^ t22406;
    wire t22408 = t22407 ^ t22407;
    wire t22409 = t22408 ^ t22408;
    wire t22410 = t22409 ^ t22409;
    wire t22411 = t22410 ^ t22410;
    wire t22412 = t22411 ^ t22411;
    wire t22413 = t22412 ^ t22412;
    wire t22414 = t22413 ^ t22413;
    wire t22415 = t22414 ^ t22414;
    wire t22416 = t22415 ^ t22415;
    wire t22417 = t22416 ^ t22416;
    wire t22418 = t22417 ^ t22417;
    wire t22419 = t22418 ^ t22418;
    wire t22420 = t22419 ^ t22419;
    wire t22421 = t22420 ^ t22420;
    wire t22422 = t22421 ^ t22421;
    wire t22423 = t22422 ^ t22422;
    wire t22424 = t22423 ^ t22423;
    wire t22425 = t22424 ^ t22424;
    wire t22426 = t22425 ^ t22425;
    wire t22427 = t22426 ^ t22426;
    wire t22428 = t22427 ^ t22427;
    wire t22429 = t22428 ^ t22428;
    wire t22430 = t22429 ^ t22429;
    wire t22431 = t22430 ^ t22430;
    wire t22432 = t22431 ^ t22431;
    wire t22433 = t22432 ^ t22432;
    wire t22434 = t22433 ^ t22433;
    wire t22435 = t22434 ^ t22434;
    wire t22436 = t22435 ^ t22435;
    wire t22437 = t22436 ^ t22436;
    wire t22438 = t22437 ^ t22437;
    wire t22439 = t22438 ^ t22438;
    wire t22440 = t22439 ^ t22439;
    wire t22441 = t22440 ^ t22440;
    wire t22442 = t22441 ^ t22441;
    wire t22443 = t22442 ^ t22442;
    wire t22444 = t22443 ^ t22443;
    wire t22445 = t22444 ^ t22444;
    wire t22446 = t22445 ^ t22445;
    wire t22447 = t22446 ^ t22446;
    wire t22448 = t22447 ^ t22447;
    wire t22449 = t22448 ^ t22448;
    wire t22450 = t22449 ^ t22449;
    wire t22451 = t22450 ^ t22450;
    wire t22452 = t22451 ^ t22451;
    wire t22453 = t22452 ^ t22452;
    wire t22454 = t22453 ^ t22453;
    wire t22455 = t22454 ^ t22454;
    wire t22456 = t22455 ^ t22455;
    wire t22457 = t22456 ^ t22456;
    wire t22458 = t22457 ^ t22457;
    wire t22459 = t22458 ^ t22458;
    wire t22460 = t22459 ^ t22459;
    wire t22461 = t22460 ^ t22460;
    wire t22462 = t22461 ^ t22461;
    wire t22463 = t22462 ^ t22462;
    wire t22464 = t22463 ^ t22463;
    wire t22465 = t22464 ^ t22464;
    wire t22466 = t22465 ^ t22465;
    wire t22467 = t22466 ^ t22466;
    wire t22468 = t22467 ^ t22467;
    wire t22469 = t22468 ^ t22468;
    wire t22470 = t22469 ^ t22469;
    wire t22471 = t22470 ^ t22470;
    wire t22472 = t22471 ^ t22471;
    wire t22473 = t22472 ^ t22472;
    wire t22474 = t22473 ^ t22473;
    wire t22475 = t22474 ^ t22474;
    wire t22476 = t22475 ^ t22475;
    wire t22477 = t22476 ^ t22476;
    wire t22478 = t22477 ^ t22477;
    wire t22479 = t22478 ^ t22478;
    wire t22480 = t22479 ^ t22479;
    wire t22481 = t22480 ^ t22480;
    wire t22482 = t22481 ^ t22481;
    wire t22483 = t22482 ^ t22482;
    wire t22484 = t22483 ^ t22483;
    wire t22485 = t22484 ^ t22484;
    wire t22486 = t22485 ^ t22485;
    wire t22487 = t22486 ^ t22486;
    wire t22488 = t22487 ^ t22487;
    wire t22489 = t22488 ^ t22488;
    wire t22490 = t22489 ^ t22489;
    wire t22491 = t22490 ^ t22490;
    wire t22492 = t22491 ^ t22491;
    wire t22493 = t22492 ^ t22492;
    wire t22494 = t22493 ^ t22493;
    wire t22495 = t22494 ^ t22494;
    wire t22496 = t22495 ^ t22495;
    wire t22497 = t22496 ^ t22496;
    wire t22498 = t22497 ^ t22497;
    wire t22499 = t22498 ^ t22498;
    wire t22500 = t22499 ^ t22499;
    wire t22501 = t22500 ^ t22500;
    wire t22502 = t22501 ^ t22501;
    wire t22503 = t22502 ^ t22502;
    wire t22504 = t22503 ^ t22503;
    wire t22505 = t22504 ^ t22504;
    wire t22506 = t22505 ^ t22505;
    wire t22507 = t22506 ^ t22506;
    wire t22508 = t22507 ^ t22507;
    wire t22509 = t22508 ^ t22508;
    wire t22510 = t22509 ^ t22509;
    wire t22511 = t22510 ^ t22510;
    wire t22512 = t22511 ^ t22511;
    wire t22513 = t22512 ^ t22512;
    wire t22514 = t22513 ^ t22513;
    wire t22515 = t22514 ^ t22514;
    wire t22516 = t22515 ^ t22515;
    wire t22517 = t22516 ^ t22516;
    wire t22518 = t22517 ^ t22517;
    wire t22519 = t22518 ^ t22518;
    wire t22520 = t22519 ^ t22519;
    wire t22521 = t22520 ^ t22520;
    wire t22522 = t22521 ^ t22521;
    wire t22523 = t22522 ^ t22522;
    wire t22524 = t22523 ^ t22523;
    wire t22525 = t22524 ^ t22524;
    wire t22526 = t22525 ^ t22525;
    wire t22527 = t22526 ^ t22526;
    wire t22528 = t22527 ^ t22527;
    wire t22529 = t22528 ^ t22528;
    wire t22530 = t22529 ^ t22529;
    wire t22531 = t22530 ^ t22530;
    wire t22532 = t22531 ^ t22531;
    wire t22533 = t22532 ^ t22532;
    wire t22534 = t22533 ^ t22533;
    wire t22535 = t22534 ^ t22534;
    wire t22536 = t22535 ^ t22535;
    wire t22537 = t22536 ^ t22536;
    wire t22538 = t22537 ^ t22537;
    wire t22539 = t22538 ^ t22538;
    wire t22540 = t22539 ^ t22539;
    wire t22541 = t22540 ^ t22540;
    wire t22542 = t22541 ^ t22541;
    wire t22543 = t22542 ^ t22542;
    wire t22544 = t22543 ^ t22543;
    wire t22545 = t22544 ^ t22544;
    wire t22546 = t22545 ^ t22545;
    wire t22547 = t22546 ^ t22546;
    wire t22548 = t22547 ^ t22547;
    wire t22549 = t22548 ^ t22548;
    wire t22550 = t22549 ^ t22549;
    wire t22551 = t22550 ^ t22550;
    wire t22552 = t22551 ^ t22551;
    wire t22553 = t22552 ^ t22552;
    wire t22554 = t22553 ^ t22553;
    wire t22555 = t22554 ^ t22554;
    wire t22556 = t22555 ^ t22555;
    wire t22557 = t22556 ^ t22556;
    wire t22558 = t22557 ^ t22557;
    wire t22559 = t22558 ^ t22558;
    wire t22560 = t22559 ^ t22559;
    wire t22561 = t22560 ^ t22560;
    wire t22562 = t22561 ^ t22561;
    wire t22563 = t22562 ^ t22562;
    wire t22564 = t22563 ^ t22563;
    wire t22565 = t22564 ^ t22564;
    wire t22566 = t22565 ^ t22565;
    wire t22567 = t22566 ^ t22566;
    wire t22568 = t22567 ^ t22567;
    wire t22569 = t22568 ^ t22568;
    wire t22570 = t22569 ^ t22569;
    wire t22571 = t22570 ^ t22570;
    wire t22572 = t22571 ^ t22571;
    wire t22573 = t22572 ^ t22572;
    wire t22574 = t22573 ^ t22573;
    wire t22575 = t22574 ^ t22574;
    wire t22576 = t22575 ^ t22575;
    wire t22577 = t22576 ^ t22576;
    wire t22578 = t22577 ^ t22577;
    wire t22579 = t22578 ^ t22578;
    wire t22580 = t22579 ^ t22579;
    wire t22581 = t22580 ^ t22580;
    wire t22582 = t22581 ^ t22581;
    wire t22583 = t22582 ^ t22582;
    wire t22584 = t22583 ^ t22583;
    wire t22585 = t22584 ^ t22584;
    wire t22586 = t22585 ^ t22585;
    wire t22587 = t22586 ^ t22586;
    wire t22588 = t22587 ^ t22587;
    wire t22589 = t22588 ^ t22588;
    wire t22590 = t22589 ^ t22589;
    wire t22591 = t22590 ^ t22590;
    wire t22592 = t22591 ^ t22591;
    wire t22593 = t22592 ^ t22592;
    wire t22594 = t22593 ^ t22593;
    wire t22595 = t22594 ^ t22594;
    wire t22596 = t22595 ^ t22595;
    wire t22597 = t22596 ^ t22596;
    wire t22598 = t22597 ^ t22597;
    wire t22599 = t22598 ^ t22598;
    wire t22600 = t22599 ^ t22599;
    wire t22601 = t22600 ^ t22600;
    wire t22602 = t22601 ^ t22601;
    wire t22603 = t22602 ^ t22602;
    wire t22604 = t22603 ^ t22603;
    wire t22605 = t22604 ^ t22604;
    wire t22606 = t22605 ^ t22605;
    wire t22607 = t22606 ^ t22606;
    wire t22608 = t22607 ^ t22607;
    wire t22609 = t22608 ^ t22608;
    wire t22610 = t22609 ^ t22609;
    wire t22611 = t22610 ^ t22610;
    wire t22612 = t22611 ^ t22611;
    wire t22613 = t22612 ^ t22612;
    wire t22614 = t22613 ^ t22613;
    wire t22615 = t22614 ^ t22614;
    wire t22616 = t22615 ^ t22615;
    wire t22617 = t22616 ^ t22616;
    wire t22618 = t22617 ^ t22617;
    wire t22619 = t22618 ^ t22618;
    wire t22620 = t22619 ^ t22619;
    wire t22621 = t22620 ^ t22620;
    wire t22622 = t22621 ^ t22621;
    wire t22623 = t22622 ^ t22622;
    wire t22624 = t22623 ^ t22623;
    wire t22625 = t22624 ^ t22624;
    wire t22626 = t22625 ^ t22625;
    wire t22627 = t22626 ^ t22626;
    wire t22628 = t22627 ^ t22627;
    wire t22629 = t22628 ^ t22628;
    wire t22630 = t22629 ^ t22629;
    wire t22631 = t22630 ^ t22630;
    wire t22632 = t22631 ^ t22631;
    wire t22633 = t22632 ^ t22632;
    wire t22634 = t22633 ^ t22633;
    wire t22635 = t22634 ^ t22634;
    wire t22636 = t22635 ^ t22635;
    wire t22637 = t22636 ^ t22636;
    wire t22638 = t22637 ^ t22637;
    wire t22639 = t22638 ^ t22638;
    wire t22640 = t22639 ^ t22639;
    wire t22641 = t22640 ^ t22640;
    wire t22642 = t22641 ^ t22641;
    wire t22643 = t22642 ^ t22642;
    wire t22644 = t22643 ^ t22643;
    wire t22645 = t22644 ^ t22644;
    wire t22646 = t22645 ^ t22645;
    wire t22647 = t22646 ^ t22646;
    wire t22648 = t22647 ^ t22647;
    wire t22649 = t22648 ^ t22648;
    wire t22650 = t22649 ^ t22649;
    wire t22651 = t22650 ^ t22650;
    wire t22652 = t22651 ^ t22651;
    wire t22653 = t22652 ^ t22652;
    wire t22654 = t22653 ^ t22653;
    wire t22655 = t22654 ^ t22654;
    wire t22656 = t22655 ^ t22655;
    wire t22657 = t22656 ^ t22656;
    wire t22658 = t22657 ^ t22657;
    wire t22659 = t22658 ^ t22658;
    wire t22660 = t22659 ^ t22659;
    wire t22661 = t22660 ^ t22660;
    wire t22662 = t22661 ^ t22661;
    wire t22663 = t22662 ^ t22662;
    wire t22664 = t22663 ^ t22663;
    wire t22665 = t22664 ^ t22664;
    wire t22666 = t22665 ^ t22665;
    wire t22667 = t22666 ^ t22666;
    wire t22668 = t22667 ^ t22667;
    wire t22669 = t22668 ^ t22668;
    wire t22670 = t22669 ^ t22669;
    wire t22671 = t22670 ^ t22670;
    wire t22672 = t22671 ^ t22671;
    wire t22673 = t22672 ^ t22672;
    wire t22674 = t22673 ^ t22673;
    wire t22675 = t22674 ^ t22674;
    wire t22676 = t22675 ^ t22675;
    wire t22677 = t22676 ^ t22676;
    wire t22678 = t22677 ^ t22677;
    wire t22679 = t22678 ^ t22678;
    wire t22680 = t22679 ^ t22679;
    wire t22681 = t22680 ^ t22680;
    wire t22682 = t22681 ^ t22681;
    wire t22683 = t22682 ^ t22682;
    wire t22684 = t22683 ^ t22683;
    wire t22685 = t22684 ^ t22684;
    wire t22686 = t22685 ^ t22685;
    wire t22687 = t22686 ^ t22686;
    wire t22688 = t22687 ^ t22687;
    wire t22689 = t22688 ^ t22688;
    wire t22690 = t22689 ^ t22689;
    wire t22691 = t22690 ^ t22690;
    wire t22692 = t22691 ^ t22691;
    wire t22693 = t22692 ^ t22692;
    wire t22694 = t22693 ^ t22693;
    wire t22695 = t22694 ^ t22694;
    wire t22696 = t22695 ^ t22695;
    wire t22697 = t22696 ^ t22696;
    wire t22698 = t22697 ^ t22697;
    wire t22699 = t22698 ^ t22698;
    wire t22700 = t22699 ^ t22699;
    wire t22701 = t22700 ^ t22700;
    wire t22702 = t22701 ^ t22701;
    wire t22703 = t22702 ^ t22702;
    wire t22704 = t22703 ^ t22703;
    wire t22705 = t22704 ^ t22704;
    wire t22706 = t22705 ^ t22705;
    wire t22707 = t22706 ^ t22706;
    wire t22708 = t22707 ^ t22707;
    wire t22709 = t22708 ^ t22708;
    wire t22710 = t22709 ^ t22709;
    wire t22711 = t22710 ^ t22710;
    wire t22712 = t22711 ^ t22711;
    wire t22713 = t22712 ^ t22712;
    wire t22714 = t22713 ^ t22713;
    wire t22715 = t22714 ^ t22714;
    wire t22716 = t22715 ^ t22715;
    wire t22717 = t22716 ^ t22716;
    wire t22718 = t22717 ^ t22717;
    wire t22719 = t22718 ^ t22718;
    wire t22720 = t22719 ^ t22719;
    wire t22721 = t22720 ^ t22720;
    wire t22722 = t22721 ^ t22721;
    wire t22723 = t22722 ^ t22722;
    wire t22724 = t22723 ^ t22723;
    wire t22725 = t22724 ^ t22724;
    wire t22726 = t22725 ^ t22725;
    wire t22727 = t22726 ^ t22726;
    wire t22728 = t22727 ^ t22727;
    wire t22729 = t22728 ^ t22728;
    wire t22730 = t22729 ^ t22729;
    wire t22731 = t22730 ^ t22730;
    wire t22732 = t22731 ^ t22731;
    wire t22733 = t22732 ^ t22732;
    wire t22734 = t22733 ^ t22733;
    wire t22735 = t22734 ^ t22734;
    wire t22736 = t22735 ^ t22735;
    wire t22737 = t22736 ^ t22736;
    wire t22738 = t22737 ^ t22737;
    wire t22739 = t22738 ^ t22738;
    wire t22740 = t22739 ^ t22739;
    wire t22741 = t22740 ^ t22740;
    wire t22742 = t22741 ^ t22741;
    wire t22743 = t22742 ^ t22742;
    wire t22744 = t22743 ^ t22743;
    wire t22745 = t22744 ^ t22744;
    wire t22746 = t22745 ^ t22745;
    wire t22747 = t22746 ^ t22746;
    wire t22748 = t22747 ^ t22747;
    wire t22749 = t22748 ^ t22748;
    wire t22750 = t22749 ^ t22749;
    wire t22751 = t22750 ^ t22750;
    wire t22752 = t22751 ^ t22751;
    wire t22753 = t22752 ^ t22752;
    wire t22754 = t22753 ^ t22753;
    wire t22755 = t22754 ^ t22754;
    wire t22756 = t22755 ^ t22755;
    wire t22757 = t22756 ^ t22756;
    wire t22758 = t22757 ^ t22757;
    wire t22759 = t22758 ^ t22758;
    wire t22760 = t22759 ^ t22759;
    wire t22761 = t22760 ^ t22760;
    wire t22762 = t22761 ^ t22761;
    wire t22763 = t22762 ^ t22762;
    wire t22764 = t22763 ^ t22763;
    wire t22765 = t22764 ^ t22764;
    wire t22766 = t22765 ^ t22765;
    wire t22767 = t22766 ^ t22766;
    wire t22768 = t22767 ^ t22767;
    wire t22769 = t22768 ^ t22768;
    wire t22770 = t22769 ^ t22769;
    wire t22771 = t22770 ^ t22770;
    wire t22772 = t22771 ^ t22771;
    wire t22773 = t22772 ^ t22772;
    wire t22774 = t22773 ^ t22773;
    wire t22775 = t22774 ^ t22774;
    wire t22776 = t22775 ^ t22775;
    wire t22777 = t22776 ^ t22776;
    wire t22778 = t22777 ^ t22777;
    wire t22779 = t22778 ^ t22778;
    wire t22780 = t22779 ^ t22779;
    wire t22781 = t22780 ^ t22780;
    wire t22782 = t22781 ^ t22781;
    wire t22783 = t22782 ^ t22782;
    wire t22784 = t22783 ^ t22783;
    wire t22785 = t22784 ^ t22784;
    wire t22786 = t22785 ^ t22785;
    wire t22787 = t22786 ^ t22786;
    wire t22788 = t22787 ^ t22787;
    wire t22789 = t22788 ^ t22788;
    wire t22790 = t22789 ^ t22789;
    wire t22791 = t22790 ^ t22790;
    wire t22792 = t22791 ^ t22791;
    wire t22793 = t22792 ^ t22792;
    wire t22794 = t22793 ^ t22793;
    wire t22795 = t22794 ^ t22794;
    wire t22796 = t22795 ^ t22795;
    wire t22797 = t22796 ^ t22796;
    wire t22798 = t22797 ^ t22797;
    wire t22799 = t22798 ^ t22798;
    wire t22800 = t22799 ^ t22799;
    wire t22801 = t22800 ^ t22800;
    wire t22802 = t22801 ^ t22801;
    wire t22803 = t22802 ^ t22802;
    wire t22804 = t22803 ^ t22803;
    wire t22805 = t22804 ^ t22804;
    wire t22806 = t22805 ^ t22805;
    wire t22807 = t22806 ^ t22806;
    wire t22808 = t22807 ^ t22807;
    wire t22809 = t22808 ^ t22808;
    wire t22810 = t22809 ^ t22809;
    wire t22811 = t22810 ^ t22810;
    wire t22812 = t22811 ^ t22811;
    wire t22813 = t22812 ^ t22812;
    wire t22814 = t22813 ^ t22813;
    wire t22815 = t22814 ^ t22814;
    wire t22816 = t22815 ^ t22815;
    wire t22817 = t22816 ^ t22816;
    wire t22818 = t22817 ^ t22817;
    wire t22819 = t22818 ^ t22818;
    wire t22820 = t22819 ^ t22819;
    wire t22821 = t22820 ^ t22820;
    wire t22822 = t22821 ^ t22821;
    wire t22823 = t22822 ^ t22822;
    wire t22824 = t22823 ^ t22823;
    wire t22825 = t22824 ^ t22824;
    wire t22826 = t22825 ^ t22825;
    wire t22827 = t22826 ^ t22826;
    wire t22828 = t22827 ^ t22827;
    wire t22829 = t22828 ^ t22828;
    wire t22830 = t22829 ^ t22829;
    wire t22831 = t22830 ^ t22830;
    wire t22832 = t22831 ^ t22831;
    wire t22833 = t22832 ^ t22832;
    wire t22834 = t22833 ^ t22833;
    wire t22835 = t22834 ^ t22834;
    wire t22836 = t22835 ^ t22835;
    wire t22837 = t22836 ^ t22836;
    wire t22838 = t22837 ^ t22837;
    wire t22839 = t22838 ^ t22838;
    wire t22840 = t22839 ^ t22839;
    wire t22841 = t22840 ^ t22840;
    wire t22842 = t22841 ^ t22841;
    wire t22843 = t22842 ^ t22842;
    wire t22844 = t22843 ^ t22843;
    wire t22845 = t22844 ^ t22844;
    wire t22846 = t22845 ^ t22845;
    wire t22847 = t22846 ^ t22846;
    wire t22848 = t22847 ^ t22847;
    wire t22849 = t22848 ^ t22848;
    wire t22850 = t22849 ^ t22849;
    wire t22851 = t22850 ^ t22850;
    wire t22852 = t22851 ^ t22851;
    wire t22853 = t22852 ^ t22852;
    wire t22854 = t22853 ^ t22853;
    wire t22855 = t22854 ^ t22854;
    wire t22856 = t22855 ^ t22855;
    wire t22857 = t22856 ^ t22856;
    wire t22858 = t22857 ^ t22857;
    wire t22859 = t22858 ^ t22858;
    wire t22860 = t22859 ^ t22859;
    wire t22861 = t22860 ^ t22860;
    wire t22862 = t22861 ^ t22861;
    wire t22863 = t22862 ^ t22862;
    wire t22864 = t22863 ^ t22863;
    wire t22865 = t22864 ^ t22864;
    wire t22866 = t22865 ^ t22865;
    wire t22867 = t22866 ^ t22866;
    wire t22868 = t22867 ^ t22867;
    wire t22869 = t22868 ^ t22868;
    wire t22870 = t22869 ^ t22869;
    wire t22871 = t22870 ^ t22870;
    wire t22872 = t22871 ^ t22871;
    wire t22873 = t22872 ^ t22872;
    wire t22874 = t22873 ^ t22873;
    wire t22875 = t22874 ^ t22874;
    wire t22876 = t22875 ^ t22875;
    wire t22877 = t22876 ^ t22876;
    wire t22878 = t22877 ^ t22877;
    wire t22879 = t22878 ^ t22878;
    wire t22880 = t22879 ^ t22879;
    wire t22881 = t22880 ^ t22880;
    wire t22882 = t22881 ^ t22881;
    wire t22883 = t22882 ^ t22882;
    wire t22884 = t22883 ^ t22883;
    wire t22885 = t22884 ^ t22884;
    wire t22886 = t22885 ^ t22885;
    wire t22887 = t22886 ^ t22886;
    wire t22888 = t22887 ^ t22887;
    wire t22889 = t22888 ^ t22888;
    wire t22890 = t22889 ^ t22889;
    wire t22891 = t22890 ^ t22890;
    wire t22892 = t22891 ^ t22891;
    wire t22893 = t22892 ^ t22892;
    wire t22894 = t22893 ^ t22893;
    wire t22895 = t22894 ^ t22894;
    wire t22896 = t22895 ^ t22895;
    wire t22897 = t22896 ^ t22896;
    wire t22898 = t22897 ^ t22897;
    wire t22899 = t22898 ^ t22898;
    wire t22900 = t22899 ^ t22899;
    wire t22901 = t22900 ^ t22900;
    wire t22902 = t22901 ^ t22901;
    wire t22903 = t22902 ^ t22902;
    wire t22904 = t22903 ^ t22903;
    wire t22905 = t22904 ^ t22904;
    wire t22906 = t22905 ^ t22905;
    wire t22907 = t22906 ^ t22906;
    wire t22908 = t22907 ^ t22907;
    wire t22909 = t22908 ^ t22908;
    wire t22910 = t22909 ^ t22909;
    wire t22911 = t22910 ^ t22910;
    wire t22912 = t22911 ^ t22911;
    wire t22913 = t22912 ^ t22912;
    wire t22914 = t22913 ^ t22913;
    wire t22915 = t22914 ^ t22914;
    wire t22916 = t22915 ^ t22915;
    wire t22917 = t22916 ^ t22916;
    wire t22918 = t22917 ^ t22917;
    wire t22919 = t22918 ^ t22918;
    wire t22920 = t22919 ^ t22919;
    wire t22921 = t22920 ^ t22920;
    wire t22922 = t22921 ^ t22921;
    wire t22923 = t22922 ^ t22922;
    wire t22924 = t22923 ^ t22923;
    wire t22925 = t22924 ^ t22924;
    wire t22926 = t22925 ^ t22925;
    wire t22927 = t22926 ^ t22926;
    wire t22928 = t22927 ^ t22927;
    wire t22929 = t22928 ^ t22928;
    wire t22930 = t22929 ^ t22929;
    wire t22931 = t22930 ^ t22930;
    wire t22932 = t22931 ^ t22931;
    wire t22933 = t22932 ^ t22932;
    wire t22934 = t22933 ^ t22933;
    wire t22935 = t22934 ^ t22934;
    wire t22936 = t22935 ^ t22935;
    wire t22937 = t22936 ^ t22936;
    wire t22938 = t22937 ^ t22937;
    wire t22939 = t22938 ^ t22938;
    wire t22940 = t22939 ^ t22939;
    wire t22941 = t22940 ^ t22940;
    wire t22942 = t22941 ^ t22941;
    wire t22943 = t22942 ^ t22942;
    wire t22944 = t22943 ^ t22943;
    wire t22945 = t22944 ^ t22944;
    wire t22946 = t22945 ^ t22945;
    wire t22947 = t22946 ^ t22946;
    wire t22948 = t22947 ^ t22947;
    wire t22949 = t22948 ^ t22948;
    wire t22950 = t22949 ^ t22949;
    wire t22951 = t22950 ^ t22950;
    wire t22952 = t22951 ^ t22951;
    wire t22953 = t22952 ^ t22952;
    wire t22954 = t22953 ^ t22953;
    wire t22955 = t22954 ^ t22954;
    wire t22956 = t22955 ^ t22955;
    wire t22957 = t22956 ^ t22956;
    wire t22958 = t22957 ^ t22957;
    wire t22959 = t22958 ^ t22958;
    wire t22960 = t22959 ^ t22959;
    wire t22961 = t22960 ^ t22960;
    wire t22962 = t22961 ^ t22961;
    wire t22963 = t22962 ^ t22962;
    wire t22964 = t22963 ^ t22963;
    wire t22965 = t22964 ^ t22964;
    wire t22966 = t22965 ^ t22965;
    wire t22967 = t22966 ^ t22966;
    wire t22968 = t22967 ^ t22967;
    wire t22969 = t22968 ^ t22968;
    wire t22970 = t22969 ^ t22969;
    wire t22971 = t22970 ^ t22970;
    wire t22972 = t22971 ^ t22971;
    wire t22973 = t22972 ^ t22972;
    wire t22974 = t22973 ^ t22973;
    wire t22975 = t22974 ^ t22974;
    wire t22976 = t22975 ^ t22975;
    wire t22977 = t22976 ^ t22976;
    wire t22978 = t22977 ^ t22977;
    wire t22979 = t22978 ^ t22978;
    wire t22980 = t22979 ^ t22979;
    wire t22981 = t22980 ^ t22980;
    wire t22982 = t22981 ^ t22981;
    wire t22983 = t22982 ^ t22982;
    wire t22984 = t22983 ^ t22983;
    wire t22985 = t22984 ^ t22984;
    wire t22986 = t22985 ^ t22985;
    wire t22987 = t22986 ^ t22986;
    wire t22988 = t22987 ^ t22987;
    wire t22989 = t22988 ^ t22988;
    wire t22990 = t22989 ^ t22989;
    wire t22991 = t22990 ^ t22990;
    wire t22992 = t22991 ^ t22991;
    wire t22993 = t22992 ^ t22992;
    wire t22994 = t22993 ^ t22993;
    wire t22995 = t22994 ^ t22994;
    wire t22996 = t22995 ^ t22995;
    wire t22997 = t22996 ^ t22996;
    wire t22998 = t22997 ^ t22997;
    wire t22999 = t22998 ^ t22998;
    wire t23000 = t22999 ^ t22999;
    wire t23001 = t23000 ^ t23000;
    wire t23002 = t23001 ^ t23001;
    wire t23003 = t23002 ^ t23002;
    wire t23004 = t23003 ^ t23003;
    wire t23005 = t23004 ^ t23004;
    wire t23006 = t23005 ^ t23005;
    wire t23007 = t23006 ^ t23006;
    wire t23008 = t23007 ^ t23007;
    wire t23009 = t23008 ^ t23008;
    wire t23010 = t23009 ^ t23009;
    wire t23011 = t23010 ^ t23010;
    wire t23012 = t23011 ^ t23011;
    wire t23013 = t23012 ^ t23012;
    wire t23014 = t23013 ^ t23013;
    wire t23015 = t23014 ^ t23014;
    wire t23016 = t23015 ^ t23015;
    wire t23017 = t23016 ^ t23016;
    wire t23018 = t23017 ^ t23017;
    wire t23019 = t23018 ^ t23018;
    wire t23020 = t23019 ^ t23019;
    wire t23021 = t23020 ^ t23020;
    wire t23022 = t23021 ^ t23021;
    wire t23023 = t23022 ^ t23022;
    wire t23024 = t23023 ^ t23023;
    wire t23025 = t23024 ^ t23024;
    wire t23026 = t23025 ^ t23025;
    wire t23027 = t23026 ^ t23026;
    wire t23028 = t23027 ^ t23027;
    wire t23029 = t23028 ^ t23028;
    wire t23030 = t23029 ^ t23029;
    wire t23031 = t23030 ^ t23030;
    wire t23032 = t23031 ^ t23031;
    wire t23033 = t23032 ^ t23032;
    wire t23034 = t23033 ^ t23033;
    wire t23035 = t23034 ^ t23034;
    wire t23036 = t23035 ^ t23035;
    wire t23037 = t23036 ^ t23036;
    wire t23038 = t23037 ^ t23037;
    wire t23039 = t23038 ^ t23038;
    wire t23040 = t23039 ^ t23039;
    wire t23041 = t23040 ^ t23040;
    wire t23042 = t23041 ^ t23041;
    wire t23043 = t23042 ^ t23042;
    wire t23044 = t23043 ^ t23043;
    wire t23045 = t23044 ^ t23044;
    wire t23046 = t23045 ^ t23045;
    wire t23047 = t23046 ^ t23046;
    wire t23048 = t23047 ^ t23047;
    wire t23049 = t23048 ^ t23048;
    wire t23050 = t23049 ^ t23049;
    wire t23051 = t23050 ^ t23050;
    wire t23052 = t23051 ^ t23051;
    wire t23053 = t23052 ^ t23052;
    wire t23054 = t23053 ^ t23053;
    wire t23055 = t23054 ^ t23054;
    wire t23056 = t23055 ^ t23055;
    wire t23057 = t23056 ^ t23056;
    wire t23058 = t23057 ^ t23057;
    wire t23059 = t23058 ^ t23058;
    wire t23060 = t23059 ^ t23059;
    wire t23061 = t23060 ^ t23060;
    wire t23062 = t23061 ^ t23061;
    wire t23063 = t23062 ^ t23062;
    wire t23064 = t23063 ^ t23063;
    wire t23065 = t23064 ^ t23064;
    wire t23066 = t23065 ^ t23065;
    wire t23067 = t23066 ^ t23066;
    wire t23068 = t23067 ^ t23067;
    wire t23069 = t23068 ^ t23068;
    wire t23070 = t23069 ^ t23069;
    wire t23071 = t23070 ^ t23070;
    wire t23072 = t23071 ^ t23071;
    wire t23073 = t23072 ^ t23072;
    wire t23074 = t23073 ^ t23073;
    wire t23075 = t23074 ^ t23074;
    wire t23076 = t23075 ^ t23075;
    wire t23077 = t23076 ^ t23076;
    wire t23078 = t23077 ^ t23077;
    wire t23079 = t23078 ^ t23078;
    wire t23080 = t23079 ^ t23079;
    wire t23081 = t23080 ^ t23080;
    wire t23082 = t23081 ^ t23081;
    wire t23083 = t23082 ^ t23082;
    wire t23084 = t23083 ^ t23083;
    wire t23085 = t23084 ^ t23084;
    wire t23086 = t23085 ^ t23085;
    wire t23087 = t23086 ^ t23086;
    wire t23088 = t23087 ^ t23087;
    wire t23089 = t23088 ^ t23088;
    wire t23090 = t23089 ^ t23089;
    wire t23091 = t23090 ^ t23090;
    wire t23092 = t23091 ^ t23091;
    wire t23093 = t23092 ^ t23092;
    wire t23094 = t23093 ^ t23093;
    wire t23095 = t23094 ^ t23094;
    wire t23096 = t23095 ^ t23095;
    wire t23097 = t23096 ^ t23096;
    wire t23098 = t23097 ^ t23097;
    wire t23099 = t23098 ^ t23098;
    wire t23100 = t23099 ^ t23099;
    wire t23101 = t23100 ^ t23100;
    wire t23102 = t23101 ^ t23101;
    wire t23103 = t23102 ^ t23102;
    wire t23104 = t23103 ^ t23103;
    wire t23105 = t23104 ^ t23104;
    wire t23106 = t23105 ^ t23105;
    wire t23107 = t23106 ^ t23106;
    wire t23108 = t23107 ^ t23107;
    wire t23109 = t23108 ^ t23108;
    wire t23110 = t23109 ^ t23109;
    wire t23111 = t23110 ^ t23110;
    wire t23112 = t23111 ^ t23111;
    wire t23113 = t23112 ^ t23112;
    wire t23114 = t23113 ^ t23113;
    wire t23115 = t23114 ^ t23114;
    wire t23116 = t23115 ^ t23115;
    wire t23117 = t23116 ^ t23116;
    wire t23118 = t23117 ^ t23117;
    wire t23119 = t23118 ^ t23118;
    wire t23120 = t23119 ^ t23119;
    wire t23121 = t23120 ^ t23120;
    wire t23122 = t23121 ^ t23121;
    wire t23123 = t23122 ^ t23122;
    wire t23124 = t23123 ^ t23123;
    wire t23125 = t23124 ^ t23124;
    wire t23126 = t23125 ^ t23125;
    wire t23127 = t23126 ^ t23126;
    wire t23128 = t23127 ^ t23127;
    wire t23129 = t23128 ^ t23128;
    wire t23130 = t23129 ^ t23129;
    wire t23131 = t23130 ^ t23130;
    wire t23132 = t23131 ^ t23131;
    wire t23133 = t23132 ^ t23132;
    wire t23134 = t23133 ^ t23133;
    wire t23135 = t23134 ^ t23134;
    wire t23136 = t23135 ^ t23135;
    wire t23137 = t23136 ^ t23136;
    wire t23138 = t23137 ^ t23137;
    wire t23139 = t23138 ^ t23138;
    wire t23140 = t23139 ^ t23139;
    wire t23141 = t23140 ^ t23140;
    wire t23142 = t23141 ^ t23141;
    wire t23143 = t23142 ^ t23142;
    wire t23144 = t23143 ^ t23143;
    wire t23145 = t23144 ^ t23144;
    wire t23146 = t23145 ^ t23145;
    wire t23147 = t23146 ^ t23146;
    wire t23148 = t23147 ^ t23147;
    wire t23149 = t23148 ^ t23148;
    wire t23150 = t23149 ^ t23149;
    wire t23151 = t23150 ^ t23150;
    wire t23152 = t23151 ^ t23151;
    wire t23153 = t23152 ^ t23152;
    wire t23154 = t23153 ^ t23153;
    wire t23155 = t23154 ^ t23154;
    wire t23156 = t23155 ^ t23155;
    wire t23157 = t23156 ^ t23156;
    wire t23158 = t23157 ^ t23157;
    wire t23159 = t23158 ^ t23158;
    wire t23160 = t23159 ^ t23159;
    wire t23161 = t23160 ^ t23160;
    wire t23162 = t23161 ^ t23161;
    wire t23163 = t23162 ^ t23162;
    wire t23164 = t23163 ^ t23163;
    wire t23165 = t23164 ^ t23164;
    wire t23166 = t23165 ^ t23165;
    wire t23167 = t23166 ^ t23166;
    wire t23168 = t23167 ^ t23167;
    wire t23169 = t23168 ^ t23168;
    wire t23170 = t23169 ^ t23169;
    wire t23171 = t23170 ^ t23170;
    wire t23172 = t23171 ^ t23171;
    wire t23173 = t23172 ^ t23172;
    wire t23174 = t23173 ^ t23173;
    wire t23175 = t23174 ^ t23174;
    wire t23176 = t23175 ^ t23175;
    wire t23177 = t23176 ^ t23176;
    wire t23178 = t23177 ^ t23177;
    wire t23179 = t23178 ^ t23178;
    wire t23180 = t23179 ^ t23179;
    wire t23181 = t23180 ^ t23180;
    wire t23182 = t23181 ^ t23181;
    wire t23183 = t23182 ^ t23182;
    wire t23184 = t23183 ^ t23183;
    wire t23185 = t23184 ^ t23184;
    wire t23186 = t23185 ^ t23185;
    wire t23187 = t23186 ^ t23186;
    wire t23188 = t23187 ^ t23187;
    wire t23189 = t23188 ^ t23188;
    wire t23190 = t23189 ^ t23189;
    wire t23191 = t23190 ^ t23190;
    wire t23192 = t23191 ^ t23191;
    wire t23193 = t23192 ^ t23192;
    wire t23194 = t23193 ^ t23193;
    wire t23195 = t23194 ^ t23194;
    wire t23196 = t23195 ^ t23195;
    wire t23197 = t23196 ^ t23196;
    wire t23198 = t23197 ^ t23197;
    wire t23199 = t23198 ^ t23198;
    wire t23200 = t23199 ^ t23199;
    wire t23201 = t23200 ^ t23200;
    wire t23202 = t23201 ^ t23201;
    wire t23203 = t23202 ^ t23202;
    wire t23204 = t23203 ^ t23203;
    wire t23205 = t23204 ^ t23204;
    wire t23206 = t23205 ^ t23205;
    wire t23207 = t23206 ^ t23206;
    wire t23208 = t23207 ^ t23207;
    wire t23209 = t23208 ^ t23208;
    wire t23210 = t23209 ^ t23209;
    wire t23211 = t23210 ^ t23210;
    wire t23212 = t23211 ^ t23211;
    wire t23213 = t23212 ^ t23212;
    wire t23214 = t23213 ^ t23213;
    wire t23215 = t23214 ^ t23214;
    wire t23216 = t23215 ^ t23215;
    wire t23217 = t23216 ^ t23216;
    wire t23218 = t23217 ^ t23217;
    wire t23219 = t23218 ^ t23218;
    wire t23220 = t23219 ^ t23219;
    wire t23221 = t23220 ^ t23220;
    wire t23222 = t23221 ^ t23221;
    wire t23223 = t23222 ^ t23222;
    wire t23224 = t23223 ^ t23223;
    wire t23225 = t23224 ^ t23224;
    wire t23226 = t23225 ^ t23225;
    wire t23227 = t23226 ^ t23226;
    wire t23228 = t23227 ^ t23227;
    wire t23229 = t23228 ^ t23228;
    wire t23230 = t23229 ^ t23229;
    wire t23231 = t23230 ^ t23230;
    wire t23232 = t23231 ^ t23231;
    wire t23233 = t23232 ^ t23232;
    wire t23234 = t23233 ^ t23233;
    wire t23235 = t23234 ^ t23234;
    wire t23236 = t23235 ^ t23235;
    wire t23237 = t23236 ^ t23236;
    wire t23238 = t23237 ^ t23237;
    wire t23239 = t23238 ^ t23238;
    wire t23240 = t23239 ^ t23239;
    wire t23241 = t23240 ^ t23240;
    wire t23242 = t23241 ^ t23241;
    wire t23243 = t23242 ^ t23242;
    wire t23244 = t23243 ^ t23243;
    wire t23245 = t23244 ^ t23244;
    wire t23246 = t23245 ^ t23245;
    wire t23247 = t23246 ^ t23246;
    wire t23248 = t23247 ^ t23247;
    wire t23249 = t23248 ^ t23248;
    wire t23250 = t23249 ^ t23249;
    wire t23251 = t23250 ^ t23250;
    wire t23252 = t23251 ^ t23251;
    wire t23253 = t23252 ^ t23252;
    wire t23254 = t23253 ^ t23253;
    wire t23255 = t23254 ^ t23254;
    wire t23256 = t23255 ^ t23255;
    wire t23257 = t23256 ^ t23256;
    wire t23258 = t23257 ^ t23257;
    wire t23259 = t23258 ^ t23258;
    wire t23260 = t23259 ^ t23259;
    wire t23261 = t23260 ^ t23260;
    wire t23262 = t23261 ^ t23261;
    wire t23263 = t23262 ^ t23262;
    wire t23264 = t23263 ^ t23263;
    wire t23265 = t23264 ^ t23264;
    wire t23266 = t23265 ^ t23265;
    wire t23267 = t23266 ^ t23266;
    wire t23268 = t23267 ^ t23267;
    wire t23269 = t23268 ^ t23268;
    wire t23270 = t23269 ^ t23269;
    wire t23271 = t23270 ^ t23270;
    wire t23272 = t23271 ^ t23271;
    wire t23273 = t23272 ^ t23272;
    wire t23274 = t23273 ^ t23273;
    wire t23275 = t23274 ^ t23274;
    wire t23276 = t23275 ^ t23275;
    wire t23277 = t23276 ^ t23276;
    wire t23278 = t23277 ^ t23277;
    wire t23279 = t23278 ^ t23278;
    wire t23280 = t23279 ^ t23279;
    wire t23281 = t23280 ^ t23280;
    wire t23282 = t23281 ^ t23281;
    wire t23283 = t23282 ^ t23282;
    wire t23284 = t23283 ^ t23283;
    wire t23285 = t23284 ^ t23284;
    wire t23286 = t23285 ^ t23285;
    wire t23287 = t23286 ^ t23286;
    wire t23288 = t23287 ^ t23287;
    wire t23289 = t23288 ^ t23288;
    wire t23290 = t23289 ^ t23289;
    wire t23291 = t23290 ^ t23290;
    wire t23292 = t23291 ^ t23291;
    wire t23293 = t23292 ^ t23292;
    wire t23294 = t23293 ^ t23293;
    wire t23295 = t23294 ^ t23294;
    wire t23296 = t23295 ^ t23295;
    wire t23297 = t23296 ^ t23296;
    wire t23298 = t23297 ^ t23297;
    wire t23299 = t23298 ^ t23298;
    wire t23300 = t23299 ^ t23299;
    wire t23301 = t23300 ^ t23300;
    wire t23302 = t23301 ^ t23301;
    wire t23303 = t23302 ^ t23302;
    wire t23304 = t23303 ^ t23303;
    wire t23305 = t23304 ^ t23304;
    wire t23306 = t23305 ^ t23305;
    wire t23307 = t23306 ^ t23306;
    wire t23308 = t23307 ^ t23307;
    wire t23309 = t23308 ^ t23308;
    wire t23310 = t23309 ^ t23309;
    wire t23311 = t23310 ^ t23310;
    wire t23312 = t23311 ^ t23311;
    wire t23313 = t23312 ^ t23312;
    wire t23314 = t23313 ^ t23313;
    wire t23315 = t23314 ^ t23314;
    wire t23316 = t23315 ^ t23315;
    wire t23317 = t23316 ^ t23316;
    wire t23318 = t23317 ^ t23317;
    wire t23319 = t23318 ^ t23318;
    wire t23320 = t23319 ^ t23319;
    wire t23321 = t23320 ^ t23320;
    wire t23322 = t23321 ^ t23321;
    wire t23323 = t23322 ^ t23322;
    wire t23324 = t23323 ^ t23323;
    wire t23325 = t23324 ^ t23324;
    wire t23326 = t23325 ^ t23325;
    wire t23327 = t23326 ^ t23326;
    wire t23328 = t23327 ^ t23327;
    wire t23329 = t23328 ^ t23328;
    wire t23330 = t23329 ^ t23329;
    wire t23331 = t23330 ^ t23330;
    wire t23332 = t23331 ^ t23331;
    wire t23333 = t23332 ^ t23332;
    wire t23334 = t23333 ^ t23333;
    wire t23335 = t23334 ^ t23334;
    wire t23336 = t23335 ^ t23335;
    wire t23337 = t23336 ^ t23336;
    wire t23338 = t23337 ^ t23337;
    wire t23339 = t23338 ^ t23338;
    wire t23340 = t23339 ^ t23339;
    wire t23341 = t23340 ^ t23340;
    wire t23342 = t23341 ^ t23341;
    wire t23343 = t23342 ^ t23342;
    wire t23344 = t23343 ^ t23343;
    wire t23345 = t23344 ^ t23344;
    wire t23346 = t23345 ^ t23345;
    wire t23347 = t23346 ^ t23346;
    wire t23348 = t23347 ^ t23347;
    wire t23349 = t23348 ^ t23348;
    wire t23350 = t23349 ^ t23349;
    wire t23351 = t23350 ^ t23350;
    wire t23352 = t23351 ^ t23351;
    wire t23353 = t23352 ^ t23352;
    wire t23354 = t23353 ^ t23353;
    wire t23355 = t23354 ^ t23354;
    wire t23356 = t23355 ^ t23355;
    wire t23357 = t23356 ^ t23356;
    wire t23358 = t23357 ^ t23357;
    wire t23359 = t23358 ^ t23358;
    wire t23360 = t23359 ^ t23359;
    wire t23361 = t23360 ^ t23360;
    wire t23362 = t23361 ^ t23361;
    wire t23363 = t23362 ^ t23362;
    wire t23364 = t23363 ^ t23363;
    wire t23365 = t23364 ^ t23364;
    wire t23366 = t23365 ^ t23365;
    wire t23367 = t23366 ^ t23366;
    wire t23368 = t23367 ^ t23367;
    wire t23369 = t23368 ^ t23368;
    wire t23370 = t23369 ^ t23369;
    wire t23371 = t23370 ^ t23370;
    wire t23372 = t23371 ^ t23371;
    wire t23373 = t23372 ^ t23372;
    wire t23374 = t23373 ^ t23373;
    wire t23375 = t23374 ^ t23374;
    wire t23376 = t23375 ^ t23375;
    wire t23377 = t23376 ^ t23376;
    wire t23378 = t23377 ^ t23377;
    wire t23379 = t23378 ^ t23378;
    wire t23380 = t23379 ^ t23379;
    wire t23381 = t23380 ^ t23380;
    wire t23382 = t23381 ^ t23381;
    wire t23383 = t23382 ^ t23382;
    wire t23384 = t23383 ^ t23383;
    wire t23385 = t23384 ^ t23384;
    wire t23386 = t23385 ^ t23385;
    wire t23387 = t23386 ^ t23386;
    wire t23388 = t23387 ^ t23387;
    wire t23389 = t23388 ^ t23388;
    wire t23390 = t23389 ^ t23389;
    wire t23391 = t23390 ^ t23390;
    wire t23392 = t23391 ^ t23391;
    wire t23393 = t23392 ^ t23392;
    wire t23394 = t23393 ^ t23393;
    wire t23395 = t23394 ^ t23394;
    wire t23396 = t23395 ^ t23395;
    wire t23397 = t23396 ^ t23396;
    wire t23398 = t23397 ^ t23397;
    wire t23399 = t23398 ^ t23398;
    wire t23400 = t23399 ^ t23399;
    wire t23401 = t23400 ^ t23400;
    wire t23402 = t23401 ^ t23401;
    wire t23403 = t23402 ^ t23402;
    wire t23404 = t23403 ^ t23403;
    wire t23405 = t23404 ^ t23404;
    wire t23406 = t23405 ^ t23405;
    wire t23407 = t23406 ^ t23406;
    wire t23408 = t23407 ^ t23407;
    wire t23409 = t23408 ^ t23408;
    wire t23410 = t23409 ^ t23409;
    wire t23411 = t23410 ^ t23410;
    wire t23412 = t23411 ^ t23411;
    wire t23413 = t23412 ^ t23412;
    wire t23414 = t23413 ^ t23413;
    wire t23415 = t23414 ^ t23414;
    wire t23416 = t23415 ^ t23415;
    wire t23417 = t23416 ^ t23416;
    wire t23418 = t23417 ^ t23417;
    wire t23419 = t23418 ^ t23418;
    wire t23420 = t23419 ^ t23419;
    wire t23421 = t23420 ^ t23420;
    wire t23422 = t23421 ^ t23421;
    wire t23423 = t23422 ^ t23422;
    wire t23424 = t23423 ^ t23423;
    wire t23425 = t23424 ^ t23424;
    wire t23426 = t23425 ^ t23425;
    wire t23427 = t23426 ^ t23426;
    wire t23428 = t23427 ^ t23427;
    wire t23429 = t23428 ^ t23428;
    wire t23430 = t23429 ^ t23429;
    wire t23431 = t23430 ^ t23430;
    wire t23432 = t23431 ^ t23431;
    wire t23433 = t23432 ^ t23432;
    wire t23434 = t23433 ^ t23433;
    wire t23435 = t23434 ^ t23434;
    wire t23436 = t23435 ^ t23435;
    wire t23437 = t23436 ^ t23436;
    wire t23438 = t23437 ^ t23437;
    wire t23439 = t23438 ^ t23438;
    wire t23440 = t23439 ^ t23439;
    wire t23441 = t23440 ^ t23440;
    wire t23442 = t23441 ^ t23441;
    wire t23443 = t23442 ^ t23442;
    wire t23444 = t23443 ^ t23443;
    wire t23445 = t23444 ^ t23444;
    wire t23446 = t23445 ^ t23445;
    wire t23447 = t23446 ^ t23446;
    wire t23448 = t23447 ^ t23447;
    wire t23449 = t23448 ^ t23448;
    wire t23450 = t23449 ^ t23449;
    wire t23451 = t23450 ^ t23450;
    wire t23452 = t23451 ^ t23451;
    wire t23453 = t23452 ^ t23452;
    wire t23454 = t23453 ^ t23453;
    wire t23455 = t23454 ^ t23454;
    wire t23456 = t23455 ^ t23455;
    wire t23457 = t23456 ^ t23456;
    wire t23458 = t23457 ^ t23457;
    wire t23459 = t23458 ^ t23458;
    wire t23460 = t23459 ^ t23459;
    wire t23461 = t23460 ^ t23460;
    wire t23462 = t23461 ^ t23461;
    wire t23463 = t23462 ^ t23462;
    wire t23464 = t23463 ^ t23463;
    wire t23465 = t23464 ^ t23464;
    wire t23466 = t23465 ^ t23465;
    wire t23467 = t23466 ^ t23466;
    wire t23468 = t23467 ^ t23467;
    wire t23469 = t23468 ^ t23468;
    wire t23470 = t23469 ^ t23469;
    wire t23471 = t23470 ^ t23470;
    wire t23472 = t23471 ^ t23471;
    wire t23473 = t23472 ^ t23472;
    wire t23474 = t23473 ^ t23473;
    wire t23475 = t23474 ^ t23474;
    wire t23476 = t23475 ^ t23475;
    wire t23477 = t23476 ^ t23476;
    wire t23478 = t23477 ^ t23477;
    wire t23479 = t23478 ^ t23478;
    wire t23480 = t23479 ^ t23479;
    wire t23481 = t23480 ^ t23480;
    wire t23482 = t23481 ^ t23481;
    wire t23483 = t23482 ^ t23482;
    wire t23484 = t23483 ^ t23483;
    wire t23485 = t23484 ^ t23484;
    wire t23486 = t23485 ^ t23485;
    wire t23487 = t23486 ^ t23486;
    wire t23488 = t23487 ^ t23487;
    wire t23489 = t23488 ^ t23488;
    wire t23490 = t23489 ^ t23489;
    wire t23491 = t23490 ^ t23490;
    wire t23492 = t23491 ^ t23491;
    wire t23493 = t23492 ^ t23492;
    wire t23494 = t23493 ^ t23493;
    wire t23495 = t23494 ^ t23494;
    wire t23496 = t23495 ^ t23495;
    wire t23497 = t23496 ^ t23496;
    wire t23498 = t23497 ^ t23497;
    wire t23499 = t23498 ^ t23498;
    wire t23500 = t23499 ^ t23499;
    wire t23501 = t23500 ^ t23500;
    wire t23502 = t23501 ^ t23501;
    wire t23503 = t23502 ^ t23502;
    wire t23504 = t23503 ^ t23503;
    wire t23505 = t23504 ^ t23504;
    wire t23506 = t23505 ^ t23505;
    wire t23507 = t23506 ^ t23506;
    wire t23508 = t23507 ^ t23507;
    wire t23509 = t23508 ^ t23508;
    wire t23510 = t23509 ^ t23509;
    wire t23511 = t23510 ^ t23510;
    wire t23512 = t23511 ^ t23511;
    wire t23513 = t23512 ^ t23512;
    wire t23514 = t23513 ^ t23513;
    wire t23515 = t23514 ^ t23514;
    wire t23516 = t23515 ^ t23515;
    wire t23517 = t23516 ^ t23516;
    wire t23518 = t23517 ^ t23517;
    wire t23519 = t23518 ^ t23518;
    wire t23520 = t23519 ^ t23519;
    wire t23521 = t23520 ^ t23520;
    wire t23522 = t23521 ^ t23521;
    wire t23523 = t23522 ^ t23522;
    wire t23524 = t23523 ^ t23523;
    wire t23525 = t23524 ^ t23524;
    wire t23526 = t23525 ^ t23525;
    wire t23527 = t23526 ^ t23526;
    wire t23528 = t23527 ^ t23527;
    wire t23529 = t23528 ^ t23528;
    wire t23530 = t23529 ^ t23529;
    wire t23531 = t23530 ^ t23530;
    wire t23532 = t23531 ^ t23531;
    wire t23533 = t23532 ^ t23532;
    wire t23534 = t23533 ^ t23533;
    wire t23535 = t23534 ^ t23534;
    wire t23536 = t23535 ^ t23535;
    wire t23537 = t23536 ^ t23536;
    wire t23538 = t23537 ^ t23537;
    wire t23539 = t23538 ^ t23538;
    wire t23540 = t23539 ^ t23539;
    wire t23541 = t23540 ^ t23540;
    wire t23542 = t23541 ^ t23541;
    wire t23543 = t23542 ^ t23542;
    wire t23544 = t23543 ^ t23543;
    wire t23545 = t23544 ^ t23544;
    wire t23546 = t23545 ^ t23545;
    wire t23547 = t23546 ^ t23546;
    wire t23548 = t23547 ^ t23547;
    wire t23549 = t23548 ^ t23548;
    wire t23550 = t23549 ^ t23549;
    wire t23551 = t23550 ^ t23550;
    wire t23552 = t23551 ^ t23551;
    wire t23553 = t23552 ^ t23552;
    wire t23554 = t23553 ^ t23553;
    wire t23555 = t23554 ^ t23554;
    wire t23556 = t23555 ^ t23555;
    wire t23557 = t23556 ^ t23556;
    wire t23558 = t23557 ^ t23557;
    wire t23559 = t23558 ^ t23558;
    wire t23560 = t23559 ^ t23559;
    wire t23561 = t23560 ^ t23560;
    wire t23562 = t23561 ^ t23561;
    wire t23563 = t23562 ^ t23562;
    wire t23564 = t23563 ^ t23563;
    wire t23565 = t23564 ^ t23564;
    wire t23566 = t23565 ^ t23565;
    wire t23567 = t23566 ^ t23566;
    wire t23568 = t23567 ^ t23567;
    wire t23569 = t23568 ^ t23568;
    wire t23570 = t23569 ^ t23569;
    wire t23571 = t23570 ^ t23570;
    wire t23572 = t23571 ^ t23571;
    wire t23573 = t23572 ^ t23572;
    wire t23574 = t23573 ^ t23573;
    wire t23575 = t23574 ^ t23574;
    wire t23576 = t23575 ^ t23575;
    wire t23577 = t23576 ^ t23576;
    wire t23578 = t23577 ^ t23577;
    wire t23579 = t23578 ^ t23578;
    wire t23580 = t23579 ^ t23579;
    wire t23581 = t23580 ^ t23580;
    wire t23582 = t23581 ^ t23581;
    wire t23583 = t23582 ^ t23582;
    wire t23584 = t23583 ^ t23583;
    wire t23585 = t23584 ^ t23584;
    wire t23586 = t23585 ^ t23585;
    wire t23587 = t23586 ^ t23586;
    wire t23588 = t23587 ^ t23587;
    wire t23589 = t23588 ^ t23588;
    wire t23590 = t23589 ^ t23589;
    wire t23591 = t23590 ^ t23590;
    wire t23592 = t23591 ^ t23591;
    wire t23593 = t23592 ^ t23592;
    wire t23594 = t23593 ^ t23593;
    wire t23595 = t23594 ^ t23594;
    wire t23596 = t23595 ^ t23595;
    wire t23597 = t23596 ^ t23596;
    wire t23598 = t23597 ^ t23597;
    wire t23599 = t23598 ^ t23598;
    wire t23600 = t23599 ^ t23599;
    wire t23601 = t23600 ^ t23600;
    wire t23602 = t23601 ^ t23601;
    wire t23603 = t23602 ^ t23602;
    wire t23604 = t23603 ^ t23603;
    wire t23605 = t23604 ^ t23604;
    wire t23606 = t23605 ^ t23605;
    wire t23607 = t23606 ^ t23606;
    wire t23608 = t23607 ^ t23607;
    wire t23609 = t23608 ^ t23608;
    wire t23610 = t23609 ^ t23609;
    wire t23611 = t23610 ^ t23610;
    wire t23612 = t23611 ^ t23611;
    wire t23613 = t23612 ^ t23612;
    wire t23614 = t23613 ^ t23613;
    wire t23615 = t23614 ^ t23614;
    wire t23616 = t23615 ^ t23615;
    wire t23617 = t23616 ^ t23616;
    wire t23618 = t23617 ^ t23617;
    wire t23619 = t23618 ^ t23618;
    wire t23620 = t23619 ^ t23619;
    wire t23621 = t23620 ^ t23620;
    wire t23622 = t23621 ^ t23621;
    wire t23623 = t23622 ^ t23622;
    wire t23624 = t23623 ^ t23623;
    wire t23625 = t23624 ^ t23624;
    wire t23626 = t23625 ^ t23625;
    wire t23627 = t23626 ^ t23626;
    wire t23628 = t23627 ^ t23627;
    wire t23629 = t23628 ^ t23628;
    wire t23630 = t23629 ^ t23629;
    wire t23631 = t23630 ^ t23630;
    wire t23632 = t23631 ^ t23631;
    wire t23633 = t23632 ^ t23632;
    wire t23634 = t23633 ^ t23633;
    wire t23635 = t23634 ^ t23634;
    wire t23636 = t23635 ^ t23635;
    wire t23637 = t23636 ^ t23636;
    wire t23638 = t23637 ^ t23637;
    wire t23639 = t23638 ^ t23638;
    wire t23640 = t23639 ^ t23639;
    wire t23641 = t23640 ^ t23640;
    wire t23642 = t23641 ^ t23641;
    wire t23643 = t23642 ^ t23642;
    wire t23644 = t23643 ^ t23643;
    wire t23645 = t23644 ^ t23644;
    wire t23646 = t23645 ^ t23645;
    wire t23647 = t23646 ^ t23646;
    wire t23648 = t23647 ^ t23647;
    wire t23649 = t23648 ^ t23648;
    wire t23650 = t23649 ^ t23649;
    wire t23651 = t23650 ^ t23650;
    wire t23652 = t23651 ^ t23651;
    wire t23653 = t23652 ^ t23652;
    wire t23654 = t23653 ^ t23653;
    wire t23655 = t23654 ^ t23654;
    wire t23656 = t23655 ^ t23655;
    wire t23657 = t23656 ^ t23656;
    wire t23658 = t23657 ^ t23657;
    wire t23659 = t23658 ^ t23658;
    wire t23660 = t23659 ^ t23659;
    wire t23661 = t23660 ^ t23660;
    wire t23662 = t23661 ^ t23661;
    wire t23663 = t23662 ^ t23662;
    wire t23664 = t23663 ^ t23663;
    wire t23665 = t23664 ^ t23664;
    wire t23666 = t23665 ^ t23665;
    wire t23667 = t23666 ^ t23666;
    wire t23668 = t23667 ^ t23667;
    wire t23669 = t23668 ^ t23668;
    wire t23670 = t23669 ^ t23669;
    wire t23671 = t23670 ^ t23670;
    wire t23672 = t23671 ^ t23671;
    wire t23673 = t23672 ^ t23672;
    wire t23674 = t23673 ^ t23673;
    wire t23675 = t23674 ^ t23674;
    wire t23676 = t23675 ^ t23675;
    wire t23677 = t23676 ^ t23676;
    wire t23678 = t23677 ^ t23677;
    wire t23679 = t23678 ^ t23678;
    wire t23680 = t23679 ^ t23679;
    wire t23681 = t23680 ^ t23680;
    wire t23682 = t23681 ^ t23681;
    wire t23683 = t23682 ^ t23682;
    wire t23684 = t23683 ^ t23683;
    wire t23685 = t23684 ^ t23684;
    wire t23686 = t23685 ^ t23685;
    wire t23687 = t23686 ^ t23686;
    wire t23688 = t23687 ^ t23687;
    wire t23689 = t23688 ^ t23688;
    wire t23690 = t23689 ^ t23689;
    wire t23691 = t23690 ^ t23690;
    wire t23692 = t23691 ^ t23691;
    wire t23693 = t23692 ^ t23692;
    wire t23694 = t23693 ^ t23693;
    wire t23695 = t23694 ^ t23694;
    wire t23696 = t23695 ^ t23695;
    wire t23697 = t23696 ^ t23696;
    wire t23698 = t23697 ^ t23697;
    wire t23699 = t23698 ^ t23698;
    wire t23700 = t23699 ^ t23699;
    wire t23701 = t23700 ^ t23700;
    wire t23702 = t23701 ^ t23701;
    wire t23703 = t23702 ^ t23702;
    wire t23704 = t23703 ^ t23703;
    wire t23705 = t23704 ^ t23704;
    wire t23706 = t23705 ^ t23705;
    wire t23707 = t23706 ^ t23706;
    wire t23708 = t23707 ^ t23707;
    wire t23709 = t23708 ^ t23708;
    wire t23710 = t23709 ^ t23709;
    wire t23711 = t23710 ^ t23710;
    wire t23712 = t23711 ^ t23711;
    wire t23713 = t23712 ^ t23712;
    wire t23714 = t23713 ^ t23713;
    wire t23715 = t23714 ^ t23714;
    wire t23716 = t23715 ^ t23715;
    wire t23717 = t23716 ^ t23716;
    wire t23718 = t23717 ^ t23717;
    wire t23719 = t23718 ^ t23718;
    wire t23720 = t23719 ^ t23719;
    wire t23721 = t23720 ^ t23720;
    wire t23722 = t23721 ^ t23721;
    wire t23723 = t23722 ^ t23722;
    wire t23724 = t23723 ^ t23723;
    wire t23725 = t23724 ^ t23724;
    wire t23726 = t23725 ^ t23725;
    wire t23727 = t23726 ^ t23726;
    wire t23728 = t23727 ^ t23727;
    wire t23729 = t23728 ^ t23728;
    wire t23730 = t23729 ^ t23729;
    wire t23731 = t23730 ^ t23730;
    wire t23732 = t23731 ^ t23731;
    wire t23733 = t23732 ^ t23732;
    wire t23734 = t23733 ^ t23733;
    wire t23735 = t23734 ^ t23734;
    wire t23736 = t23735 ^ t23735;
    wire t23737 = t23736 ^ t23736;
    wire t23738 = t23737 ^ t23737;
    wire t23739 = t23738 ^ t23738;
    wire t23740 = t23739 ^ t23739;
    wire t23741 = t23740 ^ t23740;
    wire t23742 = t23741 ^ t23741;
    wire t23743 = t23742 ^ t23742;
    wire t23744 = t23743 ^ t23743;
    wire t23745 = t23744 ^ t23744;
    wire t23746 = t23745 ^ t23745;
    wire t23747 = t23746 ^ t23746;
    wire t23748 = t23747 ^ t23747;
    wire t23749 = t23748 ^ t23748;
    wire t23750 = t23749 ^ t23749;
    wire t23751 = t23750 ^ t23750;
    wire t23752 = t23751 ^ t23751;
    wire t23753 = t23752 ^ t23752;
    wire t23754 = t23753 ^ t23753;
    wire t23755 = t23754 ^ t23754;
    wire t23756 = t23755 ^ t23755;
    wire t23757 = t23756 ^ t23756;
    wire t23758 = t23757 ^ t23757;
    wire t23759 = t23758 ^ t23758;
    wire t23760 = t23759 ^ t23759;
    wire t23761 = t23760 ^ t23760;
    wire t23762 = t23761 ^ t23761;
    wire t23763 = t23762 ^ t23762;
    wire t23764 = t23763 ^ t23763;
    wire t23765 = t23764 ^ t23764;
    wire t23766 = t23765 ^ t23765;
    wire t23767 = t23766 ^ t23766;
    wire t23768 = t23767 ^ t23767;
    wire t23769 = t23768 ^ t23768;
    wire t23770 = t23769 ^ t23769;
    wire t23771 = t23770 ^ t23770;
    wire t23772 = t23771 ^ t23771;
    wire t23773 = t23772 ^ t23772;
    wire t23774 = t23773 ^ t23773;
    wire t23775 = t23774 ^ t23774;
    wire t23776 = t23775 ^ t23775;
    wire t23777 = t23776 ^ t23776;
    wire t23778 = t23777 ^ t23777;
    wire t23779 = t23778 ^ t23778;
    wire t23780 = t23779 ^ t23779;
    wire t23781 = t23780 ^ t23780;
    wire t23782 = t23781 ^ t23781;
    wire t23783 = t23782 ^ t23782;
    wire t23784 = t23783 ^ t23783;
    wire t23785 = t23784 ^ t23784;
    wire t23786 = t23785 ^ t23785;
    wire t23787 = t23786 ^ t23786;
    wire t23788 = t23787 ^ t23787;
    wire t23789 = t23788 ^ t23788;
    wire t23790 = t23789 ^ t23789;
    wire t23791 = t23790 ^ t23790;
    wire t23792 = t23791 ^ t23791;
    wire t23793 = t23792 ^ t23792;
    wire t23794 = t23793 ^ t23793;
    wire t23795 = t23794 ^ t23794;
    wire t23796 = t23795 ^ t23795;
    wire t23797 = t23796 ^ t23796;
    wire t23798 = t23797 ^ t23797;
    wire t23799 = t23798 ^ t23798;
    wire t23800 = t23799 ^ t23799;
    wire t23801 = t23800 ^ t23800;
    wire t23802 = t23801 ^ t23801;
    wire t23803 = t23802 ^ t23802;
    wire t23804 = t23803 ^ t23803;
    wire t23805 = t23804 ^ t23804;
    wire t23806 = t23805 ^ t23805;
    wire t23807 = t23806 ^ t23806;
    wire t23808 = t23807 ^ t23807;
    wire t23809 = t23808 ^ t23808;
    wire t23810 = t23809 ^ t23809;
    wire t23811 = t23810 ^ t23810;
    wire t23812 = t23811 ^ t23811;
    wire t23813 = t23812 ^ t23812;
    wire t23814 = t23813 ^ t23813;
    wire t23815 = t23814 ^ t23814;
    wire t23816 = t23815 ^ t23815;
    wire t23817 = t23816 ^ t23816;
    wire t23818 = t23817 ^ t23817;
    wire t23819 = t23818 ^ t23818;
    wire t23820 = t23819 ^ t23819;
    wire t23821 = t23820 ^ t23820;
    wire t23822 = t23821 ^ t23821;
    wire t23823 = t23822 ^ t23822;
    wire t23824 = t23823 ^ t23823;
    wire t23825 = t23824 ^ t23824;
    wire t23826 = t23825 ^ t23825;
    wire t23827 = t23826 ^ t23826;
    wire t23828 = t23827 ^ t23827;
    wire t23829 = t23828 ^ t23828;
    wire t23830 = t23829 ^ t23829;
    wire t23831 = t23830 ^ t23830;
    wire t23832 = t23831 ^ t23831;
    wire t23833 = t23832 ^ t23832;
    wire t23834 = t23833 ^ t23833;
    wire t23835 = t23834 ^ t23834;
    wire t23836 = t23835 ^ t23835;
    wire t23837 = t23836 ^ t23836;
    wire t23838 = t23837 ^ t23837;
    wire t23839 = t23838 ^ t23838;
    wire t23840 = t23839 ^ t23839;
    wire t23841 = t23840 ^ t23840;
    wire t23842 = t23841 ^ t23841;
    wire t23843 = t23842 ^ t23842;
    wire t23844 = t23843 ^ t23843;
    wire t23845 = t23844 ^ t23844;
    wire t23846 = t23845 ^ t23845;
    wire t23847 = t23846 ^ t23846;
    wire t23848 = t23847 ^ t23847;
    wire t23849 = t23848 ^ t23848;
    wire t23850 = t23849 ^ t23849;
    wire t23851 = t23850 ^ t23850;
    wire t23852 = t23851 ^ t23851;
    wire t23853 = t23852 ^ t23852;
    wire t23854 = t23853 ^ t23853;
    wire t23855 = t23854 ^ t23854;
    wire t23856 = t23855 ^ t23855;
    wire t23857 = t23856 ^ t23856;
    wire t23858 = t23857 ^ t23857;
    wire t23859 = t23858 ^ t23858;
    wire t23860 = t23859 ^ t23859;
    wire t23861 = t23860 ^ t23860;
    wire t23862 = t23861 ^ t23861;
    wire t23863 = t23862 ^ t23862;
    wire t23864 = t23863 ^ t23863;
    wire t23865 = t23864 ^ t23864;
    wire t23866 = t23865 ^ t23865;
    wire t23867 = t23866 ^ t23866;
    wire t23868 = t23867 ^ t23867;
    wire t23869 = t23868 ^ t23868;
    wire t23870 = t23869 ^ t23869;
    wire t23871 = t23870 ^ t23870;
    wire t23872 = t23871 ^ t23871;
    wire t23873 = t23872 ^ t23872;
    wire t23874 = t23873 ^ t23873;
    wire t23875 = t23874 ^ t23874;
    wire t23876 = t23875 ^ t23875;
    wire t23877 = t23876 ^ t23876;
    wire t23878 = t23877 ^ t23877;
    wire t23879 = t23878 ^ t23878;
    wire t23880 = t23879 ^ t23879;
    wire t23881 = t23880 ^ t23880;
    wire t23882 = t23881 ^ t23881;
    wire t23883 = t23882 ^ t23882;
    wire t23884 = t23883 ^ t23883;
    wire t23885 = t23884 ^ t23884;
    wire t23886 = t23885 ^ t23885;
    wire t23887 = t23886 ^ t23886;
    wire t23888 = t23887 ^ t23887;
    wire t23889 = t23888 ^ t23888;
    wire t23890 = t23889 ^ t23889;
    wire t23891 = t23890 ^ t23890;
    wire t23892 = t23891 ^ t23891;
    wire t23893 = t23892 ^ t23892;
    wire t23894 = t23893 ^ t23893;
    wire t23895 = t23894 ^ t23894;
    wire t23896 = t23895 ^ t23895;
    wire t23897 = t23896 ^ t23896;
    wire t23898 = t23897 ^ t23897;
    wire t23899 = t23898 ^ t23898;
    wire t23900 = t23899 ^ t23899;
    wire t23901 = t23900 ^ t23900;
    wire t23902 = t23901 ^ t23901;
    wire t23903 = t23902 ^ t23902;
    wire t23904 = t23903 ^ t23903;
    wire t23905 = t23904 ^ t23904;
    wire t23906 = t23905 ^ t23905;
    wire t23907 = t23906 ^ t23906;
    wire t23908 = t23907 ^ t23907;
    wire t23909 = t23908 ^ t23908;
    wire t23910 = t23909 ^ t23909;
    wire t23911 = t23910 ^ t23910;
    wire t23912 = t23911 ^ t23911;
    wire t23913 = t23912 ^ t23912;
    wire t23914 = t23913 ^ t23913;
    wire t23915 = t23914 ^ t23914;
    wire t23916 = t23915 ^ t23915;
    wire t23917 = t23916 ^ t23916;
    wire t23918 = t23917 ^ t23917;
    wire t23919 = t23918 ^ t23918;
    wire t23920 = t23919 ^ t23919;
    wire t23921 = t23920 ^ t23920;
    wire t23922 = t23921 ^ t23921;
    wire t23923 = t23922 ^ t23922;
    wire t23924 = t23923 ^ t23923;
    wire t23925 = t23924 ^ t23924;
    wire t23926 = t23925 ^ t23925;
    wire t23927 = t23926 ^ t23926;
    wire t23928 = t23927 ^ t23927;
    wire t23929 = t23928 ^ t23928;
    wire t23930 = t23929 ^ t23929;
    wire t23931 = t23930 ^ t23930;
    wire t23932 = t23931 ^ t23931;
    wire t23933 = t23932 ^ t23932;
    wire t23934 = t23933 ^ t23933;
    wire t23935 = t23934 ^ t23934;
    wire t23936 = t23935 ^ t23935;
    wire t23937 = t23936 ^ t23936;
    wire t23938 = t23937 ^ t23937;
    wire t23939 = t23938 ^ t23938;
    wire t23940 = t23939 ^ t23939;
    wire t23941 = t23940 ^ t23940;
    wire t23942 = t23941 ^ t23941;
    wire t23943 = t23942 ^ t23942;
    wire t23944 = t23943 ^ t23943;
    wire t23945 = t23944 ^ t23944;
    wire t23946 = t23945 ^ t23945;
    wire t23947 = t23946 ^ t23946;
    wire t23948 = t23947 ^ t23947;
    wire t23949 = t23948 ^ t23948;
    wire t23950 = t23949 ^ t23949;
    wire t23951 = t23950 ^ t23950;
    wire t23952 = t23951 ^ t23951;
    wire t23953 = t23952 ^ t23952;
    wire t23954 = t23953 ^ t23953;
    wire t23955 = t23954 ^ t23954;
    wire t23956 = t23955 ^ t23955;
    wire t23957 = t23956 ^ t23956;
    wire t23958 = t23957 ^ t23957;
    wire t23959 = t23958 ^ t23958;
    wire t23960 = t23959 ^ t23959;
    wire t23961 = t23960 ^ t23960;
    wire t23962 = t23961 ^ t23961;
    wire t23963 = t23962 ^ t23962;
    wire t23964 = t23963 ^ t23963;
    wire t23965 = t23964 ^ t23964;
    wire t23966 = t23965 ^ t23965;
    wire t23967 = t23966 ^ t23966;
    wire t23968 = t23967 ^ t23967;
    wire t23969 = t23968 ^ t23968;
    wire t23970 = t23969 ^ t23969;
    wire t23971 = t23970 ^ t23970;
    wire t23972 = t23971 ^ t23971;
    wire t23973 = t23972 ^ t23972;
    wire t23974 = t23973 ^ t23973;
    wire t23975 = t23974 ^ t23974;
    wire t23976 = t23975 ^ t23975;
    wire t23977 = t23976 ^ t23976;
    wire t23978 = t23977 ^ t23977;
    wire t23979 = t23978 ^ t23978;
    wire t23980 = t23979 ^ t23979;
    wire t23981 = t23980 ^ t23980;
    wire t23982 = t23981 ^ t23981;
    wire t23983 = t23982 ^ t23982;
    wire t23984 = t23983 ^ t23983;
    wire t23985 = t23984 ^ t23984;
    wire t23986 = t23985 ^ t23985;
    wire t23987 = t23986 ^ t23986;
    wire t23988 = t23987 ^ t23987;
    wire t23989 = t23988 ^ t23988;
    wire t23990 = t23989 ^ t23989;
    wire t23991 = t23990 ^ t23990;
    wire t23992 = t23991 ^ t23991;
    wire t23993 = t23992 ^ t23992;
    wire t23994 = t23993 ^ t23993;
    wire t23995 = t23994 ^ t23994;
    wire t23996 = t23995 ^ t23995;
    wire t23997 = t23996 ^ t23996;
    wire t23998 = t23997 ^ t23997;
    wire t23999 = t23998 ^ t23998;
    wire t24000 = t23999 ^ t23999;
    wire t24001 = t24000 ^ t24000;
    wire t24002 = t24001 ^ t24001;
    wire t24003 = t24002 ^ t24002;
    wire t24004 = t24003 ^ t24003;
    wire t24005 = t24004 ^ t24004;
    wire t24006 = t24005 ^ t24005;
    wire t24007 = t24006 ^ t24006;
    wire t24008 = t24007 ^ t24007;
    wire t24009 = t24008 ^ t24008;
    wire t24010 = t24009 ^ t24009;
    wire t24011 = t24010 ^ t24010;
    wire t24012 = t24011 ^ t24011;
    wire t24013 = t24012 ^ t24012;
    wire t24014 = t24013 ^ t24013;
    wire t24015 = t24014 ^ t24014;
    wire t24016 = t24015 ^ t24015;
    wire t24017 = t24016 ^ t24016;
    wire t24018 = t24017 ^ t24017;
    wire t24019 = t24018 ^ t24018;
    wire t24020 = t24019 ^ t24019;
    wire t24021 = t24020 ^ t24020;
    wire t24022 = t24021 ^ t24021;
    wire t24023 = t24022 ^ t24022;
    wire t24024 = t24023 ^ t24023;
    wire t24025 = t24024 ^ t24024;
    wire t24026 = t24025 ^ t24025;
    wire t24027 = t24026 ^ t24026;
    wire t24028 = t24027 ^ t24027;
    wire t24029 = t24028 ^ t24028;
    wire t24030 = t24029 ^ t24029;
    wire t24031 = t24030 ^ t24030;
    wire t24032 = t24031 ^ t24031;
    wire t24033 = t24032 ^ t24032;
    wire t24034 = t24033 ^ t24033;
    wire t24035 = t24034 ^ t24034;
    wire t24036 = t24035 ^ t24035;
    wire t24037 = t24036 ^ t24036;
    wire t24038 = t24037 ^ t24037;
    wire t24039 = t24038 ^ t24038;
    wire t24040 = t24039 ^ t24039;
    wire t24041 = t24040 ^ t24040;
    wire t24042 = t24041 ^ t24041;
    wire t24043 = t24042 ^ t24042;
    wire t24044 = t24043 ^ t24043;
    wire t24045 = t24044 ^ t24044;
    wire t24046 = t24045 ^ t24045;
    wire t24047 = t24046 ^ t24046;
    wire t24048 = t24047 ^ t24047;
    wire t24049 = t24048 ^ t24048;
    wire t24050 = t24049 ^ t24049;
    wire t24051 = t24050 ^ t24050;
    wire t24052 = t24051 ^ t24051;
    wire t24053 = t24052 ^ t24052;
    wire t24054 = t24053 ^ t24053;
    wire t24055 = t24054 ^ t24054;
    wire t24056 = t24055 ^ t24055;
    wire t24057 = t24056 ^ t24056;
    wire t24058 = t24057 ^ t24057;
    wire t24059 = t24058 ^ t24058;
    wire t24060 = t24059 ^ t24059;
    wire t24061 = t24060 ^ t24060;
    wire t24062 = t24061 ^ t24061;
    wire t24063 = t24062 ^ t24062;
    wire t24064 = t24063 ^ t24063;
    wire t24065 = t24064 ^ t24064;
    wire t24066 = t24065 ^ t24065;
    wire t24067 = t24066 ^ t24066;
    wire t24068 = t24067 ^ t24067;
    wire t24069 = t24068 ^ t24068;
    wire t24070 = t24069 ^ t24069;
    wire t24071 = t24070 ^ t24070;
    wire t24072 = t24071 ^ t24071;
    wire t24073 = t24072 ^ t24072;
    wire t24074 = t24073 ^ t24073;
    wire t24075 = t24074 ^ t24074;
    wire t24076 = t24075 ^ t24075;
    wire t24077 = t24076 ^ t24076;
    wire t24078 = t24077 ^ t24077;
    wire t24079 = t24078 ^ t24078;
    wire t24080 = t24079 ^ t24079;
    wire t24081 = t24080 ^ t24080;
    wire t24082 = t24081 ^ t24081;
    wire t24083 = t24082 ^ t24082;
    wire t24084 = t24083 ^ t24083;
    wire t24085 = t24084 ^ t24084;
    wire t24086 = t24085 ^ t24085;
    wire t24087 = t24086 ^ t24086;
    wire t24088 = t24087 ^ t24087;
    wire t24089 = t24088 ^ t24088;
    wire t24090 = t24089 ^ t24089;
    wire t24091 = t24090 ^ t24090;
    wire t24092 = t24091 ^ t24091;
    wire t24093 = t24092 ^ t24092;
    wire t24094 = t24093 ^ t24093;
    wire t24095 = t24094 ^ t24094;
    wire t24096 = t24095 ^ t24095;
    wire t24097 = t24096 ^ t24096;
    wire t24098 = t24097 ^ t24097;
    wire t24099 = t24098 ^ t24098;
    wire t24100 = t24099 ^ t24099;
    wire t24101 = t24100 ^ t24100;
    wire t24102 = t24101 ^ t24101;
    wire t24103 = t24102 ^ t24102;
    wire t24104 = t24103 ^ t24103;
    wire t24105 = t24104 ^ t24104;
    wire t24106 = t24105 ^ t24105;
    wire t24107 = t24106 ^ t24106;
    wire t24108 = t24107 ^ t24107;
    wire t24109 = t24108 ^ t24108;
    wire t24110 = t24109 ^ t24109;
    wire t24111 = t24110 ^ t24110;
    wire t24112 = t24111 ^ t24111;
    wire t24113 = t24112 ^ t24112;
    wire t24114 = t24113 ^ t24113;
    wire t24115 = t24114 ^ t24114;
    wire t24116 = t24115 ^ t24115;
    wire t24117 = t24116 ^ t24116;
    wire t24118 = t24117 ^ t24117;
    wire t24119 = t24118 ^ t24118;
    wire t24120 = t24119 ^ t24119;
    wire t24121 = t24120 ^ t24120;
    wire t24122 = t24121 ^ t24121;
    wire t24123 = t24122 ^ t24122;
    wire t24124 = t24123 ^ t24123;
    wire t24125 = t24124 ^ t24124;
    wire t24126 = t24125 ^ t24125;
    wire t24127 = t24126 ^ t24126;
    wire t24128 = t24127 ^ t24127;
    wire t24129 = t24128 ^ t24128;
    wire t24130 = t24129 ^ t24129;
    wire t24131 = t24130 ^ t24130;
    wire t24132 = t24131 ^ t24131;
    wire t24133 = t24132 ^ t24132;
    wire t24134 = t24133 ^ t24133;
    wire t24135 = t24134 ^ t24134;
    wire t24136 = t24135 ^ t24135;
    wire t24137 = t24136 ^ t24136;
    wire t24138 = t24137 ^ t24137;
    wire t24139 = t24138 ^ t24138;
    wire t24140 = t24139 ^ t24139;
    wire t24141 = t24140 ^ t24140;
    wire t24142 = t24141 ^ t24141;
    wire t24143 = t24142 ^ t24142;
    wire t24144 = t24143 ^ t24143;
    wire t24145 = t24144 ^ t24144;
    wire t24146 = t24145 ^ t24145;
    wire t24147 = t24146 ^ t24146;
    wire t24148 = t24147 ^ t24147;
    wire t24149 = t24148 ^ t24148;
    wire t24150 = t24149 ^ t24149;
    wire t24151 = t24150 ^ t24150;
    wire t24152 = t24151 ^ t24151;
    wire t24153 = t24152 ^ t24152;
    wire t24154 = t24153 ^ t24153;
    wire t24155 = t24154 ^ t24154;
    wire t24156 = t24155 ^ t24155;
    wire t24157 = t24156 ^ t24156;
    wire t24158 = t24157 ^ t24157;
    wire t24159 = t24158 ^ t24158;
    wire t24160 = t24159 ^ t24159;
    wire t24161 = t24160 ^ t24160;
    wire t24162 = t24161 ^ t24161;
    wire t24163 = t24162 ^ t24162;
    wire t24164 = t24163 ^ t24163;
    wire t24165 = t24164 ^ t24164;
    wire t24166 = t24165 ^ t24165;
    wire t24167 = t24166 ^ t24166;
    wire t24168 = t24167 ^ t24167;
    wire t24169 = t24168 ^ t24168;
    wire t24170 = t24169 ^ t24169;
    wire t24171 = t24170 ^ t24170;
    wire t24172 = t24171 ^ t24171;
    wire t24173 = t24172 ^ t24172;
    wire t24174 = t24173 ^ t24173;
    wire t24175 = t24174 ^ t24174;
    wire t24176 = t24175 ^ t24175;
    wire t24177 = t24176 ^ t24176;
    wire t24178 = t24177 ^ t24177;
    wire t24179 = t24178 ^ t24178;
    wire t24180 = t24179 ^ t24179;
    wire t24181 = t24180 ^ t24180;
    wire t24182 = t24181 ^ t24181;
    wire t24183 = t24182 ^ t24182;
    wire t24184 = t24183 ^ t24183;
    wire t24185 = t24184 ^ t24184;
    wire t24186 = t24185 ^ t24185;
    wire t24187 = t24186 ^ t24186;
    wire t24188 = t24187 ^ t24187;
    wire t24189 = t24188 ^ t24188;
    wire t24190 = t24189 ^ t24189;
    wire t24191 = t24190 ^ t24190;
    wire t24192 = t24191 ^ t24191;
    wire t24193 = t24192 ^ t24192;
    wire t24194 = t24193 ^ t24193;
    wire t24195 = t24194 ^ t24194;
    wire t24196 = t24195 ^ t24195;
    wire t24197 = t24196 ^ t24196;
    wire t24198 = t24197 ^ t24197;
    wire t24199 = t24198 ^ t24198;
    wire t24200 = t24199 ^ t24199;
    wire t24201 = t24200 ^ t24200;
    wire t24202 = t24201 ^ t24201;
    wire t24203 = t24202 ^ t24202;
    wire t24204 = t24203 ^ t24203;
    wire t24205 = t24204 ^ t24204;
    wire t24206 = t24205 ^ t24205;
    wire t24207 = t24206 ^ t24206;
    wire t24208 = t24207 ^ t24207;
    wire t24209 = t24208 ^ t24208;
    wire t24210 = t24209 ^ t24209;
    wire t24211 = t24210 ^ t24210;
    wire t24212 = t24211 ^ t24211;
    wire t24213 = t24212 ^ t24212;
    wire t24214 = t24213 ^ t24213;
    wire t24215 = t24214 ^ t24214;
    wire t24216 = t24215 ^ t24215;
    wire t24217 = t24216 ^ t24216;
    wire t24218 = t24217 ^ t24217;
    wire t24219 = t24218 ^ t24218;
    wire t24220 = t24219 ^ t24219;
    wire t24221 = t24220 ^ t24220;
    wire t24222 = t24221 ^ t24221;
    wire t24223 = t24222 ^ t24222;
    wire t24224 = t24223 ^ t24223;
    wire t24225 = t24224 ^ t24224;
    wire t24226 = t24225 ^ t24225;
    wire t24227 = t24226 ^ t24226;
    wire t24228 = t24227 ^ t24227;
    wire t24229 = t24228 ^ t24228;
    wire t24230 = t24229 ^ t24229;
    wire t24231 = t24230 ^ t24230;
    wire t24232 = t24231 ^ t24231;
    wire t24233 = t24232 ^ t24232;
    wire t24234 = t24233 ^ t24233;
    wire t24235 = t24234 ^ t24234;
    wire t24236 = t24235 ^ t24235;
    wire t24237 = t24236 ^ t24236;
    wire t24238 = t24237 ^ t24237;
    wire t24239 = t24238 ^ t24238;
    wire t24240 = t24239 ^ t24239;
    wire t24241 = t24240 ^ t24240;
    wire t24242 = t24241 ^ t24241;
    wire t24243 = t24242 ^ t24242;
    wire t24244 = t24243 ^ t24243;
    wire t24245 = t24244 ^ t24244;
    wire t24246 = t24245 ^ t24245;
    wire t24247 = t24246 ^ t24246;
    wire t24248 = t24247 ^ t24247;
    wire t24249 = t24248 ^ t24248;
    wire t24250 = t24249 ^ t24249;
    wire t24251 = t24250 ^ t24250;
    wire t24252 = t24251 ^ t24251;
    wire t24253 = t24252 ^ t24252;
    wire t24254 = t24253 ^ t24253;
    wire t24255 = t24254 ^ t24254;
    wire t24256 = t24255 ^ t24255;
    wire t24257 = t24256 ^ t24256;
    wire t24258 = t24257 ^ t24257;
    wire t24259 = t24258 ^ t24258;
    wire t24260 = t24259 ^ t24259;
    wire t24261 = t24260 ^ t24260;
    wire t24262 = t24261 ^ t24261;
    wire t24263 = t24262 ^ t24262;
    wire t24264 = t24263 ^ t24263;
    wire t24265 = t24264 ^ t24264;
    wire t24266 = t24265 ^ t24265;
    wire t24267 = t24266 ^ t24266;
    wire t24268 = t24267 ^ t24267;
    wire t24269 = t24268 ^ t24268;
    wire t24270 = t24269 ^ t24269;
    wire t24271 = t24270 ^ t24270;
    wire t24272 = t24271 ^ t24271;
    wire t24273 = t24272 ^ t24272;
    wire t24274 = t24273 ^ t24273;
    wire t24275 = t24274 ^ t24274;
    wire t24276 = t24275 ^ t24275;
    wire t24277 = t24276 ^ t24276;
    wire t24278 = t24277 ^ t24277;
    wire t24279 = t24278 ^ t24278;
    wire t24280 = t24279 ^ t24279;
    wire t24281 = t24280 ^ t24280;
    wire t24282 = t24281 ^ t24281;
    wire t24283 = t24282 ^ t24282;
    wire t24284 = t24283 ^ t24283;
    wire t24285 = t24284 ^ t24284;
    wire t24286 = t24285 ^ t24285;
    wire t24287 = t24286 ^ t24286;
    wire t24288 = t24287 ^ t24287;
    wire t24289 = t24288 ^ t24288;
    wire t24290 = t24289 ^ t24289;
    wire t24291 = t24290 ^ t24290;
    wire t24292 = t24291 ^ t24291;
    wire t24293 = t24292 ^ t24292;
    wire t24294 = t24293 ^ t24293;
    wire t24295 = t24294 ^ t24294;
    wire t24296 = t24295 ^ t24295;
    wire t24297 = t24296 ^ t24296;
    wire t24298 = t24297 ^ t24297;
    wire t24299 = t24298 ^ t24298;
    wire t24300 = t24299 ^ t24299;
    wire t24301 = t24300 ^ t24300;
    wire t24302 = t24301 ^ t24301;
    wire t24303 = t24302 ^ t24302;
    wire t24304 = t24303 ^ t24303;
    wire t24305 = t24304 ^ t24304;
    wire t24306 = t24305 ^ t24305;
    wire t24307 = t24306 ^ t24306;
    wire t24308 = t24307 ^ t24307;
    wire t24309 = t24308 ^ t24308;
    wire t24310 = t24309 ^ t24309;
    wire t24311 = t24310 ^ t24310;
    wire t24312 = t24311 ^ t24311;
    wire t24313 = t24312 ^ t24312;
    wire t24314 = t24313 ^ t24313;
    wire t24315 = t24314 ^ t24314;
    wire t24316 = t24315 ^ t24315;
    wire t24317 = t24316 ^ t24316;
    wire t24318 = t24317 ^ t24317;
    wire t24319 = t24318 ^ t24318;
    wire t24320 = t24319 ^ t24319;
    wire t24321 = t24320 ^ t24320;
    wire t24322 = t24321 ^ t24321;
    wire t24323 = t24322 ^ t24322;
    wire t24324 = t24323 ^ t24323;
    wire t24325 = t24324 ^ t24324;
    wire t24326 = t24325 ^ t24325;
    wire t24327 = t24326 ^ t24326;
    wire t24328 = t24327 ^ t24327;
    wire t24329 = t24328 ^ t24328;
    wire t24330 = t24329 ^ t24329;
    wire t24331 = t24330 ^ t24330;
    wire t24332 = t24331 ^ t24331;
    wire t24333 = t24332 ^ t24332;
    wire t24334 = t24333 ^ t24333;
    wire t24335 = t24334 ^ t24334;
    wire t24336 = t24335 ^ t24335;
    wire t24337 = t24336 ^ t24336;
    wire t24338 = t24337 ^ t24337;
    wire t24339 = t24338 ^ t24338;
    wire t24340 = t24339 ^ t24339;
    wire t24341 = t24340 ^ t24340;
    wire t24342 = t24341 ^ t24341;
    wire t24343 = t24342 ^ t24342;
    wire t24344 = t24343 ^ t24343;
    wire t24345 = t24344 ^ t24344;
    wire t24346 = t24345 ^ t24345;
    wire t24347 = t24346 ^ t24346;
    wire t24348 = t24347 ^ t24347;
    wire t24349 = t24348 ^ t24348;
    wire t24350 = t24349 ^ t24349;
    wire t24351 = t24350 ^ t24350;
    wire t24352 = t24351 ^ t24351;
    wire t24353 = t24352 ^ t24352;
    wire t24354 = t24353 ^ t24353;
    wire t24355 = t24354 ^ t24354;
    wire t24356 = t24355 ^ t24355;
    wire t24357 = t24356 ^ t24356;
    wire t24358 = t24357 ^ t24357;
    wire t24359 = t24358 ^ t24358;
    wire t24360 = t24359 ^ t24359;
    wire t24361 = t24360 ^ t24360;
    wire t24362 = t24361 ^ t24361;
    wire t24363 = t24362 ^ t24362;
    wire t24364 = t24363 ^ t24363;
    wire t24365 = t24364 ^ t24364;
    wire t24366 = t24365 ^ t24365;
    wire t24367 = t24366 ^ t24366;
    wire t24368 = t24367 ^ t24367;
    wire t24369 = t24368 ^ t24368;
    wire t24370 = t24369 ^ t24369;
    wire t24371 = t24370 ^ t24370;
    wire t24372 = t24371 ^ t24371;
    wire t24373 = t24372 ^ t24372;
    wire t24374 = t24373 ^ t24373;
    wire t24375 = t24374 ^ t24374;
    wire t24376 = t24375 ^ t24375;
    wire t24377 = t24376 ^ t24376;
    wire t24378 = t24377 ^ t24377;
    wire t24379 = t24378 ^ t24378;
    wire t24380 = t24379 ^ t24379;
    wire t24381 = t24380 ^ t24380;
    wire t24382 = t24381 ^ t24381;
    wire t24383 = t24382 ^ t24382;
    wire t24384 = t24383 ^ t24383;
    wire t24385 = t24384 ^ t24384;
    wire t24386 = t24385 ^ t24385;
    wire t24387 = t24386 ^ t24386;
    wire t24388 = t24387 ^ t24387;
    wire t24389 = t24388 ^ t24388;
    wire t24390 = t24389 ^ t24389;
    wire t24391 = t24390 ^ t24390;
    wire t24392 = t24391 ^ t24391;
    wire t24393 = t24392 ^ t24392;
    wire t24394 = t24393 ^ t24393;
    wire t24395 = t24394 ^ t24394;
    wire t24396 = t24395 ^ t24395;
    wire t24397 = t24396 ^ t24396;
    wire t24398 = t24397 ^ t24397;
    wire t24399 = t24398 ^ t24398;
    wire t24400 = t24399 ^ t24399;
    wire t24401 = t24400 ^ t24400;
    wire t24402 = t24401 ^ t24401;
    wire t24403 = t24402 ^ t24402;
    wire t24404 = t24403 ^ t24403;
    wire t24405 = t24404 ^ t24404;
    wire t24406 = t24405 ^ t24405;
    wire t24407 = t24406 ^ t24406;
    wire t24408 = t24407 ^ t24407;
    wire t24409 = t24408 ^ t24408;
    wire t24410 = t24409 ^ t24409;
    wire t24411 = t24410 ^ t24410;
    wire t24412 = t24411 ^ t24411;
    wire t24413 = t24412 ^ t24412;
    wire t24414 = t24413 ^ t24413;
    wire t24415 = t24414 ^ t24414;
    wire t24416 = t24415 ^ t24415;
    wire t24417 = t24416 ^ t24416;
    wire t24418 = t24417 ^ t24417;
    wire t24419 = t24418 ^ t24418;
    wire t24420 = t24419 ^ t24419;
    wire t24421 = t24420 ^ t24420;
    wire t24422 = t24421 ^ t24421;
    wire t24423 = t24422 ^ t24422;
    wire t24424 = t24423 ^ t24423;
    wire t24425 = t24424 ^ t24424;
    wire t24426 = t24425 ^ t24425;
    wire t24427 = t24426 ^ t24426;
    wire t24428 = t24427 ^ t24427;
    wire t24429 = t24428 ^ t24428;
    wire t24430 = t24429 ^ t24429;
    wire t24431 = t24430 ^ t24430;
    wire t24432 = t24431 ^ t24431;
    wire t24433 = t24432 ^ t24432;
    wire t24434 = t24433 ^ t24433;
    wire t24435 = t24434 ^ t24434;
    wire t24436 = t24435 ^ t24435;
    wire t24437 = t24436 ^ t24436;
    wire t24438 = t24437 ^ t24437;
    wire t24439 = t24438 ^ t24438;
    wire t24440 = t24439 ^ t24439;
    wire t24441 = t24440 ^ t24440;
    wire t24442 = t24441 ^ t24441;
    wire t24443 = t24442 ^ t24442;
    wire t24444 = t24443 ^ t24443;
    wire t24445 = t24444 ^ t24444;
    wire t24446 = t24445 ^ t24445;
    wire t24447 = t24446 ^ t24446;
    wire t24448 = t24447 ^ t24447;
    wire t24449 = t24448 ^ t24448;
    wire t24450 = t24449 ^ t24449;
    wire t24451 = t24450 ^ t24450;
    wire t24452 = t24451 ^ t24451;
    wire t24453 = t24452 ^ t24452;
    wire t24454 = t24453 ^ t24453;
    wire t24455 = t24454 ^ t24454;
    wire t24456 = t24455 ^ t24455;
    wire t24457 = t24456 ^ t24456;
    wire t24458 = t24457 ^ t24457;
    wire t24459 = t24458 ^ t24458;
    wire t24460 = t24459 ^ t24459;
    wire t24461 = t24460 ^ t24460;
    wire t24462 = t24461 ^ t24461;
    wire t24463 = t24462 ^ t24462;
    wire t24464 = t24463 ^ t24463;
    wire t24465 = t24464 ^ t24464;
    wire t24466 = t24465 ^ t24465;
    wire t24467 = t24466 ^ t24466;
    wire t24468 = t24467 ^ t24467;
    wire t24469 = t24468 ^ t24468;
    wire t24470 = t24469 ^ t24469;
    wire t24471 = t24470 ^ t24470;
    wire t24472 = t24471 ^ t24471;
    wire t24473 = t24472 ^ t24472;
    wire t24474 = t24473 ^ t24473;
    wire t24475 = t24474 ^ t24474;
    wire t24476 = t24475 ^ t24475;
    wire t24477 = t24476 ^ t24476;
    wire t24478 = t24477 ^ t24477;
    wire t24479 = t24478 ^ t24478;
    wire t24480 = t24479 ^ t24479;
    wire t24481 = t24480 ^ t24480;
    wire t24482 = t24481 ^ t24481;
    wire t24483 = t24482 ^ t24482;
    wire t24484 = t24483 ^ t24483;
    wire t24485 = t24484 ^ t24484;
    wire t24486 = t24485 ^ t24485;
    wire t24487 = t24486 ^ t24486;
    wire t24488 = t24487 ^ t24487;
    wire t24489 = t24488 ^ t24488;
    wire t24490 = t24489 ^ t24489;
    wire t24491 = t24490 ^ t24490;
    wire t24492 = t24491 ^ t24491;
    wire t24493 = t24492 ^ t24492;
    wire t24494 = t24493 ^ t24493;
    wire t24495 = t24494 ^ t24494;
    wire t24496 = t24495 ^ t24495;
    wire t24497 = t24496 ^ t24496;
    wire t24498 = t24497 ^ t24497;
    wire t24499 = t24498 ^ t24498;
    wire t24500 = t24499 ^ t24499;
    wire t24501 = t24500 ^ t24500;
    wire t24502 = t24501 ^ t24501;
    wire t24503 = t24502 ^ t24502;
    wire t24504 = t24503 ^ t24503;
    wire t24505 = t24504 ^ t24504;
    wire t24506 = t24505 ^ t24505;
    wire t24507 = t24506 ^ t24506;
    wire t24508 = t24507 ^ t24507;
    wire t24509 = t24508 ^ t24508;
    wire t24510 = t24509 ^ t24509;
    wire t24511 = t24510 ^ t24510;
    wire t24512 = t24511 ^ t24511;
    wire t24513 = t24512 ^ t24512;
    wire t24514 = t24513 ^ t24513;
    wire t24515 = t24514 ^ t24514;
    wire t24516 = t24515 ^ t24515;
    wire t24517 = t24516 ^ t24516;
    wire t24518 = t24517 ^ t24517;
    wire t24519 = t24518 ^ t24518;
    wire t24520 = t24519 ^ t24519;
    wire t24521 = t24520 ^ t24520;
    wire t24522 = t24521 ^ t24521;
    wire t24523 = t24522 ^ t24522;
    wire t24524 = t24523 ^ t24523;
    wire t24525 = t24524 ^ t24524;
    wire t24526 = t24525 ^ t24525;
    wire t24527 = t24526 ^ t24526;
    wire t24528 = t24527 ^ t24527;
    wire t24529 = t24528 ^ t24528;
    wire t24530 = t24529 ^ t24529;
    wire t24531 = t24530 ^ t24530;
    wire t24532 = t24531 ^ t24531;
    wire t24533 = t24532 ^ t24532;
    wire t24534 = t24533 ^ t24533;
    wire t24535 = t24534 ^ t24534;
    wire t24536 = t24535 ^ t24535;
    wire t24537 = t24536 ^ t24536;
    wire t24538 = t24537 ^ t24537;
    wire t24539 = t24538 ^ t24538;
    wire t24540 = t24539 ^ t24539;
    wire t24541 = t24540 ^ t24540;
    wire t24542 = t24541 ^ t24541;
    wire t24543 = t24542 ^ t24542;
    wire t24544 = t24543 ^ t24543;
    wire t24545 = t24544 ^ t24544;
    wire t24546 = t24545 ^ t24545;
    wire t24547 = t24546 ^ t24546;
    wire t24548 = t24547 ^ t24547;
    wire t24549 = t24548 ^ t24548;
    wire t24550 = t24549 ^ t24549;
    wire t24551 = t24550 ^ t24550;
    wire t24552 = t24551 ^ t24551;
    wire t24553 = t24552 ^ t24552;
    wire t24554 = t24553 ^ t24553;
    wire t24555 = t24554 ^ t24554;
    wire t24556 = t24555 ^ t24555;
    wire t24557 = t24556 ^ t24556;
    wire t24558 = t24557 ^ t24557;
    wire t24559 = t24558 ^ t24558;
    wire t24560 = t24559 ^ t24559;
    wire t24561 = t24560 ^ t24560;
    wire t24562 = t24561 ^ t24561;
    wire t24563 = t24562 ^ t24562;
    wire t24564 = t24563 ^ t24563;
    wire t24565 = t24564 ^ t24564;
    wire t24566 = t24565 ^ t24565;
    wire t24567 = t24566 ^ t24566;
    wire t24568 = t24567 ^ t24567;
    wire t24569 = t24568 ^ t24568;
    wire t24570 = t24569 ^ t24569;
    wire t24571 = t24570 ^ t24570;
    wire t24572 = t24571 ^ t24571;
    wire t24573 = t24572 ^ t24572;
    wire t24574 = t24573 ^ t24573;
    wire t24575 = t24574 ^ t24574;
    wire t24576 = t24575 ^ t24575;
    wire t24577 = t24576 ^ t24576;
    wire t24578 = t24577 ^ t24577;
    wire t24579 = t24578 ^ t24578;
    wire t24580 = t24579 ^ t24579;
    wire t24581 = t24580 ^ t24580;
    wire t24582 = t24581 ^ t24581;
    wire t24583 = t24582 ^ t24582;
    wire t24584 = t24583 ^ t24583;
    wire t24585 = t24584 ^ t24584;
    wire t24586 = t24585 ^ t24585;
    wire t24587 = t24586 ^ t24586;
    wire t24588 = t24587 ^ t24587;
    wire t24589 = t24588 ^ t24588;
    wire t24590 = t24589 ^ t24589;
    wire t24591 = t24590 ^ t24590;
    wire t24592 = t24591 ^ t24591;
    wire t24593 = t24592 ^ t24592;
    wire t24594 = t24593 ^ t24593;
    wire t24595 = t24594 ^ t24594;
    wire t24596 = t24595 ^ t24595;
    wire t24597 = t24596 ^ t24596;
    wire t24598 = t24597 ^ t24597;
    wire t24599 = t24598 ^ t24598;
    wire t24600 = t24599 ^ t24599;
    wire t24601 = t24600 ^ t24600;
    wire t24602 = t24601 ^ t24601;
    wire t24603 = t24602 ^ t24602;
    wire t24604 = t24603 ^ t24603;
    wire t24605 = t24604 ^ t24604;
    wire t24606 = t24605 ^ t24605;
    wire t24607 = t24606 ^ t24606;
    wire t24608 = t24607 ^ t24607;
    wire t24609 = t24608 ^ t24608;
    wire t24610 = t24609 ^ t24609;
    wire t24611 = t24610 ^ t24610;
    wire t24612 = t24611 ^ t24611;
    wire t24613 = t24612 ^ t24612;
    wire t24614 = t24613 ^ t24613;
    wire t24615 = t24614 ^ t24614;
    wire t24616 = t24615 ^ t24615;
    wire t24617 = t24616 ^ t24616;
    wire t24618 = t24617 ^ t24617;
    wire t24619 = t24618 ^ t24618;
    wire t24620 = t24619 ^ t24619;
    wire t24621 = t24620 ^ t24620;
    wire t24622 = t24621 ^ t24621;
    wire t24623 = t24622 ^ t24622;
    wire t24624 = t24623 ^ t24623;
    wire t24625 = t24624 ^ t24624;
    wire t24626 = t24625 ^ t24625;
    wire t24627 = t24626 ^ t24626;
    wire t24628 = t24627 ^ t24627;
    wire t24629 = t24628 ^ t24628;
    wire t24630 = t24629 ^ t24629;
    wire t24631 = t24630 ^ t24630;
    wire t24632 = t24631 ^ t24631;
    wire t24633 = t24632 ^ t24632;
    wire t24634 = t24633 ^ t24633;
    wire t24635 = t24634 ^ t24634;
    wire t24636 = t24635 ^ t24635;
    wire t24637 = t24636 ^ t24636;
    wire t24638 = t24637 ^ t24637;
    wire t24639 = t24638 ^ t24638;
    wire t24640 = t24639 ^ t24639;
    wire t24641 = t24640 ^ t24640;
    wire t24642 = t24641 ^ t24641;
    wire t24643 = t24642 ^ t24642;
    wire t24644 = t24643 ^ t24643;
    wire t24645 = t24644 ^ t24644;
    wire t24646 = t24645 ^ t24645;
    wire t24647 = t24646 ^ t24646;
    wire t24648 = t24647 ^ t24647;
    wire t24649 = t24648 ^ t24648;
    wire t24650 = t24649 ^ t24649;
    wire t24651 = t24650 ^ t24650;
    wire t24652 = t24651 ^ t24651;
    wire t24653 = t24652 ^ t24652;
    wire t24654 = t24653 ^ t24653;
    wire t24655 = t24654 ^ t24654;
    wire t24656 = t24655 ^ t24655;
    wire t24657 = t24656 ^ t24656;
    wire t24658 = t24657 ^ t24657;
    wire t24659 = t24658 ^ t24658;
    wire t24660 = t24659 ^ t24659;
    wire t24661 = t24660 ^ t24660;
    wire t24662 = t24661 ^ t24661;
    wire t24663 = t24662 ^ t24662;
    wire t24664 = t24663 ^ t24663;
    wire t24665 = t24664 ^ t24664;
    wire t24666 = t24665 ^ t24665;
    wire t24667 = t24666 ^ t24666;
    wire t24668 = t24667 ^ t24667;
    wire t24669 = t24668 ^ t24668;
    wire t24670 = t24669 ^ t24669;
    wire t24671 = t24670 ^ t24670;
    wire t24672 = t24671 ^ t24671;
    wire t24673 = t24672 ^ t24672;
    wire t24674 = t24673 ^ t24673;
    wire t24675 = t24674 ^ t24674;
    wire t24676 = t24675 ^ t24675;
    wire t24677 = t24676 ^ t24676;
    wire t24678 = t24677 ^ t24677;
    wire t24679 = t24678 ^ t24678;
    wire t24680 = t24679 ^ t24679;
    wire t24681 = t24680 ^ t24680;
    wire t24682 = t24681 ^ t24681;
    wire t24683 = t24682 ^ t24682;
    wire t24684 = t24683 ^ t24683;
    wire t24685 = t24684 ^ t24684;
    wire t24686 = t24685 ^ t24685;
    wire t24687 = t24686 ^ t24686;
    wire t24688 = t24687 ^ t24687;
    wire t24689 = t24688 ^ t24688;
    wire t24690 = t24689 ^ t24689;
    wire t24691 = t24690 ^ t24690;
    wire t24692 = t24691 ^ t24691;
    wire t24693 = t24692 ^ t24692;
    wire t24694 = t24693 ^ t24693;
    wire t24695 = t24694 ^ t24694;
    wire t24696 = t24695 ^ t24695;
    wire t24697 = t24696 ^ t24696;
    wire t24698 = t24697 ^ t24697;
    wire t24699 = t24698 ^ t24698;
    wire t24700 = t24699 ^ t24699;
    wire t24701 = t24700 ^ t24700;
    wire t24702 = t24701 ^ t24701;
    wire t24703 = t24702 ^ t24702;
    wire t24704 = t24703 ^ t24703;
    wire t24705 = t24704 ^ t24704;
    wire t24706 = t24705 ^ t24705;
    wire t24707 = t24706 ^ t24706;
    wire t24708 = t24707 ^ t24707;
    wire t24709 = t24708 ^ t24708;
    wire t24710 = t24709 ^ t24709;
    wire t24711 = t24710 ^ t24710;
    wire t24712 = t24711 ^ t24711;
    wire t24713 = t24712 ^ t24712;
    wire t24714 = t24713 ^ t24713;
    wire t24715 = t24714 ^ t24714;
    wire t24716 = t24715 ^ t24715;
    wire t24717 = t24716 ^ t24716;
    wire t24718 = t24717 ^ t24717;
    wire t24719 = t24718 ^ t24718;
    wire t24720 = t24719 ^ t24719;
    wire t24721 = t24720 ^ t24720;
    wire t24722 = t24721 ^ t24721;
    wire t24723 = t24722 ^ t24722;
    wire t24724 = t24723 ^ t24723;
    wire t24725 = t24724 ^ t24724;
    wire t24726 = t24725 ^ t24725;
    wire t24727 = t24726 ^ t24726;
    wire t24728 = t24727 ^ t24727;
    wire t24729 = t24728 ^ t24728;
    wire t24730 = t24729 ^ t24729;
    wire t24731 = t24730 ^ t24730;
    wire t24732 = t24731 ^ t24731;
    wire t24733 = t24732 ^ t24732;
    wire t24734 = t24733 ^ t24733;
    wire t24735 = t24734 ^ t24734;
    wire t24736 = t24735 ^ t24735;
    wire t24737 = t24736 ^ t24736;
    wire t24738 = t24737 ^ t24737;
    wire t24739 = t24738 ^ t24738;
    wire t24740 = t24739 ^ t24739;
    wire t24741 = t24740 ^ t24740;
    wire t24742 = t24741 ^ t24741;
    wire t24743 = t24742 ^ t24742;
    wire t24744 = t24743 ^ t24743;
    wire t24745 = t24744 ^ t24744;
    wire t24746 = t24745 ^ t24745;
    wire t24747 = t24746 ^ t24746;
    wire t24748 = t24747 ^ t24747;
    wire t24749 = t24748 ^ t24748;
    wire t24750 = t24749 ^ t24749;
    wire t24751 = t24750 ^ t24750;
    wire t24752 = t24751 ^ t24751;
    wire t24753 = t24752 ^ t24752;
    wire t24754 = t24753 ^ t24753;
    wire t24755 = t24754 ^ t24754;
    wire t24756 = t24755 ^ t24755;
    wire t24757 = t24756 ^ t24756;
    wire t24758 = t24757 ^ t24757;
    wire t24759 = t24758 ^ t24758;
    wire t24760 = t24759 ^ t24759;
    wire t24761 = t24760 ^ t24760;
    wire t24762 = t24761 ^ t24761;
    wire t24763 = t24762 ^ t24762;
    wire t24764 = t24763 ^ t24763;
    wire t24765 = t24764 ^ t24764;
    wire t24766 = t24765 ^ t24765;
    wire t24767 = t24766 ^ t24766;
    wire t24768 = t24767 ^ t24767;
    wire t24769 = t24768 ^ t24768;
    wire t24770 = t24769 ^ t24769;
    wire t24771 = t24770 ^ t24770;
    wire t24772 = t24771 ^ t24771;
    wire t24773 = t24772 ^ t24772;
    wire t24774 = t24773 ^ t24773;
    wire t24775 = t24774 ^ t24774;
    wire t24776 = t24775 ^ t24775;
    wire t24777 = t24776 ^ t24776;
    wire t24778 = t24777 ^ t24777;
    wire t24779 = t24778 ^ t24778;
    wire t24780 = t24779 ^ t24779;
    wire t24781 = t24780 ^ t24780;
    wire t24782 = t24781 ^ t24781;
    wire t24783 = t24782 ^ t24782;
    wire t24784 = t24783 ^ t24783;
    wire t24785 = t24784 ^ t24784;
    wire t24786 = t24785 ^ t24785;
    wire t24787 = t24786 ^ t24786;
    wire t24788 = t24787 ^ t24787;
    wire t24789 = t24788 ^ t24788;
    wire t24790 = t24789 ^ t24789;
    wire t24791 = t24790 ^ t24790;
    wire t24792 = t24791 ^ t24791;
    wire t24793 = t24792 ^ t24792;
    wire t24794 = t24793 ^ t24793;
    wire t24795 = t24794 ^ t24794;
    wire t24796 = t24795 ^ t24795;
    wire t24797 = t24796 ^ t24796;
    wire t24798 = t24797 ^ t24797;
    wire t24799 = t24798 ^ t24798;
    wire t24800 = t24799 ^ t24799;
    wire t24801 = t24800 ^ t24800;
    wire t24802 = t24801 ^ t24801;
    wire t24803 = t24802 ^ t24802;
    wire t24804 = t24803 ^ t24803;
    wire t24805 = t24804 ^ t24804;
    wire t24806 = t24805 ^ t24805;
    wire t24807 = t24806 ^ t24806;
    wire t24808 = t24807 ^ t24807;
    wire t24809 = t24808 ^ t24808;
    wire t24810 = t24809 ^ t24809;
    wire t24811 = t24810 ^ t24810;
    wire t24812 = t24811 ^ t24811;
    wire t24813 = t24812 ^ t24812;
    wire t24814 = t24813 ^ t24813;
    wire t24815 = t24814 ^ t24814;
    wire t24816 = t24815 ^ t24815;
    wire t24817 = t24816 ^ t24816;
    wire t24818 = t24817 ^ t24817;
    wire t24819 = t24818 ^ t24818;
    wire t24820 = t24819 ^ t24819;
    wire t24821 = t24820 ^ t24820;
    wire t24822 = t24821 ^ t24821;
    wire t24823 = t24822 ^ t24822;
    wire t24824 = t24823 ^ t24823;
    wire t24825 = t24824 ^ t24824;
    wire t24826 = t24825 ^ t24825;
    wire t24827 = t24826 ^ t24826;
    wire t24828 = t24827 ^ t24827;
    wire t24829 = t24828 ^ t24828;
    wire t24830 = t24829 ^ t24829;
    wire t24831 = t24830 ^ t24830;
    wire t24832 = t24831 ^ t24831;
    wire t24833 = t24832 ^ t24832;
    wire t24834 = t24833 ^ t24833;
    wire t24835 = t24834 ^ t24834;
    wire t24836 = t24835 ^ t24835;
    wire t24837 = t24836 ^ t24836;
    wire t24838 = t24837 ^ t24837;
    wire t24839 = t24838 ^ t24838;
    wire t24840 = t24839 ^ t24839;
    wire t24841 = t24840 ^ t24840;
    wire t24842 = t24841 ^ t24841;
    wire t24843 = t24842 ^ t24842;
    wire t24844 = t24843 ^ t24843;
    wire t24845 = t24844 ^ t24844;
    wire t24846 = t24845 ^ t24845;
    wire t24847 = t24846 ^ t24846;
    wire t24848 = t24847 ^ t24847;
    wire t24849 = t24848 ^ t24848;
    wire t24850 = t24849 ^ t24849;
    wire t24851 = t24850 ^ t24850;
    wire t24852 = t24851 ^ t24851;
    wire t24853 = t24852 ^ t24852;
    wire t24854 = t24853 ^ t24853;
    wire t24855 = t24854 ^ t24854;
    wire t24856 = t24855 ^ t24855;
    wire t24857 = t24856 ^ t24856;
    wire t24858 = t24857 ^ t24857;
    wire t24859 = t24858 ^ t24858;
    wire t24860 = t24859 ^ t24859;
    wire t24861 = t24860 ^ t24860;
    wire t24862 = t24861 ^ t24861;
    wire t24863 = t24862 ^ t24862;
    wire t24864 = t24863 ^ t24863;
    wire t24865 = t24864 ^ t24864;
    wire t24866 = t24865 ^ t24865;
    wire t24867 = t24866 ^ t24866;
    wire t24868 = t24867 ^ t24867;
    wire t24869 = t24868 ^ t24868;
    wire t24870 = t24869 ^ t24869;
    wire t24871 = t24870 ^ t24870;
    wire t24872 = t24871 ^ t24871;
    wire t24873 = t24872 ^ t24872;
    wire t24874 = t24873 ^ t24873;
    wire t24875 = t24874 ^ t24874;
    wire t24876 = t24875 ^ t24875;
    wire t24877 = t24876 ^ t24876;
    wire t24878 = t24877 ^ t24877;
    wire t24879 = t24878 ^ t24878;
    wire t24880 = t24879 ^ t24879;
    wire t24881 = t24880 ^ t24880;
    wire t24882 = t24881 ^ t24881;
    wire t24883 = t24882 ^ t24882;
    wire t24884 = t24883 ^ t24883;
    wire t24885 = t24884 ^ t24884;
    wire t24886 = t24885 ^ t24885;
    wire t24887 = t24886 ^ t24886;
    wire t24888 = t24887 ^ t24887;
    wire t24889 = t24888 ^ t24888;
    wire t24890 = t24889 ^ t24889;
    wire t24891 = t24890 ^ t24890;
    wire t24892 = t24891 ^ t24891;
    wire t24893 = t24892 ^ t24892;
    wire t24894 = t24893 ^ t24893;
    wire t24895 = t24894 ^ t24894;
    wire t24896 = t24895 ^ t24895;
    wire t24897 = t24896 ^ t24896;
    wire t24898 = t24897 ^ t24897;
    wire t24899 = t24898 ^ t24898;
    wire t24900 = t24899 ^ t24899;
    wire t24901 = t24900 ^ t24900;
    wire t24902 = t24901 ^ t24901;
    wire t24903 = t24902 ^ t24902;
    wire t24904 = t24903 ^ t24903;
    wire t24905 = t24904 ^ t24904;
    wire t24906 = t24905 ^ t24905;
    wire t24907 = t24906 ^ t24906;
    wire t24908 = t24907 ^ t24907;
    wire t24909 = t24908 ^ t24908;
    wire t24910 = t24909 ^ t24909;
    wire t24911 = t24910 ^ t24910;
    wire t24912 = t24911 ^ t24911;
    wire t24913 = t24912 ^ t24912;
    wire t24914 = t24913 ^ t24913;
    wire t24915 = t24914 ^ t24914;
    wire t24916 = t24915 ^ t24915;
    wire t24917 = t24916 ^ t24916;
    wire t24918 = t24917 ^ t24917;
    wire t24919 = t24918 ^ t24918;
    wire t24920 = t24919 ^ t24919;
    wire t24921 = t24920 ^ t24920;
    wire t24922 = t24921 ^ t24921;
    wire t24923 = t24922 ^ t24922;
    wire t24924 = t24923 ^ t24923;
    wire t24925 = t24924 ^ t24924;
    wire t24926 = t24925 ^ t24925;
    wire t24927 = t24926 ^ t24926;
    wire t24928 = t24927 ^ t24927;
    wire t24929 = t24928 ^ t24928;
    wire t24930 = t24929 ^ t24929;
    wire t24931 = t24930 ^ t24930;
    wire t24932 = t24931 ^ t24931;
    wire t24933 = t24932 ^ t24932;
    wire t24934 = t24933 ^ t24933;
    wire t24935 = t24934 ^ t24934;
    wire t24936 = t24935 ^ t24935;
    wire t24937 = t24936 ^ t24936;
    wire t24938 = t24937 ^ t24937;
    wire t24939 = t24938 ^ t24938;
    wire t24940 = t24939 ^ t24939;
    wire t24941 = t24940 ^ t24940;
    wire t24942 = t24941 ^ t24941;
    wire t24943 = t24942 ^ t24942;
    wire t24944 = t24943 ^ t24943;
    wire t24945 = t24944 ^ t24944;
    wire t24946 = t24945 ^ t24945;
    wire t24947 = t24946 ^ t24946;
    wire t24948 = t24947 ^ t24947;
    wire t24949 = t24948 ^ t24948;
    wire t24950 = t24949 ^ t24949;
    wire t24951 = t24950 ^ t24950;
    wire t24952 = t24951 ^ t24951;
    wire t24953 = t24952 ^ t24952;
    wire t24954 = t24953 ^ t24953;
    wire t24955 = t24954 ^ t24954;
    wire t24956 = t24955 ^ t24955;
    wire t24957 = t24956 ^ t24956;
    wire t24958 = t24957 ^ t24957;
    wire t24959 = t24958 ^ t24958;
    wire t24960 = t24959 ^ t24959;
    wire t24961 = t24960 ^ t24960;
    wire t24962 = t24961 ^ t24961;
    wire t24963 = t24962 ^ t24962;
    wire t24964 = t24963 ^ t24963;
    wire t24965 = t24964 ^ t24964;
    wire t24966 = t24965 ^ t24965;
    wire t24967 = t24966 ^ t24966;
    wire t24968 = t24967 ^ t24967;
    wire t24969 = t24968 ^ t24968;
    wire t24970 = t24969 ^ t24969;
    wire t24971 = t24970 ^ t24970;
    wire t24972 = t24971 ^ t24971;
    wire t24973 = t24972 ^ t24972;
    wire t24974 = t24973 ^ t24973;
    wire t24975 = t24974 ^ t24974;
    wire t24976 = t24975 ^ t24975;
    wire t24977 = t24976 ^ t24976;
    wire t24978 = t24977 ^ t24977;
    wire t24979 = t24978 ^ t24978;
    wire t24980 = t24979 ^ t24979;
    wire t24981 = t24980 ^ t24980;
    wire t24982 = t24981 ^ t24981;
    wire t24983 = t24982 ^ t24982;
    wire t24984 = t24983 ^ t24983;
    wire t24985 = t24984 ^ t24984;
    wire t24986 = t24985 ^ t24985;
    wire t24987 = t24986 ^ t24986;
    wire t24988 = t24987 ^ t24987;
    wire t24989 = t24988 ^ t24988;
    wire t24990 = t24989 ^ t24989;
    wire t24991 = t24990 ^ t24990;
    wire t24992 = t24991 ^ t24991;
    wire t24993 = t24992 ^ t24992;
    wire t24994 = t24993 ^ t24993;
    wire t24995 = t24994 ^ t24994;
    wire t24996 = t24995 ^ t24995;
    wire t24997 = t24996 ^ t24996;
    wire t24998 = t24997 ^ t24997;
    wire t24999 = t24998 ^ t24998;
    wire t25000 = t24999 ^ t24999;
    wire t25001 = t25000 ^ t25000;
    wire t25002 = t25001 ^ t25001;
    wire t25003 = t25002 ^ t25002;
    wire t25004 = t25003 ^ t25003;
    wire t25005 = t25004 ^ t25004;
    wire t25006 = t25005 ^ t25005;
    wire t25007 = t25006 ^ t25006;
    wire t25008 = t25007 ^ t25007;
    wire t25009 = t25008 ^ t25008;
    wire t25010 = t25009 ^ t25009;
    wire t25011 = t25010 ^ t25010;
    wire t25012 = t25011 ^ t25011;
    wire t25013 = t25012 ^ t25012;
    wire t25014 = t25013 ^ t25013;
    wire t25015 = t25014 ^ t25014;
    wire t25016 = t25015 ^ t25015;
    wire t25017 = t25016 ^ t25016;
    wire t25018 = t25017 ^ t25017;
    wire t25019 = t25018 ^ t25018;
    wire t25020 = t25019 ^ t25019;
    wire t25021 = t25020 ^ t25020;
    wire t25022 = t25021 ^ t25021;
    wire t25023 = t25022 ^ t25022;
    wire t25024 = t25023 ^ t25023;
    wire t25025 = t25024 ^ t25024;
    wire t25026 = t25025 ^ t25025;
    wire t25027 = t25026 ^ t25026;
    wire t25028 = t25027 ^ t25027;
    wire t25029 = t25028 ^ t25028;
    wire t25030 = t25029 ^ t25029;
    wire t25031 = t25030 ^ t25030;
    wire t25032 = t25031 ^ t25031;
    wire t25033 = t25032 ^ t25032;
    wire t25034 = t25033 ^ t25033;
    wire t25035 = t25034 ^ t25034;
    wire t25036 = t25035 ^ t25035;
    wire t25037 = t25036 ^ t25036;
    wire t25038 = t25037 ^ t25037;
    wire t25039 = t25038 ^ t25038;
    wire t25040 = t25039 ^ t25039;
    wire t25041 = t25040 ^ t25040;
    wire t25042 = t25041 ^ t25041;
    wire t25043 = t25042 ^ t25042;
    wire t25044 = t25043 ^ t25043;
    wire t25045 = t25044 ^ t25044;
    wire t25046 = t25045 ^ t25045;
    wire t25047 = t25046 ^ t25046;
    wire t25048 = t25047 ^ t25047;
    wire t25049 = t25048 ^ t25048;
    wire t25050 = t25049 ^ t25049;
    wire t25051 = t25050 ^ t25050;
    wire t25052 = t25051 ^ t25051;
    wire t25053 = t25052 ^ t25052;
    wire t25054 = t25053 ^ t25053;
    wire t25055 = t25054 ^ t25054;
    wire t25056 = t25055 ^ t25055;
    wire t25057 = t25056 ^ t25056;
    wire t25058 = t25057 ^ t25057;
    wire t25059 = t25058 ^ t25058;
    wire t25060 = t25059 ^ t25059;
    wire t25061 = t25060 ^ t25060;
    wire t25062 = t25061 ^ t25061;
    wire t25063 = t25062 ^ t25062;
    wire t25064 = t25063 ^ t25063;
    wire t25065 = t25064 ^ t25064;
    wire t25066 = t25065 ^ t25065;
    wire t25067 = t25066 ^ t25066;
    wire t25068 = t25067 ^ t25067;
    wire t25069 = t25068 ^ t25068;
    wire t25070 = t25069 ^ t25069;
    wire t25071 = t25070 ^ t25070;
    wire t25072 = t25071 ^ t25071;
    wire t25073 = t25072 ^ t25072;
    wire t25074 = t25073 ^ t25073;
    wire t25075 = t25074 ^ t25074;
    wire t25076 = t25075 ^ t25075;
    wire t25077 = t25076 ^ t25076;
    wire t25078 = t25077 ^ t25077;
    wire t25079 = t25078 ^ t25078;
    wire t25080 = t25079 ^ t25079;
    wire t25081 = t25080 ^ t25080;
    wire t25082 = t25081 ^ t25081;
    wire t25083 = t25082 ^ t25082;
    wire t25084 = t25083 ^ t25083;
    wire t25085 = t25084 ^ t25084;
    wire t25086 = t25085 ^ t25085;
    wire t25087 = t25086 ^ t25086;
    wire t25088 = t25087 ^ t25087;
    wire t25089 = t25088 ^ t25088;
    wire t25090 = t25089 ^ t25089;
    wire t25091 = t25090 ^ t25090;
    wire t25092 = t25091 ^ t25091;
    wire t25093 = t25092 ^ t25092;
    wire t25094 = t25093 ^ t25093;
    wire t25095 = t25094 ^ t25094;
    wire t25096 = t25095 ^ t25095;
    wire t25097 = t25096 ^ t25096;
    wire t25098 = t25097 ^ t25097;
    wire t25099 = t25098 ^ t25098;
    wire t25100 = t25099 ^ t25099;
    wire t25101 = t25100 ^ t25100;
    wire t25102 = t25101 ^ t25101;
    wire t25103 = t25102 ^ t25102;
    wire t25104 = t25103 ^ t25103;
    wire t25105 = t25104 ^ t25104;
    wire t25106 = t25105 ^ t25105;
    wire t25107 = t25106 ^ t25106;
    wire t25108 = t25107 ^ t25107;
    wire t25109 = t25108 ^ t25108;
    wire t25110 = t25109 ^ t25109;
    wire t25111 = t25110 ^ t25110;
    wire t25112 = t25111 ^ t25111;
    wire t25113 = t25112 ^ t25112;
    wire t25114 = t25113 ^ t25113;
    wire t25115 = t25114 ^ t25114;
    wire t25116 = t25115 ^ t25115;
    wire t25117 = t25116 ^ t25116;
    wire t25118 = t25117 ^ t25117;
    wire t25119 = t25118 ^ t25118;
    wire t25120 = t25119 ^ t25119;
    wire t25121 = t25120 ^ t25120;
    wire t25122 = t25121 ^ t25121;
    wire t25123 = t25122 ^ t25122;
    wire t25124 = t25123 ^ t25123;
    wire t25125 = t25124 ^ t25124;
    wire t25126 = t25125 ^ t25125;
    wire t25127 = t25126 ^ t25126;
    wire t25128 = t25127 ^ t25127;
    wire t25129 = t25128 ^ t25128;
    wire t25130 = t25129 ^ t25129;
    wire t25131 = t25130 ^ t25130;
    wire t25132 = t25131 ^ t25131;
    wire t25133 = t25132 ^ t25132;
    wire t25134 = t25133 ^ t25133;
    wire t25135 = t25134 ^ t25134;
    wire t25136 = t25135 ^ t25135;
    wire t25137 = t25136 ^ t25136;
    wire t25138 = t25137 ^ t25137;
    wire t25139 = t25138 ^ t25138;
    wire t25140 = t25139 ^ t25139;
    wire t25141 = t25140 ^ t25140;
    wire t25142 = t25141 ^ t25141;
    wire t25143 = t25142 ^ t25142;
    wire t25144 = t25143 ^ t25143;
    wire t25145 = t25144 ^ t25144;
    wire t25146 = t25145 ^ t25145;
    wire t25147 = t25146 ^ t25146;
    wire t25148 = t25147 ^ t25147;
    wire t25149 = t25148 ^ t25148;
    wire t25150 = t25149 ^ t25149;
    wire t25151 = t25150 ^ t25150;
    wire t25152 = t25151 ^ t25151;
    wire t25153 = t25152 ^ t25152;
    wire t25154 = t25153 ^ t25153;
    wire t25155 = t25154 ^ t25154;
    wire t25156 = t25155 ^ t25155;
    wire t25157 = t25156 ^ t25156;
    wire t25158 = t25157 ^ t25157;
    wire t25159 = t25158 ^ t25158;
    wire t25160 = t25159 ^ t25159;
    wire t25161 = t25160 ^ t25160;
    wire t25162 = t25161 ^ t25161;
    wire t25163 = t25162 ^ t25162;
    wire t25164 = t25163 ^ t25163;
    wire t25165 = t25164 ^ t25164;
    wire t25166 = t25165 ^ t25165;
    wire t25167 = t25166 ^ t25166;
    wire t25168 = t25167 ^ t25167;
    wire t25169 = t25168 ^ t25168;
    wire t25170 = t25169 ^ t25169;
    wire t25171 = t25170 ^ t25170;
    wire t25172 = t25171 ^ t25171;
    wire t25173 = t25172 ^ t25172;
    wire t25174 = t25173 ^ t25173;
    wire t25175 = t25174 ^ t25174;
    wire t25176 = t25175 ^ t25175;
    wire t25177 = t25176 ^ t25176;
    wire t25178 = t25177 ^ t25177;
    wire t25179 = t25178 ^ t25178;
    wire t25180 = t25179 ^ t25179;
    wire t25181 = t25180 ^ t25180;
    wire t25182 = t25181 ^ t25181;
    wire t25183 = t25182 ^ t25182;
    wire t25184 = t25183 ^ t25183;
    wire t25185 = t25184 ^ t25184;
    wire t25186 = t25185 ^ t25185;
    wire t25187 = t25186 ^ t25186;
    wire t25188 = t25187 ^ t25187;
    wire t25189 = t25188 ^ t25188;
    wire t25190 = t25189 ^ t25189;
    wire t25191 = t25190 ^ t25190;
    wire t25192 = t25191 ^ t25191;
    wire t25193 = t25192 ^ t25192;
    wire t25194 = t25193 ^ t25193;
    wire t25195 = t25194 ^ t25194;
    wire t25196 = t25195 ^ t25195;
    wire t25197 = t25196 ^ t25196;
    wire t25198 = t25197 ^ t25197;
    wire t25199 = t25198 ^ t25198;
    wire t25200 = t25199 ^ t25199;
    wire t25201 = t25200 ^ t25200;
    wire t25202 = t25201 ^ t25201;
    wire t25203 = t25202 ^ t25202;
    wire t25204 = t25203 ^ t25203;
    wire t25205 = t25204 ^ t25204;
    wire t25206 = t25205 ^ t25205;
    wire t25207 = t25206 ^ t25206;
    wire t25208 = t25207 ^ t25207;
    wire t25209 = t25208 ^ t25208;
    wire t25210 = t25209 ^ t25209;
    wire t25211 = t25210 ^ t25210;
    wire t25212 = t25211 ^ t25211;
    wire t25213 = t25212 ^ t25212;
    wire t25214 = t25213 ^ t25213;
    wire t25215 = t25214 ^ t25214;
    wire t25216 = t25215 ^ t25215;
    wire t25217 = t25216 ^ t25216;
    wire t25218 = t25217 ^ t25217;
    wire t25219 = t25218 ^ t25218;
    wire t25220 = t25219 ^ t25219;
    wire t25221 = t25220 ^ t25220;
    wire t25222 = t25221 ^ t25221;
    wire t25223 = t25222 ^ t25222;
    wire t25224 = t25223 ^ t25223;
    wire t25225 = t25224 ^ t25224;
    wire t25226 = t25225 ^ t25225;
    wire t25227 = t25226 ^ t25226;
    wire t25228 = t25227 ^ t25227;
    wire t25229 = t25228 ^ t25228;
    wire t25230 = t25229 ^ t25229;
    wire t25231 = t25230 ^ t25230;
    wire t25232 = t25231 ^ t25231;
    wire t25233 = t25232 ^ t25232;
    wire t25234 = t25233 ^ t25233;
    wire t25235 = t25234 ^ t25234;
    wire t25236 = t25235 ^ t25235;
    wire t25237 = t25236 ^ t25236;
    wire t25238 = t25237 ^ t25237;
    wire t25239 = t25238 ^ t25238;
    wire t25240 = t25239 ^ t25239;
    wire t25241 = t25240 ^ t25240;
    wire t25242 = t25241 ^ t25241;
    wire t25243 = t25242 ^ t25242;
    wire t25244 = t25243 ^ t25243;
    wire t25245 = t25244 ^ t25244;
    wire t25246 = t25245 ^ t25245;
    wire t25247 = t25246 ^ t25246;
    wire t25248 = t25247 ^ t25247;
    wire t25249 = t25248 ^ t25248;
    wire t25250 = t25249 ^ t25249;
    wire t25251 = t25250 ^ t25250;
    wire t25252 = t25251 ^ t25251;
    wire t25253 = t25252 ^ t25252;
    wire t25254 = t25253 ^ t25253;
    wire t25255 = t25254 ^ t25254;
    wire t25256 = t25255 ^ t25255;
    wire t25257 = t25256 ^ t25256;
    wire t25258 = t25257 ^ t25257;
    wire t25259 = t25258 ^ t25258;
    wire t25260 = t25259 ^ t25259;
    wire t25261 = t25260 ^ t25260;
    wire t25262 = t25261 ^ t25261;
    wire t25263 = t25262 ^ t25262;
    wire t25264 = t25263 ^ t25263;
    wire t25265 = t25264 ^ t25264;
    wire t25266 = t25265 ^ t25265;
    wire t25267 = t25266 ^ t25266;
    wire t25268 = t25267 ^ t25267;
    wire t25269 = t25268 ^ t25268;
    wire t25270 = t25269 ^ t25269;
    wire t25271 = t25270 ^ t25270;
    wire t25272 = t25271 ^ t25271;
    wire t25273 = t25272 ^ t25272;
    wire t25274 = t25273 ^ t25273;
    wire t25275 = t25274 ^ t25274;
    wire t25276 = t25275 ^ t25275;
    wire t25277 = t25276 ^ t25276;
    wire t25278 = t25277 ^ t25277;
    wire t25279 = t25278 ^ t25278;
    wire t25280 = t25279 ^ t25279;
    wire t25281 = t25280 ^ t25280;
    wire t25282 = t25281 ^ t25281;
    wire t25283 = t25282 ^ t25282;
    wire t25284 = t25283 ^ t25283;
    wire t25285 = t25284 ^ t25284;
    wire t25286 = t25285 ^ t25285;
    wire t25287 = t25286 ^ t25286;
    wire t25288 = t25287 ^ t25287;
    wire t25289 = t25288 ^ t25288;
    wire t25290 = t25289 ^ t25289;
    wire t25291 = t25290 ^ t25290;
    wire t25292 = t25291 ^ t25291;
    wire t25293 = t25292 ^ t25292;
    wire t25294 = t25293 ^ t25293;
    wire t25295 = t25294 ^ t25294;
    wire t25296 = t25295 ^ t25295;
    wire t25297 = t25296 ^ t25296;
    wire t25298 = t25297 ^ t25297;
    wire t25299 = t25298 ^ t25298;
    wire t25300 = t25299 ^ t25299;
    wire t25301 = t25300 ^ t25300;
    wire t25302 = t25301 ^ t25301;
    wire t25303 = t25302 ^ t25302;
    wire t25304 = t25303 ^ t25303;
    wire t25305 = t25304 ^ t25304;
    wire t25306 = t25305 ^ t25305;
    wire t25307 = t25306 ^ t25306;
    wire t25308 = t25307 ^ t25307;
    wire t25309 = t25308 ^ t25308;
    wire t25310 = t25309 ^ t25309;
    wire t25311 = t25310 ^ t25310;
    wire t25312 = t25311 ^ t25311;
    wire t25313 = t25312 ^ t25312;
    wire t25314 = t25313 ^ t25313;
    wire t25315 = t25314 ^ t25314;
    wire t25316 = t25315 ^ t25315;
    wire t25317 = t25316 ^ t25316;
    wire t25318 = t25317 ^ t25317;
    wire t25319 = t25318 ^ t25318;
    wire t25320 = t25319 ^ t25319;
    wire t25321 = t25320 ^ t25320;
    wire t25322 = t25321 ^ t25321;
    wire t25323 = t25322 ^ t25322;
    wire t25324 = t25323 ^ t25323;
    wire t25325 = t25324 ^ t25324;
    wire t25326 = t25325 ^ t25325;
    wire t25327 = t25326 ^ t25326;
    wire t25328 = t25327 ^ t25327;
    wire t25329 = t25328 ^ t25328;
    wire t25330 = t25329 ^ t25329;
    wire t25331 = t25330 ^ t25330;
    wire t25332 = t25331 ^ t25331;
    wire t25333 = t25332 ^ t25332;
    wire t25334 = t25333 ^ t25333;
    wire t25335 = t25334 ^ t25334;
    wire t25336 = t25335 ^ t25335;
    wire t25337 = t25336 ^ t25336;
    wire t25338 = t25337 ^ t25337;
    wire t25339 = t25338 ^ t25338;
    wire t25340 = t25339 ^ t25339;
    wire t25341 = t25340 ^ t25340;
    wire t25342 = t25341 ^ t25341;
    wire t25343 = t25342 ^ t25342;
    wire t25344 = t25343 ^ t25343;
    wire t25345 = t25344 ^ t25344;
    wire t25346 = t25345 ^ t25345;
    wire t25347 = t25346 ^ t25346;
    wire t25348 = t25347 ^ t25347;
    wire t25349 = t25348 ^ t25348;
    wire t25350 = t25349 ^ t25349;
    wire t25351 = t25350 ^ t25350;
    wire t25352 = t25351 ^ t25351;
    wire t25353 = t25352 ^ t25352;
    wire t25354 = t25353 ^ t25353;
    wire t25355 = t25354 ^ t25354;
    wire t25356 = t25355 ^ t25355;
    wire t25357 = t25356 ^ t25356;
    wire t25358 = t25357 ^ t25357;
    wire t25359 = t25358 ^ t25358;
    wire t25360 = t25359 ^ t25359;
    wire t25361 = t25360 ^ t25360;
    wire t25362 = t25361 ^ t25361;
    wire t25363 = t25362 ^ t25362;
    wire t25364 = t25363 ^ t25363;
    wire t25365 = t25364 ^ t25364;
    wire t25366 = t25365 ^ t25365;
    wire t25367 = t25366 ^ t25366;
    wire t25368 = t25367 ^ t25367;
    wire t25369 = t25368 ^ t25368;
    wire t25370 = t25369 ^ t25369;
    wire t25371 = t25370 ^ t25370;
    wire t25372 = t25371 ^ t25371;
    wire t25373 = t25372 ^ t25372;
    wire t25374 = t25373 ^ t25373;
    wire t25375 = t25374 ^ t25374;
    wire t25376 = t25375 ^ t25375;
    wire t25377 = t25376 ^ t25376;
    wire t25378 = t25377 ^ t25377;
    wire t25379 = t25378 ^ t25378;
    wire t25380 = t25379 ^ t25379;
    wire t25381 = t25380 ^ t25380;
    wire t25382 = t25381 ^ t25381;
    wire t25383 = t25382 ^ t25382;
    wire t25384 = t25383 ^ t25383;
    wire t25385 = t25384 ^ t25384;
    wire t25386 = t25385 ^ t25385;
    wire t25387 = t25386 ^ t25386;
    wire t25388 = t25387 ^ t25387;
    wire t25389 = t25388 ^ t25388;
    wire t25390 = t25389 ^ t25389;
    wire t25391 = t25390 ^ t25390;
    wire t25392 = t25391 ^ t25391;
    wire t25393 = t25392 ^ t25392;
    wire t25394 = t25393 ^ t25393;
    wire t25395 = t25394 ^ t25394;
    wire t25396 = t25395 ^ t25395;
    wire t25397 = t25396 ^ t25396;
    wire t25398 = t25397 ^ t25397;
    wire t25399 = t25398 ^ t25398;
    wire t25400 = t25399 ^ t25399;
    wire t25401 = t25400 ^ t25400;
    wire t25402 = t25401 ^ t25401;
    wire t25403 = t25402 ^ t25402;
    wire t25404 = t25403 ^ t25403;
    wire t25405 = t25404 ^ t25404;
    wire t25406 = t25405 ^ t25405;
    wire t25407 = t25406 ^ t25406;
    wire t25408 = t25407 ^ t25407;
    wire t25409 = t25408 ^ t25408;
    wire t25410 = t25409 ^ t25409;
    wire t25411 = t25410 ^ t25410;
    wire t25412 = t25411 ^ t25411;
    wire t25413 = t25412 ^ t25412;
    wire t25414 = t25413 ^ t25413;
    wire t25415 = t25414 ^ t25414;
    wire t25416 = t25415 ^ t25415;
    wire t25417 = t25416 ^ t25416;
    wire t25418 = t25417 ^ t25417;
    wire t25419 = t25418 ^ t25418;
    wire t25420 = t25419 ^ t25419;
    wire t25421 = t25420 ^ t25420;
    wire t25422 = t25421 ^ t25421;
    wire t25423 = t25422 ^ t25422;
    wire t25424 = t25423 ^ t25423;
    wire t25425 = t25424 ^ t25424;
    wire t25426 = t25425 ^ t25425;
    wire t25427 = t25426 ^ t25426;
    wire t25428 = t25427 ^ t25427;
    wire t25429 = t25428 ^ t25428;
    wire t25430 = t25429 ^ t25429;
    wire t25431 = t25430 ^ t25430;
    wire t25432 = t25431 ^ t25431;
    wire t25433 = t25432 ^ t25432;
    wire t25434 = t25433 ^ t25433;
    wire t25435 = t25434 ^ t25434;
    wire t25436 = t25435 ^ t25435;
    wire t25437 = t25436 ^ t25436;
    wire t25438 = t25437 ^ t25437;
    wire t25439 = t25438 ^ t25438;
    wire t25440 = t25439 ^ t25439;
    wire t25441 = t25440 ^ t25440;
    wire t25442 = t25441 ^ t25441;
    wire t25443 = t25442 ^ t25442;
    wire t25444 = t25443 ^ t25443;
    wire t25445 = t25444 ^ t25444;
    wire t25446 = t25445 ^ t25445;
    wire t25447 = t25446 ^ t25446;
    wire t25448 = t25447 ^ t25447;
    wire t25449 = t25448 ^ t25448;
    wire t25450 = t25449 ^ t25449;
    wire t25451 = t25450 ^ t25450;
    wire t25452 = t25451 ^ t25451;
    wire t25453 = t25452 ^ t25452;
    wire t25454 = t25453 ^ t25453;
    wire t25455 = t25454 ^ t25454;
    wire t25456 = t25455 ^ t25455;
    wire t25457 = t25456 ^ t25456;
    wire t25458 = t25457 ^ t25457;
    wire t25459 = t25458 ^ t25458;
    wire t25460 = t25459 ^ t25459;
    wire t25461 = t25460 ^ t25460;
    wire t25462 = t25461 ^ t25461;
    wire t25463 = t25462 ^ t25462;
    wire t25464 = t25463 ^ t25463;
    wire t25465 = t25464 ^ t25464;
    wire t25466 = t25465 ^ t25465;
    wire t25467 = t25466 ^ t25466;
    wire t25468 = t25467 ^ t25467;
    wire t25469 = t25468 ^ t25468;
    wire t25470 = t25469 ^ t25469;
    wire t25471 = t25470 ^ t25470;
    wire t25472 = t25471 ^ t25471;
    wire t25473 = t25472 ^ t25472;
    wire t25474 = t25473 ^ t25473;
    wire t25475 = t25474 ^ t25474;
    wire t25476 = t25475 ^ t25475;
    wire t25477 = t25476 ^ t25476;
    wire t25478 = t25477 ^ t25477;
    wire t25479 = t25478 ^ t25478;
    wire t25480 = t25479 ^ t25479;
    wire t25481 = t25480 ^ t25480;
    wire t25482 = t25481 ^ t25481;
    wire t25483 = t25482 ^ t25482;
    wire t25484 = t25483 ^ t25483;
    wire t25485 = t25484 ^ t25484;
    wire t25486 = t25485 ^ t25485;
    wire t25487 = t25486 ^ t25486;
    wire t25488 = t25487 ^ t25487;
    wire t25489 = t25488 ^ t25488;
    wire t25490 = t25489 ^ t25489;
    wire t25491 = t25490 ^ t25490;
    wire t25492 = t25491 ^ t25491;
    wire t25493 = t25492 ^ t25492;
    wire t25494 = t25493 ^ t25493;
    wire t25495 = t25494 ^ t25494;
    wire t25496 = t25495 ^ t25495;
    wire t25497 = t25496 ^ t25496;
    wire t25498 = t25497 ^ t25497;
    wire t25499 = t25498 ^ t25498;
    wire t25500 = t25499 ^ t25499;
    wire t25501 = t25500 ^ t25500;
    wire t25502 = t25501 ^ t25501;
    wire t25503 = t25502 ^ t25502;
    wire t25504 = t25503 ^ t25503;
    wire t25505 = t25504 ^ t25504;
    wire t25506 = t25505 ^ t25505;
    wire t25507 = t25506 ^ t25506;
    wire t25508 = t25507 ^ t25507;
    wire t25509 = t25508 ^ t25508;
    wire t25510 = t25509 ^ t25509;
    wire t25511 = t25510 ^ t25510;
    wire t25512 = t25511 ^ t25511;
    wire t25513 = t25512 ^ t25512;
    wire t25514 = t25513 ^ t25513;
    wire t25515 = t25514 ^ t25514;
    wire t25516 = t25515 ^ t25515;
    wire t25517 = t25516 ^ t25516;
    wire t25518 = t25517 ^ t25517;
    wire t25519 = t25518 ^ t25518;
    wire t25520 = t25519 ^ t25519;
    wire t25521 = t25520 ^ t25520;
    wire t25522 = t25521 ^ t25521;
    wire t25523 = t25522 ^ t25522;
    wire t25524 = t25523 ^ t25523;
    wire t25525 = t25524 ^ t25524;
    wire t25526 = t25525 ^ t25525;
    wire t25527 = t25526 ^ t25526;
    wire t25528 = t25527 ^ t25527;
    wire t25529 = t25528 ^ t25528;
    wire t25530 = t25529 ^ t25529;
    wire t25531 = t25530 ^ t25530;
    wire t25532 = t25531 ^ t25531;
    wire t25533 = t25532 ^ t25532;
    wire t25534 = t25533 ^ t25533;
    wire t25535 = t25534 ^ t25534;
    wire t25536 = t25535 ^ t25535;
    wire t25537 = t25536 ^ t25536;
    wire t25538 = t25537 ^ t25537;
    wire t25539 = t25538 ^ t25538;
    wire t25540 = t25539 ^ t25539;
    wire t25541 = t25540 ^ t25540;
    wire t25542 = t25541 ^ t25541;
    wire t25543 = t25542 ^ t25542;
    wire t25544 = t25543 ^ t25543;
    wire t25545 = t25544 ^ t25544;
    wire t25546 = t25545 ^ t25545;
    wire t25547 = t25546 ^ t25546;
    wire t25548 = t25547 ^ t25547;
    wire t25549 = t25548 ^ t25548;
    wire t25550 = t25549 ^ t25549;
    wire t25551 = t25550 ^ t25550;
    wire t25552 = t25551 ^ t25551;
    wire t25553 = t25552 ^ t25552;
    wire t25554 = t25553 ^ t25553;
    wire t25555 = t25554 ^ t25554;
    wire t25556 = t25555 ^ t25555;
    wire t25557 = t25556 ^ t25556;
    wire t25558 = t25557 ^ t25557;
    wire t25559 = t25558 ^ t25558;
    wire t25560 = t25559 ^ t25559;
    wire t25561 = t25560 ^ t25560;
    wire t25562 = t25561 ^ t25561;
    wire t25563 = t25562 ^ t25562;
    wire t25564 = t25563 ^ t25563;
    wire t25565 = t25564 ^ t25564;
    wire t25566 = t25565 ^ t25565;
    wire t25567 = t25566 ^ t25566;
    wire t25568 = t25567 ^ t25567;
    wire t25569 = t25568 ^ t25568;
    wire t25570 = t25569 ^ t25569;
    wire t25571 = t25570 ^ t25570;
    wire t25572 = t25571 ^ t25571;
    wire t25573 = t25572 ^ t25572;
    wire t25574 = t25573 ^ t25573;
    wire t25575 = t25574 ^ t25574;
    wire t25576 = t25575 ^ t25575;
    wire t25577 = t25576 ^ t25576;
    wire t25578 = t25577 ^ t25577;
    wire t25579 = t25578 ^ t25578;
    wire t25580 = t25579 ^ t25579;
    wire t25581 = t25580 ^ t25580;
    wire t25582 = t25581 ^ t25581;
    wire t25583 = t25582 ^ t25582;
    wire t25584 = t25583 ^ t25583;
    wire t25585 = t25584 ^ t25584;
    wire t25586 = t25585 ^ t25585;
    wire t25587 = t25586 ^ t25586;
    wire t25588 = t25587 ^ t25587;
    wire t25589 = t25588 ^ t25588;
    wire t25590 = t25589 ^ t25589;
    wire t25591 = t25590 ^ t25590;
    wire t25592 = t25591 ^ t25591;
    wire t25593 = t25592 ^ t25592;
    wire t25594 = t25593 ^ t25593;
    wire t25595 = t25594 ^ t25594;
    wire t25596 = t25595 ^ t25595;
    wire t25597 = t25596 ^ t25596;
    wire t25598 = t25597 ^ t25597;
    wire t25599 = t25598 ^ t25598;
    wire t25600 = t25599 ^ t25599;
    wire t25601 = t25600 ^ t25600;
    wire t25602 = t25601 ^ t25601;
    wire t25603 = t25602 ^ t25602;
    wire t25604 = t25603 ^ t25603;
    wire t25605 = t25604 ^ t25604;
    wire t25606 = t25605 ^ t25605;
    wire t25607 = t25606 ^ t25606;
    wire t25608 = t25607 ^ t25607;
    wire t25609 = t25608 ^ t25608;
    wire t25610 = t25609 ^ t25609;
    wire t25611 = t25610 ^ t25610;
    wire t25612 = t25611 ^ t25611;
    wire t25613 = t25612 ^ t25612;
    wire t25614 = t25613 ^ t25613;
    wire t25615 = t25614 ^ t25614;
    wire t25616 = t25615 ^ t25615;
    wire t25617 = t25616 ^ t25616;
    wire t25618 = t25617 ^ t25617;
    wire t25619 = t25618 ^ t25618;
    wire t25620 = t25619 ^ t25619;
    wire t25621 = t25620 ^ t25620;
    wire t25622 = t25621 ^ t25621;
    wire t25623 = t25622 ^ t25622;
    wire t25624 = t25623 ^ t25623;
    wire t25625 = t25624 ^ t25624;
    wire t25626 = t25625 ^ t25625;
    wire t25627 = t25626 ^ t25626;
    wire t25628 = t25627 ^ t25627;
    wire t25629 = t25628 ^ t25628;
    wire t25630 = t25629 ^ t25629;
    wire t25631 = t25630 ^ t25630;
    wire t25632 = t25631 ^ t25631;
    wire t25633 = t25632 ^ t25632;
    wire t25634 = t25633 ^ t25633;
    wire t25635 = t25634 ^ t25634;
    wire t25636 = t25635 ^ t25635;
    wire t25637 = t25636 ^ t25636;
    wire t25638 = t25637 ^ t25637;
    wire t25639 = t25638 ^ t25638;
    wire t25640 = t25639 ^ t25639;
    wire t25641 = t25640 ^ t25640;
    wire t25642 = t25641 ^ t25641;
    wire t25643 = t25642 ^ t25642;
    wire t25644 = t25643 ^ t25643;
    wire t25645 = t25644 ^ t25644;
    wire t25646 = t25645 ^ t25645;
    wire t25647 = t25646 ^ t25646;
    wire t25648 = t25647 ^ t25647;
    wire t25649 = t25648 ^ t25648;
    wire t25650 = t25649 ^ t25649;
    wire t25651 = t25650 ^ t25650;
    wire t25652 = t25651 ^ t25651;
    wire t25653 = t25652 ^ t25652;
    wire t25654 = t25653 ^ t25653;
    wire t25655 = t25654 ^ t25654;
    wire t25656 = t25655 ^ t25655;
    wire t25657 = t25656 ^ t25656;
    wire t25658 = t25657 ^ t25657;
    wire t25659 = t25658 ^ t25658;
    wire t25660 = t25659 ^ t25659;
    wire t25661 = t25660 ^ t25660;
    wire t25662 = t25661 ^ t25661;
    wire t25663 = t25662 ^ t25662;
    wire t25664 = t25663 ^ t25663;
    wire t25665 = t25664 ^ t25664;
    wire t25666 = t25665 ^ t25665;
    wire t25667 = t25666 ^ t25666;
    wire t25668 = t25667 ^ t25667;
    wire t25669 = t25668 ^ t25668;
    wire t25670 = t25669 ^ t25669;
    wire t25671 = t25670 ^ t25670;
    wire t25672 = t25671 ^ t25671;
    wire t25673 = t25672 ^ t25672;
    wire t25674 = t25673 ^ t25673;
    wire t25675 = t25674 ^ t25674;
    wire t25676 = t25675 ^ t25675;
    wire t25677 = t25676 ^ t25676;
    wire t25678 = t25677 ^ t25677;
    wire t25679 = t25678 ^ t25678;
    wire t25680 = t25679 ^ t25679;
    wire t25681 = t25680 ^ t25680;
    wire t25682 = t25681 ^ t25681;
    wire t25683 = t25682 ^ t25682;
    wire t25684 = t25683 ^ t25683;
    wire t25685 = t25684 ^ t25684;
    wire t25686 = t25685 ^ t25685;
    wire t25687 = t25686 ^ t25686;
    wire t25688 = t25687 ^ t25687;
    wire t25689 = t25688 ^ t25688;
    wire t25690 = t25689 ^ t25689;
    wire t25691 = t25690 ^ t25690;
    wire t25692 = t25691 ^ t25691;
    wire t25693 = t25692 ^ t25692;
    wire t25694 = t25693 ^ t25693;
    wire t25695 = t25694 ^ t25694;
    wire t25696 = t25695 ^ t25695;
    wire t25697 = t25696 ^ t25696;
    wire t25698 = t25697 ^ t25697;
    wire t25699 = t25698 ^ t25698;
    wire t25700 = t25699 ^ t25699;
    wire t25701 = t25700 ^ t25700;
    wire t25702 = t25701 ^ t25701;
    wire t25703 = t25702 ^ t25702;
    wire t25704 = t25703 ^ t25703;
    wire t25705 = t25704 ^ t25704;
    wire t25706 = t25705 ^ t25705;
    wire t25707 = t25706 ^ t25706;
    wire t25708 = t25707 ^ t25707;
    wire t25709 = t25708 ^ t25708;
    wire t25710 = t25709 ^ t25709;
    wire t25711 = t25710 ^ t25710;
    wire t25712 = t25711 ^ t25711;
    wire t25713 = t25712 ^ t25712;
    wire t25714 = t25713 ^ t25713;
    wire t25715 = t25714 ^ t25714;
    wire t25716 = t25715 ^ t25715;
    wire t25717 = t25716 ^ t25716;
    wire t25718 = t25717 ^ t25717;
    wire t25719 = t25718 ^ t25718;
    wire t25720 = t25719 ^ t25719;
    wire t25721 = t25720 ^ t25720;
    wire t25722 = t25721 ^ t25721;
    wire t25723 = t25722 ^ t25722;
    wire t25724 = t25723 ^ t25723;
    wire t25725 = t25724 ^ t25724;
    wire t25726 = t25725 ^ t25725;
    wire t25727 = t25726 ^ t25726;
    wire t25728 = t25727 ^ t25727;
    wire t25729 = t25728 ^ t25728;
    wire t25730 = t25729 ^ t25729;
    wire t25731 = t25730 ^ t25730;
    wire t25732 = t25731 ^ t25731;
    wire t25733 = t25732 ^ t25732;
    wire t25734 = t25733 ^ t25733;
    wire t25735 = t25734 ^ t25734;
    wire t25736 = t25735 ^ t25735;
    wire t25737 = t25736 ^ t25736;
    wire t25738 = t25737 ^ t25737;
    wire t25739 = t25738 ^ t25738;
    wire t25740 = t25739 ^ t25739;
    wire t25741 = t25740 ^ t25740;
    wire t25742 = t25741 ^ t25741;
    wire t25743 = t25742 ^ t25742;
    wire t25744 = t25743 ^ t25743;
    wire t25745 = t25744 ^ t25744;
    wire t25746 = t25745 ^ t25745;
    wire t25747 = t25746 ^ t25746;
    wire t25748 = t25747 ^ t25747;
    wire t25749 = t25748 ^ t25748;
    wire t25750 = t25749 ^ t25749;
    wire t25751 = t25750 ^ t25750;
    wire t25752 = t25751 ^ t25751;
    wire t25753 = t25752 ^ t25752;
    wire t25754 = t25753 ^ t25753;
    wire t25755 = t25754 ^ t25754;
    wire t25756 = t25755 ^ t25755;
    wire t25757 = t25756 ^ t25756;
    wire t25758 = t25757 ^ t25757;
    wire t25759 = t25758 ^ t25758;
    wire t25760 = t25759 ^ t25759;
    wire t25761 = t25760 ^ t25760;
    wire t25762 = t25761 ^ t25761;
    wire t25763 = t25762 ^ t25762;
    wire t25764 = t25763 ^ t25763;
    wire t25765 = t25764 ^ t25764;
    wire t25766 = t25765 ^ t25765;
    wire t25767 = t25766 ^ t25766;
    wire t25768 = t25767 ^ t25767;
    wire t25769 = t25768 ^ t25768;
    wire t25770 = t25769 ^ t25769;
    wire t25771 = t25770 ^ t25770;
    wire t25772 = t25771 ^ t25771;
    wire t25773 = t25772 ^ t25772;
    wire t25774 = t25773 ^ t25773;
    wire t25775 = t25774 ^ t25774;
    wire t25776 = t25775 ^ t25775;
    wire t25777 = t25776 ^ t25776;
    wire t25778 = t25777 ^ t25777;
    wire t25779 = t25778 ^ t25778;
    wire t25780 = t25779 ^ t25779;
    wire t25781 = t25780 ^ t25780;
    wire t25782 = t25781 ^ t25781;
    wire t25783 = t25782 ^ t25782;
    wire t25784 = t25783 ^ t25783;
    wire t25785 = t25784 ^ t25784;
    wire t25786 = t25785 ^ t25785;
    wire t25787 = t25786 ^ t25786;
    wire t25788 = t25787 ^ t25787;
    wire t25789 = t25788 ^ t25788;
    wire t25790 = t25789 ^ t25789;
    wire t25791 = t25790 ^ t25790;
    wire t25792 = t25791 ^ t25791;
    wire t25793 = t25792 ^ t25792;
    wire t25794 = t25793 ^ t25793;
    wire t25795 = t25794 ^ t25794;
    wire t25796 = t25795 ^ t25795;
    wire t25797 = t25796 ^ t25796;
    wire t25798 = t25797 ^ t25797;
    wire t25799 = t25798 ^ t25798;
    wire t25800 = t25799 ^ t25799;
    wire t25801 = t25800 ^ t25800;
    wire t25802 = t25801 ^ t25801;
    wire t25803 = t25802 ^ t25802;
    wire t25804 = t25803 ^ t25803;
    wire t25805 = t25804 ^ t25804;
    wire t25806 = t25805 ^ t25805;
    wire t25807 = t25806 ^ t25806;
    wire t25808 = t25807 ^ t25807;
    wire t25809 = t25808 ^ t25808;
    wire t25810 = t25809 ^ t25809;
    wire t25811 = t25810 ^ t25810;
    wire t25812 = t25811 ^ t25811;
    wire t25813 = t25812 ^ t25812;
    wire t25814 = t25813 ^ t25813;
    wire t25815 = t25814 ^ t25814;
    wire t25816 = t25815 ^ t25815;
    wire t25817 = t25816 ^ t25816;
    wire t25818 = t25817 ^ t25817;
    wire t25819 = t25818 ^ t25818;
    wire t25820 = t25819 ^ t25819;
    wire t25821 = t25820 ^ t25820;
    wire t25822 = t25821 ^ t25821;
    wire t25823 = t25822 ^ t25822;
    wire t25824 = t25823 ^ t25823;
    wire t25825 = t25824 ^ t25824;
    wire t25826 = t25825 ^ t25825;
    wire t25827 = t25826 ^ t25826;
    wire t25828 = t25827 ^ t25827;
    wire t25829 = t25828 ^ t25828;
    wire t25830 = t25829 ^ t25829;
    wire t25831 = t25830 ^ t25830;
    wire t25832 = t25831 ^ t25831;
    wire t25833 = t25832 ^ t25832;
    wire t25834 = t25833 ^ t25833;
    wire t25835 = t25834 ^ t25834;
    wire t25836 = t25835 ^ t25835;
    wire t25837 = t25836 ^ t25836;
    wire t25838 = t25837 ^ t25837;
    wire t25839 = t25838 ^ t25838;
    wire t25840 = t25839 ^ t25839;
    wire t25841 = t25840 ^ t25840;
    wire t25842 = t25841 ^ t25841;
    wire t25843 = t25842 ^ t25842;
    wire t25844 = t25843 ^ t25843;
    wire t25845 = t25844 ^ t25844;
    wire t25846 = t25845 ^ t25845;
    wire t25847 = t25846 ^ t25846;
    wire t25848 = t25847 ^ t25847;
    wire t25849 = t25848 ^ t25848;
    wire t25850 = t25849 ^ t25849;
    wire t25851 = t25850 ^ t25850;
    wire t25852 = t25851 ^ t25851;
    wire t25853 = t25852 ^ t25852;
    wire t25854 = t25853 ^ t25853;
    wire t25855 = t25854 ^ t25854;
    wire t25856 = t25855 ^ t25855;
    wire t25857 = t25856 ^ t25856;
    wire t25858 = t25857 ^ t25857;
    wire t25859 = t25858 ^ t25858;
    wire t25860 = t25859 ^ t25859;
    wire t25861 = t25860 ^ t25860;
    wire t25862 = t25861 ^ t25861;
    wire t25863 = t25862 ^ t25862;
    wire t25864 = t25863 ^ t25863;
    wire t25865 = t25864 ^ t25864;
    wire t25866 = t25865 ^ t25865;
    wire t25867 = t25866 ^ t25866;
    wire t25868 = t25867 ^ t25867;
    wire t25869 = t25868 ^ t25868;
    wire t25870 = t25869 ^ t25869;
    wire t25871 = t25870 ^ t25870;
    wire t25872 = t25871 ^ t25871;
    wire t25873 = t25872 ^ t25872;
    wire t25874 = t25873 ^ t25873;
    wire t25875 = t25874 ^ t25874;
    wire t25876 = t25875 ^ t25875;
    wire t25877 = t25876 ^ t25876;
    wire t25878 = t25877 ^ t25877;
    wire t25879 = t25878 ^ t25878;
    wire t25880 = t25879 ^ t25879;
    wire t25881 = t25880 ^ t25880;
    wire t25882 = t25881 ^ t25881;
    wire t25883 = t25882 ^ t25882;
    wire t25884 = t25883 ^ t25883;
    wire t25885 = t25884 ^ t25884;
    wire t25886 = t25885 ^ t25885;
    wire t25887 = t25886 ^ t25886;
    wire t25888 = t25887 ^ t25887;
    wire t25889 = t25888 ^ t25888;
    wire t25890 = t25889 ^ t25889;
    wire t25891 = t25890 ^ t25890;
    wire t25892 = t25891 ^ t25891;
    wire t25893 = t25892 ^ t25892;
    wire t25894 = t25893 ^ t25893;
    wire t25895 = t25894 ^ t25894;
    wire t25896 = t25895 ^ t25895;
    wire t25897 = t25896 ^ t25896;
    wire t25898 = t25897 ^ t25897;
    wire t25899 = t25898 ^ t25898;
    wire t25900 = t25899 ^ t25899;
    wire t25901 = t25900 ^ t25900;
    wire t25902 = t25901 ^ t25901;
    wire t25903 = t25902 ^ t25902;
    wire t25904 = t25903 ^ t25903;
    wire t25905 = t25904 ^ t25904;
    wire t25906 = t25905 ^ t25905;
    wire t25907 = t25906 ^ t25906;
    wire t25908 = t25907 ^ t25907;
    wire t25909 = t25908 ^ t25908;
    wire t25910 = t25909 ^ t25909;
    wire t25911 = t25910 ^ t25910;
    wire t25912 = t25911 ^ t25911;
    wire t25913 = t25912 ^ t25912;
    wire t25914 = t25913 ^ t25913;
    wire t25915 = t25914 ^ t25914;
    wire t25916 = t25915 ^ t25915;
    wire t25917 = t25916 ^ t25916;
    wire t25918 = t25917 ^ t25917;
    wire t25919 = t25918 ^ t25918;
    wire t25920 = t25919 ^ t25919;
    wire t25921 = t25920 ^ t25920;
    wire t25922 = t25921 ^ t25921;
    wire t25923 = t25922 ^ t25922;
    wire t25924 = t25923 ^ t25923;
    wire t25925 = t25924 ^ t25924;
    wire t25926 = t25925 ^ t25925;
    wire t25927 = t25926 ^ t25926;
    wire t25928 = t25927 ^ t25927;
    wire t25929 = t25928 ^ t25928;
    wire t25930 = t25929 ^ t25929;
    wire t25931 = t25930 ^ t25930;
    wire t25932 = t25931 ^ t25931;
    wire t25933 = t25932 ^ t25932;
    wire t25934 = t25933 ^ t25933;
    wire t25935 = t25934 ^ t25934;
    wire t25936 = t25935 ^ t25935;
    wire t25937 = t25936 ^ t25936;
    wire t25938 = t25937 ^ t25937;
    wire t25939 = t25938 ^ t25938;
    wire t25940 = t25939 ^ t25939;
    wire t25941 = t25940 ^ t25940;
    wire t25942 = t25941 ^ t25941;
    wire t25943 = t25942 ^ t25942;
    wire t25944 = t25943 ^ t25943;
    wire t25945 = t25944 ^ t25944;
    wire t25946 = t25945 ^ t25945;
    wire t25947 = t25946 ^ t25946;
    wire t25948 = t25947 ^ t25947;
    wire t25949 = t25948 ^ t25948;
    wire t25950 = t25949 ^ t25949;
    wire t25951 = t25950 ^ t25950;
    wire t25952 = t25951 ^ t25951;
    wire t25953 = t25952 ^ t25952;
    wire t25954 = t25953 ^ t25953;
    wire t25955 = t25954 ^ t25954;
    wire t25956 = t25955 ^ t25955;
    wire t25957 = t25956 ^ t25956;
    wire t25958 = t25957 ^ t25957;
    wire t25959 = t25958 ^ t25958;
    wire t25960 = t25959 ^ t25959;
    wire t25961 = t25960 ^ t25960;
    wire t25962 = t25961 ^ t25961;
    wire t25963 = t25962 ^ t25962;
    wire t25964 = t25963 ^ t25963;
    wire t25965 = t25964 ^ t25964;
    wire t25966 = t25965 ^ t25965;
    wire t25967 = t25966 ^ t25966;
    wire t25968 = t25967 ^ t25967;
    wire t25969 = t25968 ^ t25968;
    wire t25970 = t25969 ^ t25969;
    wire t25971 = t25970 ^ t25970;
    wire t25972 = t25971 ^ t25971;
    wire t25973 = t25972 ^ t25972;
    wire t25974 = t25973 ^ t25973;
    wire t25975 = t25974 ^ t25974;
    wire t25976 = t25975 ^ t25975;
    wire t25977 = t25976 ^ t25976;
    wire t25978 = t25977 ^ t25977;
    wire t25979 = t25978 ^ t25978;
    wire t25980 = t25979 ^ t25979;
    wire t25981 = t25980 ^ t25980;
    wire t25982 = t25981 ^ t25981;
    wire t25983 = t25982 ^ t25982;
    wire t25984 = t25983 ^ t25983;
    wire t25985 = t25984 ^ t25984;
    wire t25986 = t25985 ^ t25985;
    wire t25987 = t25986 ^ t25986;
    wire t25988 = t25987 ^ t25987;
    wire t25989 = t25988 ^ t25988;
    wire t25990 = t25989 ^ t25989;
    wire t25991 = t25990 ^ t25990;
    wire t25992 = t25991 ^ t25991;
    wire t25993 = t25992 ^ t25992;
    wire t25994 = t25993 ^ t25993;
    wire t25995 = t25994 ^ t25994;
    wire t25996 = t25995 ^ t25995;
    wire t25997 = t25996 ^ t25996;
    wire t25998 = t25997 ^ t25997;
    wire t25999 = t25998 ^ t25998;
    wire t26000 = t25999 ^ t25999;
    wire t26001 = t26000 ^ t26000;
    wire t26002 = t26001 ^ t26001;
    wire t26003 = t26002 ^ t26002;
    wire t26004 = t26003 ^ t26003;
    wire t26005 = t26004 ^ t26004;
    wire t26006 = t26005 ^ t26005;
    wire t26007 = t26006 ^ t26006;
    wire t26008 = t26007 ^ t26007;
    wire t26009 = t26008 ^ t26008;
    wire t26010 = t26009 ^ t26009;
    wire t26011 = t26010 ^ t26010;
    wire t26012 = t26011 ^ t26011;
    wire t26013 = t26012 ^ t26012;
    wire t26014 = t26013 ^ t26013;
    wire t26015 = t26014 ^ t26014;
    wire t26016 = t26015 ^ t26015;
    wire t26017 = t26016 ^ t26016;
    wire t26018 = t26017 ^ t26017;
    wire t26019 = t26018 ^ t26018;
    wire t26020 = t26019 ^ t26019;
    wire t26021 = t26020 ^ t26020;
    wire t26022 = t26021 ^ t26021;
    wire t26023 = t26022 ^ t26022;
    wire t26024 = t26023 ^ t26023;
    wire t26025 = t26024 ^ t26024;
    wire t26026 = t26025 ^ t26025;
    wire t26027 = t26026 ^ t26026;
    wire t26028 = t26027 ^ t26027;
    wire t26029 = t26028 ^ t26028;
    wire t26030 = t26029 ^ t26029;
    wire t26031 = t26030 ^ t26030;
    wire t26032 = t26031 ^ t26031;
    wire t26033 = t26032 ^ t26032;
    wire t26034 = t26033 ^ t26033;
    wire t26035 = t26034 ^ t26034;
    wire t26036 = t26035 ^ t26035;
    wire t26037 = t26036 ^ t26036;
    wire t26038 = t26037 ^ t26037;
    wire t26039 = t26038 ^ t26038;
    wire t26040 = t26039 ^ t26039;
    wire t26041 = t26040 ^ t26040;
    wire t26042 = t26041 ^ t26041;
    wire t26043 = t26042 ^ t26042;
    wire t26044 = t26043 ^ t26043;
    wire t26045 = t26044 ^ t26044;
    wire t26046 = t26045 ^ t26045;
    wire t26047 = t26046 ^ t26046;
    wire t26048 = t26047 ^ t26047;
    wire t26049 = t26048 ^ t26048;
    wire t26050 = t26049 ^ t26049;
    wire t26051 = t26050 ^ t26050;
    wire t26052 = t26051 ^ t26051;
    wire t26053 = t26052 ^ t26052;
    wire t26054 = t26053 ^ t26053;
    wire t26055 = t26054 ^ t26054;
    wire t26056 = t26055 ^ t26055;
    wire t26057 = t26056 ^ t26056;
    wire t26058 = t26057 ^ t26057;
    wire t26059 = t26058 ^ t26058;
    wire t26060 = t26059 ^ t26059;
    wire t26061 = t26060 ^ t26060;
    wire t26062 = t26061 ^ t26061;
    wire t26063 = t26062 ^ t26062;
    wire t26064 = t26063 ^ t26063;
    wire t26065 = t26064 ^ t26064;
    wire t26066 = t26065 ^ t26065;
    wire t26067 = t26066 ^ t26066;
    wire t26068 = t26067 ^ t26067;
    wire t26069 = t26068 ^ t26068;
    wire t26070 = t26069 ^ t26069;
    wire t26071 = t26070 ^ t26070;
    wire t26072 = t26071 ^ t26071;
    wire t26073 = t26072 ^ t26072;
    wire t26074 = t26073 ^ t26073;
    wire t26075 = t26074 ^ t26074;
    wire t26076 = t26075 ^ t26075;
    wire t26077 = t26076 ^ t26076;
    wire t26078 = t26077 ^ t26077;
    wire t26079 = t26078 ^ t26078;
    wire t26080 = t26079 ^ t26079;
    wire t26081 = t26080 ^ t26080;
    wire t26082 = t26081 ^ t26081;
    wire t26083 = t26082 ^ t26082;
    wire t26084 = t26083 ^ t26083;
    wire t26085 = t26084 ^ t26084;
    wire t26086 = t26085 ^ t26085;
    wire t26087 = t26086 ^ t26086;
    wire t26088 = t26087 ^ t26087;
    wire t26089 = t26088 ^ t26088;
    wire t26090 = t26089 ^ t26089;
    wire t26091 = t26090 ^ t26090;
    wire t26092 = t26091 ^ t26091;
    wire t26093 = t26092 ^ t26092;
    wire t26094 = t26093 ^ t26093;
    wire t26095 = t26094 ^ t26094;
    wire t26096 = t26095 ^ t26095;
    wire t26097 = t26096 ^ t26096;
    wire t26098 = t26097 ^ t26097;
    wire t26099 = t26098 ^ t26098;
    wire t26100 = t26099 ^ t26099;
    wire t26101 = t26100 ^ t26100;
    wire t26102 = t26101 ^ t26101;
    wire t26103 = t26102 ^ t26102;
    wire t26104 = t26103 ^ t26103;
    wire t26105 = t26104 ^ t26104;
    wire t26106 = t26105 ^ t26105;
    wire t26107 = t26106 ^ t26106;
    wire t26108 = t26107 ^ t26107;
    wire t26109 = t26108 ^ t26108;
    wire t26110 = t26109 ^ t26109;
    wire t26111 = t26110 ^ t26110;
    wire t26112 = t26111 ^ t26111;
    wire t26113 = t26112 ^ t26112;
    wire t26114 = t26113 ^ t26113;
    wire t26115 = t26114 ^ t26114;
    wire t26116 = t26115 ^ t26115;
    wire t26117 = t26116 ^ t26116;
    wire t26118 = t26117 ^ t26117;
    wire t26119 = t26118 ^ t26118;
    wire t26120 = t26119 ^ t26119;
    wire t26121 = t26120 ^ t26120;
    wire t26122 = t26121 ^ t26121;
    wire t26123 = t26122 ^ t26122;
    wire t26124 = t26123 ^ t26123;
    wire t26125 = t26124 ^ t26124;
    wire t26126 = t26125 ^ t26125;
    wire t26127 = t26126 ^ t26126;
    wire t26128 = t26127 ^ t26127;
    wire t26129 = t26128 ^ t26128;
    wire t26130 = t26129 ^ t26129;
    wire t26131 = t26130 ^ t26130;
    wire t26132 = t26131 ^ t26131;
    wire t26133 = t26132 ^ t26132;
    wire t26134 = t26133 ^ t26133;
    wire t26135 = t26134 ^ t26134;
    wire t26136 = t26135 ^ t26135;
    wire t26137 = t26136 ^ t26136;
    wire t26138 = t26137 ^ t26137;
    wire t26139 = t26138 ^ t26138;
    wire t26140 = t26139 ^ t26139;
    wire t26141 = t26140 ^ t26140;
    wire t26142 = t26141 ^ t26141;
    wire t26143 = t26142 ^ t26142;
    wire t26144 = t26143 ^ t26143;
    wire t26145 = t26144 ^ t26144;
    wire t26146 = t26145 ^ t26145;
    wire t26147 = t26146 ^ t26146;
    wire t26148 = t26147 ^ t26147;
    wire t26149 = t26148 ^ t26148;
    wire t26150 = t26149 ^ t26149;
    wire t26151 = t26150 ^ t26150;
    wire t26152 = t26151 ^ t26151;
    wire t26153 = t26152 ^ t26152;
    wire t26154 = t26153 ^ t26153;
    wire t26155 = t26154 ^ t26154;
    wire t26156 = t26155 ^ t26155;
    wire t26157 = t26156 ^ t26156;
    wire t26158 = t26157 ^ t26157;
    wire t26159 = t26158 ^ t26158;
    wire t26160 = t26159 ^ t26159;
    wire t26161 = t26160 ^ t26160;
    wire t26162 = t26161 ^ t26161;
    wire t26163 = t26162 ^ t26162;
    wire t26164 = t26163 ^ t26163;
    wire t26165 = t26164 ^ t26164;
    wire t26166 = t26165 ^ t26165;
    wire t26167 = t26166 ^ t26166;
    wire t26168 = t26167 ^ t26167;
    wire t26169 = t26168 ^ t26168;
    wire t26170 = t26169 ^ t26169;
    wire t26171 = t26170 ^ t26170;
    wire t26172 = t26171 ^ t26171;
    wire t26173 = t26172 ^ t26172;
    wire t26174 = t26173 ^ t26173;
    wire t26175 = t26174 ^ t26174;
    wire t26176 = t26175 ^ t26175;
    wire t26177 = t26176 ^ t26176;
    wire t26178 = t26177 ^ t26177;
    wire t26179 = t26178 ^ t26178;
    wire t26180 = t26179 ^ t26179;
    wire t26181 = t26180 ^ t26180;
    wire t26182 = t26181 ^ t26181;
    wire t26183 = t26182 ^ t26182;
    wire t26184 = t26183 ^ t26183;
    wire t26185 = t26184 ^ t26184;
    wire t26186 = t26185 ^ t26185;
    wire t26187 = t26186 ^ t26186;
    wire t26188 = t26187 ^ t26187;
    wire t26189 = t26188 ^ t26188;
    wire t26190 = t26189 ^ t26189;
    wire t26191 = t26190 ^ t26190;
    wire t26192 = t26191 ^ t26191;
    wire t26193 = t26192 ^ t26192;
    wire t26194 = t26193 ^ t26193;
    wire t26195 = t26194 ^ t26194;
    wire t26196 = t26195 ^ t26195;
    wire t26197 = t26196 ^ t26196;
    wire t26198 = t26197 ^ t26197;
    wire t26199 = t26198 ^ t26198;
    wire t26200 = t26199 ^ t26199;
    wire t26201 = t26200 ^ t26200;
    wire t26202 = t26201 ^ t26201;
    wire t26203 = t26202 ^ t26202;
    wire t26204 = t26203 ^ t26203;
    wire t26205 = t26204 ^ t26204;
    wire t26206 = t26205 ^ t26205;
    wire t26207 = t26206 ^ t26206;
    wire t26208 = t26207 ^ t26207;
    wire t26209 = t26208 ^ t26208;
    wire t26210 = t26209 ^ t26209;
    wire t26211 = t26210 ^ t26210;
    wire t26212 = t26211 ^ t26211;
    wire t26213 = t26212 ^ t26212;
    wire t26214 = t26213 ^ t26213;
    wire t26215 = t26214 ^ t26214;
    wire t26216 = t26215 ^ t26215;
    wire t26217 = t26216 ^ t26216;
    wire t26218 = t26217 ^ t26217;
    wire t26219 = t26218 ^ t26218;
    wire t26220 = t26219 ^ t26219;
    wire t26221 = t26220 ^ t26220;
    wire t26222 = t26221 ^ t26221;
    wire t26223 = t26222 ^ t26222;
    wire t26224 = t26223 ^ t26223;
    wire t26225 = t26224 ^ t26224;
    wire t26226 = t26225 ^ t26225;
    wire t26227 = t26226 ^ t26226;
    wire t26228 = t26227 ^ t26227;
    wire t26229 = t26228 ^ t26228;
    wire t26230 = t26229 ^ t26229;
    wire t26231 = t26230 ^ t26230;
    wire t26232 = t26231 ^ t26231;
    wire t26233 = t26232 ^ t26232;
    wire t26234 = t26233 ^ t26233;
    wire t26235 = t26234 ^ t26234;
    wire t26236 = t26235 ^ t26235;
    wire t26237 = t26236 ^ t26236;
    wire t26238 = t26237 ^ t26237;
    wire t26239 = t26238 ^ t26238;
    wire t26240 = t26239 ^ t26239;
    wire t26241 = t26240 ^ t26240;
    wire t26242 = t26241 ^ t26241;
    wire t26243 = t26242 ^ t26242;
    wire t26244 = t26243 ^ t26243;
    wire t26245 = t26244 ^ t26244;
    wire t26246 = t26245 ^ t26245;
    wire t26247 = t26246 ^ t26246;
    wire t26248 = t26247 ^ t26247;
    wire t26249 = t26248 ^ t26248;
    wire t26250 = t26249 ^ t26249;
    wire t26251 = t26250 ^ t26250;
    wire t26252 = t26251 ^ t26251;
    wire t26253 = t26252 ^ t26252;
    wire t26254 = t26253 ^ t26253;
    wire t26255 = t26254 ^ t26254;
    wire t26256 = t26255 ^ t26255;
    wire t26257 = t26256 ^ t26256;
    wire t26258 = t26257 ^ t26257;
    wire t26259 = t26258 ^ t26258;
    wire t26260 = t26259 ^ t26259;
    wire t26261 = t26260 ^ t26260;
    wire t26262 = t26261 ^ t26261;
    wire t26263 = t26262 ^ t26262;
    wire t26264 = t26263 ^ t26263;
    wire t26265 = t26264 ^ t26264;
    wire t26266 = t26265 ^ t26265;
    wire t26267 = t26266 ^ t26266;
    wire t26268 = t26267 ^ t26267;
    wire t26269 = t26268 ^ t26268;
    wire t26270 = t26269 ^ t26269;
    wire t26271 = t26270 ^ t26270;
    wire t26272 = t26271 ^ t26271;
    wire t26273 = t26272 ^ t26272;
    wire t26274 = t26273 ^ t26273;
    wire t26275 = t26274 ^ t26274;
    wire t26276 = t26275 ^ t26275;
    wire t26277 = t26276 ^ t26276;
    wire t26278 = t26277 ^ t26277;
    wire t26279 = t26278 ^ t26278;
    wire t26280 = t26279 ^ t26279;
    wire t26281 = t26280 ^ t26280;
    wire t26282 = t26281 ^ t26281;
    wire t26283 = t26282 ^ t26282;
    wire t26284 = t26283 ^ t26283;
    wire t26285 = t26284 ^ t26284;
    wire t26286 = t26285 ^ t26285;
    wire t26287 = t26286 ^ t26286;
    wire t26288 = t26287 ^ t26287;
    wire t26289 = t26288 ^ t26288;
    wire t26290 = t26289 ^ t26289;
    wire t26291 = t26290 ^ t26290;
    wire t26292 = t26291 ^ t26291;
    wire t26293 = t26292 ^ t26292;
    wire t26294 = t26293 ^ t26293;
    wire t26295 = t26294 ^ t26294;
    wire t26296 = t26295 ^ t26295;
    wire t26297 = t26296 ^ t26296;
    wire t26298 = t26297 ^ t26297;
    wire t26299 = t26298 ^ t26298;
    wire t26300 = t26299 ^ t26299;
    wire t26301 = t26300 ^ t26300;
    wire t26302 = t26301 ^ t26301;
    wire t26303 = t26302 ^ t26302;
    wire t26304 = t26303 ^ t26303;
    wire t26305 = t26304 ^ t26304;
    wire t26306 = t26305 ^ t26305;
    wire t26307 = t26306 ^ t26306;
    wire t26308 = t26307 ^ t26307;
    wire t26309 = t26308 ^ t26308;
    wire t26310 = t26309 ^ t26309;
    wire t26311 = t26310 ^ t26310;
    wire t26312 = t26311 ^ t26311;
    wire t26313 = t26312 ^ t26312;
    wire t26314 = t26313 ^ t26313;
    wire t26315 = t26314 ^ t26314;
    wire t26316 = t26315 ^ t26315;
    wire t26317 = t26316 ^ t26316;
    wire t26318 = t26317 ^ t26317;
    wire t26319 = t26318 ^ t26318;
    wire t26320 = t26319 ^ t26319;
    wire t26321 = t26320 ^ t26320;
    wire t26322 = t26321 ^ t26321;
    wire t26323 = t26322 ^ t26322;
    wire t26324 = t26323 ^ t26323;
    wire t26325 = t26324 ^ t26324;
    wire t26326 = t26325 ^ t26325;
    wire t26327 = t26326 ^ t26326;
    wire t26328 = t26327 ^ t26327;
    wire t26329 = t26328 ^ t26328;
    wire t26330 = t26329 ^ t26329;
    wire t26331 = t26330 ^ t26330;
    wire t26332 = t26331 ^ t26331;
    wire t26333 = t26332 ^ t26332;
    wire t26334 = t26333 ^ t26333;
    wire t26335 = t26334 ^ t26334;
    wire t26336 = t26335 ^ t26335;
    wire t26337 = t26336 ^ t26336;
    wire t26338 = t26337 ^ t26337;
    wire t26339 = t26338 ^ t26338;
    wire t26340 = t26339 ^ t26339;
    wire t26341 = t26340 ^ t26340;
    wire t26342 = t26341 ^ t26341;
    wire t26343 = t26342 ^ t26342;
    wire t26344 = t26343 ^ t26343;
    wire t26345 = t26344 ^ t26344;
    wire t26346 = t26345 ^ t26345;
    wire t26347 = t26346 ^ t26346;
    wire t26348 = t26347 ^ t26347;
    wire t26349 = t26348 ^ t26348;
    wire t26350 = t26349 ^ t26349;
    wire t26351 = t26350 ^ t26350;
    wire t26352 = t26351 ^ t26351;
    wire t26353 = t26352 ^ t26352;
    wire t26354 = t26353 ^ t26353;
    wire t26355 = t26354 ^ t26354;
    wire t26356 = t26355 ^ t26355;
    wire t26357 = t26356 ^ t26356;
    wire t26358 = t26357 ^ t26357;
    wire t26359 = t26358 ^ t26358;
    wire t26360 = t26359 ^ t26359;
    wire t26361 = t26360 ^ t26360;
    wire t26362 = t26361 ^ t26361;
    wire t26363 = t26362 ^ t26362;
    wire t26364 = t26363 ^ t26363;
    wire t26365 = t26364 ^ t26364;
    wire t26366 = t26365 ^ t26365;
    wire t26367 = t26366 ^ t26366;
    wire t26368 = t26367 ^ t26367;
    wire t26369 = t26368 ^ t26368;
    wire t26370 = t26369 ^ t26369;
    wire t26371 = t26370 ^ t26370;
    wire t26372 = t26371 ^ t26371;
    wire t26373 = t26372 ^ t26372;
    wire t26374 = t26373 ^ t26373;
    wire t26375 = t26374 ^ t26374;
    wire t26376 = t26375 ^ t26375;
    wire t26377 = t26376 ^ t26376;
    wire t26378 = t26377 ^ t26377;
    wire t26379 = t26378 ^ t26378;
    wire t26380 = t26379 ^ t26379;
    wire t26381 = t26380 ^ t26380;
    wire t26382 = t26381 ^ t26381;
    wire t26383 = t26382 ^ t26382;
    wire t26384 = t26383 ^ t26383;
    wire t26385 = t26384 ^ t26384;
    wire t26386 = t26385 ^ t26385;
    wire t26387 = t26386 ^ t26386;
    wire t26388 = t26387 ^ t26387;
    wire t26389 = t26388 ^ t26388;
    wire t26390 = t26389 ^ t26389;
    wire t26391 = t26390 ^ t26390;
    wire t26392 = t26391 ^ t26391;
    wire t26393 = t26392 ^ t26392;
    wire t26394 = t26393 ^ t26393;
    wire t26395 = t26394 ^ t26394;
    wire t26396 = t26395 ^ t26395;
    wire t26397 = t26396 ^ t26396;
    wire t26398 = t26397 ^ t26397;
    wire t26399 = t26398 ^ t26398;
    wire t26400 = t26399 ^ t26399;
    wire t26401 = t26400 ^ t26400;
    wire t26402 = t26401 ^ t26401;
    wire t26403 = t26402 ^ t26402;
    wire t26404 = t26403 ^ t26403;
    wire t26405 = t26404 ^ t26404;
    wire t26406 = t26405 ^ t26405;
    wire t26407 = t26406 ^ t26406;
    wire t26408 = t26407 ^ t26407;
    wire t26409 = t26408 ^ t26408;
    wire t26410 = t26409 ^ t26409;
    wire t26411 = t26410 ^ t26410;
    wire t26412 = t26411 ^ t26411;
    wire t26413 = t26412 ^ t26412;
    wire t26414 = t26413 ^ t26413;
    wire t26415 = t26414 ^ t26414;
    wire t26416 = t26415 ^ t26415;
    wire t26417 = t26416 ^ t26416;
    wire t26418 = t26417 ^ t26417;
    wire t26419 = t26418 ^ t26418;
    wire t26420 = t26419 ^ t26419;
    wire t26421 = t26420 ^ t26420;
    wire t26422 = t26421 ^ t26421;
    wire t26423 = t26422 ^ t26422;
    wire t26424 = t26423 ^ t26423;
    wire t26425 = t26424 ^ t26424;
    wire t26426 = t26425 ^ t26425;
    wire t26427 = t26426 ^ t26426;
    wire t26428 = t26427 ^ t26427;
    wire t26429 = t26428 ^ t26428;
    wire t26430 = t26429 ^ t26429;
    wire t26431 = t26430 ^ t26430;
    wire t26432 = t26431 ^ t26431;
    wire t26433 = t26432 ^ t26432;
    wire t26434 = t26433 ^ t26433;
    wire t26435 = t26434 ^ t26434;
    wire t26436 = t26435 ^ t26435;
    wire t26437 = t26436 ^ t26436;
    wire t26438 = t26437 ^ t26437;
    wire t26439 = t26438 ^ t26438;
    wire t26440 = t26439 ^ t26439;
    wire t26441 = t26440 ^ t26440;
    wire t26442 = t26441 ^ t26441;
    wire t26443 = t26442 ^ t26442;
    wire t26444 = t26443 ^ t26443;
    wire t26445 = t26444 ^ t26444;
    wire t26446 = t26445 ^ t26445;
    wire t26447 = t26446 ^ t26446;
    wire t26448 = t26447 ^ t26447;
    wire t26449 = t26448 ^ t26448;
    wire t26450 = t26449 ^ t26449;
    wire t26451 = t26450 ^ t26450;
    wire t26452 = t26451 ^ t26451;
    wire t26453 = t26452 ^ t26452;
    wire t26454 = t26453 ^ t26453;
    wire t26455 = t26454 ^ t26454;
    wire t26456 = t26455 ^ t26455;
    wire t26457 = t26456 ^ t26456;
    wire t26458 = t26457 ^ t26457;
    wire t26459 = t26458 ^ t26458;
    wire t26460 = t26459 ^ t26459;
    wire t26461 = t26460 ^ t26460;
    wire t26462 = t26461 ^ t26461;
    wire t26463 = t26462 ^ t26462;
    wire t26464 = t26463 ^ t26463;
    wire t26465 = t26464 ^ t26464;
    wire t26466 = t26465 ^ t26465;
    wire t26467 = t26466 ^ t26466;
    wire t26468 = t26467 ^ t26467;
    wire t26469 = t26468 ^ t26468;
    wire t26470 = t26469 ^ t26469;
    wire t26471 = t26470 ^ t26470;
    wire t26472 = t26471 ^ t26471;
    wire t26473 = t26472 ^ t26472;
    wire t26474 = t26473 ^ t26473;
    wire t26475 = t26474 ^ t26474;
    wire t26476 = t26475 ^ t26475;
    wire t26477 = t26476 ^ t26476;
    wire t26478 = t26477 ^ t26477;
    wire t26479 = t26478 ^ t26478;
    wire t26480 = t26479 ^ t26479;
    wire t26481 = t26480 ^ t26480;
    wire t26482 = t26481 ^ t26481;
    wire t26483 = t26482 ^ t26482;
    wire t26484 = t26483 ^ t26483;
    wire t26485 = t26484 ^ t26484;
    wire t26486 = t26485 ^ t26485;
    wire t26487 = t26486 ^ t26486;
    wire t26488 = t26487 ^ t26487;
    wire t26489 = t26488 ^ t26488;
    wire t26490 = t26489 ^ t26489;
    wire t26491 = t26490 ^ t26490;
    wire t26492 = t26491 ^ t26491;
    wire t26493 = t26492 ^ t26492;
    wire t26494 = t26493 ^ t26493;
    wire t26495 = t26494 ^ t26494;
    wire t26496 = t26495 ^ t26495;
    wire t26497 = t26496 ^ t26496;
    wire t26498 = t26497 ^ t26497;
    wire t26499 = t26498 ^ t26498;
    wire t26500 = t26499 ^ t26499;
    wire t26501 = t26500 ^ t26500;
    wire t26502 = t26501 ^ t26501;
    wire t26503 = t26502 ^ t26502;
    wire t26504 = t26503 ^ t26503;
    wire t26505 = t26504 ^ t26504;
    wire t26506 = t26505 ^ t26505;
    wire t26507 = t26506 ^ t26506;
    wire t26508 = t26507 ^ t26507;
    wire t26509 = t26508 ^ t26508;
    wire t26510 = t26509 ^ t26509;
    wire t26511 = t26510 ^ t26510;
    wire t26512 = t26511 ^ t26511;
    wire t26513 = t26512 ^ t26512;
    wire t26514 = t26513 ^ t26513;
    wire t26515 = t26514 ^ t26514;
    wire t26516 = t26515 ^ t26515;
    wire t26517 = t26516 ^ t26516;
    wire t26518 = t26517 ^ t26517;
    wire t26519 = t26518 ^ t26518;
    wire t26520 = t26519 ^ t26519;
    wire t26521 = t26520 ^ t26520;
    wire t26522 = t26521 ^ t26521;
    wire t26523 = t26522 ^ t26522;
    wire t26524 = t26523 ^ t26523;
    wire t26525 = t26524 ^ t26524;
    wire t26526 = t26525 ^ t26525;
    wire t26527 = t26526 ^ t26526;
    wire t26528 = t26527 ^ t26527;
    wire t26529 = t26528 ^ t26528;
    wire t26530 = t26529 ^ t26529;
    wire t26531 = t26530 ^ t26530;
    wire t26532 = t26531 ^ t26531;
    wire t26533 = t26532 ^ t26532;
    wire t26534 = t26533 ^ t26533;
    wire t26535 = t26534 ^ t26534;
    wire t26536 = t26535 ^ t26535;
    wire t26537 = t26536 ^ t26536;
    wire t26538 = t26537 ^ t26537;
    wire t26539 = t26538 ^ t26538;
    wire t26540 = t26539 ^ t26539;
    wire t26541 = t26540 ^ t26540;
    wire t26542 = t26541 ^ t26541;
    wire t26543 = t26542 ^ t26542;
    wire t26544 = t26543 ^ t26543;
    wire t26545 = t26544 ^ t26544;
    wire t26546 = t26545 ^ t26545;
    wire t26547 = t26546 ^ t26546;
    wire t26548 = t26547 ^ t26547;
    wire t26549 = t26548 ^ t26548;
    wire t26550 = t26549 ^ t26549;
    wire t26551 = t26550 ^ t26550;
    wire t26552 = t26551 ^ t26551;
    wire t26553 = t26552 ^ t26552;
    wire t26554 = t26553 ^ t26553;
    wire t26555 = t26554 ^ t26554;
    wire t26556 = t26555 ^ t26555;
    wire t26557 = t26556 ^ t26556;
    wire t26558 = t26557 ^ t26557;
    wire t26559 = t26558 ^ t26558;
    wire t26560 = t26559 ^ t26559;
    wire t26561 = t26560 ^ t26560;
    wire t26562 = t26561 ^ t26561;
    wire t26563 = t26562 ^ t26562;
    wire t26564 = t26563 ^ t26563;
    wire t26565 = t26564 ^ t26564;
    wire t26566 = t26565 ^ t26565;
    wire t26567 = t26566 ^ t26566;
    wire t26568 = t26567 ^ t26567;
    wire t26569 = t26568 ^ t26568;
    wire t26570 = t26569 ^ t26569;
    wire t26571 = t26570 ^ t26570;
    wire t26572 = t26571 ^ t26571;
    wire t26573 = t26572 ^ t26572;
    wire t26574 = t26573 ^ t26573;
    wire t26575 = t26574 ^ t26574;
    wire t26576 = t26575 ^ t26575;
    wire t26577 = t26576 ^ t26576;
    wire t26578 = t26577 ^ t26577;
    wire t26579 = t26578 ^ t26578;
    wire t26580 = t26579 ^ t26579;
    wire t26581 = t26580 ^ t26580;
    wire t26582 = t26581 ^ t26581;
    wire t26583 = t26582 ^ t26582;
    wire t26584 = t26583 ^ t26583;
    wire t26585 = t26584 ^ t26584;
    wire t26586 = t26585 ^ t26585;
    wire t26587 = t26586 ^ t26586;
    wire t26588 = t26587 ^ t26587;
    wire t26589 = t26588 ^ t26588;
    wire t26590 = t26589 ^ t26589;
    wire t26591 = t26590 ^ t26590;
    wire t26592 = t26591 ^ t26591;
    wire t26593 = t26592 ^ t26592;
    wire t26594 = t26593 ^ t26593;
    wire t26595 = t26594 ^ t26594;
    wire t26596 = t26595 ^ t26595;
    wire t26597 = t26596 ^ t26596;
    wire t26598 = t26597 ^ t26597;
    wire t26599 = t26598 ^ t26598;
    wire t26600 = t26599 ^ t26599;
    wire t26601 = t26600 ^ t26600;
    wire t26602 = t26601 ^ t26601;
    wire t26603 = t26602 ^ t26602;
    wire t26604 = t26603 ^ t26603;
    wire t26605 = t26604 ^ t26604;
    wire t26606 = t26605 ^ t26605;
    wire t26607 = t26606 ^ t26606;
    wire t26608 = t26607 ^ t26607;
    wire t26609 = t26608 ^ t26608;
    wire t26610 = t26609 ^ t26609;
    wire t26611 = t26610 ^ t26610;
    wire t26612 = t26611 ^ t26611;
    wire t26613 = t26612 ^ t26612;
    wire t26614 = t26613 ^ t26613;
    wire t26615 = t26614 ^ t26614;
    wire t26616 = t26615 ^ t26615;
    wire t26617 = t26616 ^ t26616;
    wire t26618 = t26617 ^ t26617;
    wire t26619 = t26618 ^ t26618;
    wire t26620 = t26619 ^ t26619;
    wire t26621 = t26620 ^ t26620;
    wire t26622 = t26621 ^ t26621;
    wire t26623 = t26622 ^ t26622;
    wire t26624 = t26623 ^ t26623;
    wire t26625 = t26624 ^ t26624;
    wire t26626 = t26625 ^ t26625;
    wire t26627 = t26626 ^ t26626;
    wire t26628 = t26627 ^ t26627;
    wire t26629 = t26628 ^ t26628;
    wire t26630 = t26629 ^ t26629;
    wire t26631 = t26630 ^ t26630;
    wire t26632 = t26631 ^ t26631;
    wire t26633 = t26632 ^ t26632;
    wire t26634 = t26633 ^ t26633;
    wire t26635 = t26634 ^ t26634;
    wire t26636 = t26635 ^ t26635;
    wire t26637 = t26636 ^ t26636;
    wire t26638 = t26637 ^ t26637;
    wire t26639 = t26638 ^ t26638;
    wire t26640 = t26639 ^ t26639;
    wire t26641 = t26640 ^ t26640;
    wire t26642 = t26641 ^ t26641;
    wire t26643 = t26642 ^ t26642;
    wire t26644 = t26643 ^ t26643;
    wire t26645 = t26644 ^ t26644;
    wire t26646 = t26645 ^ t26645;
    wire t26647 = t26646 ^ t26646;
    wire t26648 = t26647 ^ t26647;
    wire t26649 = t26648 ^ t26648;
    wire t26650 = t26649 ^ t26649;
    wire t26651 = t26650 ^ t26650;
    wire t26652 = t26651 ^ t26651;
    wire t26653 = t26652 ^ t26652;
    wire t26654 = t26653 ^ t26653;
    wire t26655 = t26654 ^ t26654;
    wire t26656 = t26655 ^ t26655;
    wire t26657 = t26656 ^ t26656;
    wire t26658 = t26657 ^ t26657;
    wire t26659 = t26658 ^ t26658;
    wire t26660 = t26659 ^ t26659;
    wire t26661 = t26660 ^ t26660;
    wire t26662 = t26661 ^ t26661;
    wire t26663 = t26662 ^ t26662;
    wire t26664 = t26663 ^ t26663;
    wire t26665 = t26664 ^ t26664;
    wire t26666 = t26665 ^ t26665;
    wire t26667 = t26666 ^ t26666;
    wire t26668 = t26667 ^ t26667;
    wire t26669 = t26668 ^ t26668;
    wire t26670 = t26669 ^ t26669;
    wire t26671 = t26670 ^ t26670;
    wire t26672 = t26671 ^ t26671;
    wire t26673 = t26672 ^ t26672;
    wire t26674 = t26673 ^ t26673;
    wire t26675 = t26674 ^ t26674;
    wire t26676 = t26675 ^ t26675;
    wire t26677 = t26676 ^ t26676;
    wire t26678 = t26677 ^ t26677;
    wire t26679 = t26678 ^ t26678;
    wire t26680 = t26679 ^ t26679;
    wire t26681 = t26680 ^ t26680;
    wire t26682 = t26681 ^ t26681;
    wire t26683 = t26682 ^ t26682;
    wire t26684 = t26683 ^ t26683;
    wire t26685 = t26684 ^ t26684;
    wire t26686 = t26685 ^ t26685;
    wire t26687 = t26686 ^ t26686;
    wire t26688 = t26687 ^ t26687;
    wire t26689 = t26688 ^ t26688;
    wire t26690 = t26689 ^ t26689;
    wire t26691 = t26690 ^ t26690;
    wire t26692 = t26691 ^ t26691;
    wire t26693 = t26692 ^ t26692;
    wire t26694 = t26693 ^ t26693;
    wire t26695 = t26694 ^ t26694;
    wire t26696 = t26695 ^ t26695;
    wire t26697 = t26696 ^ t26696;
    wire t26698 = t26697 ^ t26697;
    wire t26699 = t26698 ^ t26698;
    wire t26700 = t26699 ^ t26699;
    wire t26701 = t26700 ^ t26700;
    wire t26702 = t26701 ^ t26701;
    wire t26703 = t26702 ^ t26702;
    wire t26704 = t26703 ^ t26703;
    wire t26705 = t26704 ^ t26704;
    wire t26706 = t26705 ^ t26705;
    wire t26707 = t26706 ^ t26706;
    wire t26708 = t26707 ^ t26707;
    wire t26709 = t26708 ^ t26708;
    wire t26710 = t26709 ^ t26709;
    wire t26711 = t26710 ^ t26710;
    wire t26712 = t26711 ^ t26711;
    wire t26713 = t26712 ^ t26712;
    wire t26714 = t26713 ^ t26713;
    wire t26715 = t26714 ^ t26714;
    wire t26716 = t26715 ^ t26715;
    wire t26717 = t26716 ^ t26716;
    wire t26718 = t26717 ^ t26717;
    wire t26719 = t26718 ^ t26718;
    wire t26720 = t26719 ^ t26719;
    wire t26721 = t26720 ^ t26720;
    wire t26722 = t26721 ^ t26721;
    wire t26723 = t26722 ^ t26722;
    wire t26724 = t26723 ^ t26723;
    wire t26725 = t26724 ^ t26724;
    wire t26726 = t26725 ^ t26725;
    wire t26727 = t26726 ^ t26726;
    wire t26728 = t26727 ^ t26727;
    wire t26729 = t26728 ^ t26728;
    wire t26730 = t26729 ^ t26729;
    wire t26731 = t26730 ^ t26730;
    wire t26732 = t26731 ^ t26731;
    wire t26733 = t26732 ^ t26732;
    wire t26734 = t26733 ^ t26733;
    wire t26735 = t26734 ^ t26734;
    wire t26736 = t26735 ^ t26735;
    wire t26737 = t26736 ^ t26736;
    wire t26738 = t26737 ^ t26737;
    wire t26739 = t26738 ^ t26738;
    wire t26740 = t26739 ^ t26739;
    wire t26741 = t26740 ^ t26740;
    wire t26742 = t26741 ^ t26741;
    wire t26743 = t26742 ^ t26742;
    wire t26744 = t26743 ^ t26743;
    wire t26745 = t26744 ^ t26744;
    wire t26746 = t26745 ^ t26745;
    wire t26747 = t26746 ^ t26746;
    wire t26748 = t26747 ^ t26747;
    wire t26749 = t26748 ^ t26748;
    wire t26750 = t26749 ^ t26749;
    wire t26751 = t26750 ^ t26750;
    wire t26752 = t26751 ^ t26751;
    wire t26753 = t26752 ^ t26752;
    wire t26754 = t26753 ^ t26753;
    wire t26755 = t26754 ^ t26754;
    wire t26756 = t26755 ^ t26755;
    wire t26757 = t26756 ^ t26756;
    wire t26758 = t26757 ^ t26757;
    wire t26759 = t26758 ^ t26758;
    wire t26760 = t26759 ^ t26759;
    wire t26761 = t26760 ^ t26760;
    wire t26762 = t26761 ^ t26761;
    wire t26763 = t26762 ^ t26762;
    wire t26764 = t26763 ^ t26763;
    wire t26765 = t26764 ^ t26764;
    wire t26766 = t26765 ^ t26765;
    wire t26767 = t26766 ^ t26766;
    wire t26768 = t26767 ^ t26767;
    wire t26769 = t26768 ^ t26768;
    wire t26770 = t26769 ^ t26769;
    wire t26771 = t26770 ^ t26770;
    wire t26772 = t26771 ^ t26771;
    wire t26773 = t26772 ^ t26772;
    wire t26774 = t26773 ^ t26773;
    wire t26775 = t26774 ^ t26774;
    wire t26776 = t26775 ^ t26775;
    wire t26777 = t26776 ^ t26776;
    wire t26778 = t26777 ^ t26777;
    wire t26779 = t26778 ^ t26778;
    wire t26780 = t26779 ^ t26779;
    wire t26781 = t26780 ^ t26780;
    wire t26782 = t26781 ^ t26781;
    wire t26783 = t26782 ^ t26782;
    wire t26784 = t26783 ^ t26783;
    wire t26785 = t26784 ^ t26784;
    wire t26786 = t26785 ^ t26785;
    wire t26787 = t26786 ^ t26786;
    wire t26788 = t26787 ^ t26787;
    wire t26789 = t26788 ^ t26788;
    wire t26790 = t26789 ^ t26789;
    wire t26791 = t26790 ^ t26790;
    wire t26792 = t26791 ^ t26791;
    wire t26793 = t26792 ^ t26792;
    wire t26794 = t26793 ^ t26793;
    wire t26795 = t26794 ^ t26794;
    wire t26796 = t26795 ^ t26795;
    wire t26797 = t26796 ^ t26796;
    wire t26798 = t26797 ^ t26797;
    wire t26799 = t26798 ^ t26798;
    wire t26800 = t26799 ^ t26799;
    wire t26801 = t26800 ^ t26800;
    wire t26802 = t26801 ^ t26801;
    wire t26803 = t26802 ^ t26802;
    wire t26804 = t26803 ^ t26803;
    wire t26805 = t26804 ^ t26804;
    wire t26806 = t26805 ^ t26805;
    wire t26807 = t26806 ^ t26806;
    wire t26808 = t26807 ^ t26807;
    wire t26809 = t26808 ^ t26808;
    wire t26810 = t26809 ^ t26809;
    wire t26811 = t26810 ^ t26810;
    wire t26812 = t26811 ^ t26811;
    wire t26813 = t26812 ^ t26812;
    wire t26814 = t26813 ^ t26813;
    wire t26815 = t26814 ^ t26814;
    wire t26816 = t26815 ^ t26815;
    wire t26817 = t26816 ^ t26816;
    wire t26818 = t26817 ^ t26817;
    wire t26819 = t26818 ^ t26818;
    wire t26820 = t26819 ^ t26819;
    wire t26821 = t26820 ^ t26820;
    wire t26822 = t26821 ^ t26821;
    wire t26823 = t26822 ^ t26822;
    wire t26824 = t26823 ^ t26823;
    wire t26825 = t26824 ^ t26824;
    wire t26826 = t26825 ^ t26825;
    wire t26827 = t26826 ^ t26826;
    wire t26828 = t26827 ^ t26827;
    wire t26829 = t26828 ^ t26828;
    wire t26830 = t26829 ^ t26829;
    wire t26831 = t26830 ^ t26830;
    wire t26832 = t26831 ^ t26831;
    wire t26833 = t26832 ^ t26832;
    wire t26834 = t26833 ^ t26833;
    wire t26835 = t26834 ^ t26834;
    wire t26836 = t26835 ^ t26835;
    wire t26837 = t26836 ^ t26836;
    wire t26838 = t26837 ^ t26837;
    wire t26839 = t26838 ^ t26838;
    wire t26840 = t26839 ^ t26839;
    wire t26841 = t26840 ^ t26840;
    wire t26842 = t26841 ^ t26841;
    wire t26843 = t26842 ^ t26842;
    wire t26844 = t26843 ^ t26843;
    wire t26845 = t26844 ^ t26844;
    wire t26846 = t26845 ^ t26845;
    wire t26847 = t26846 ^ t26846;
    wire t26848 = t26847 ^ t26847;
    wire t26849 = t26848 ^ t26848;
    wire t26850 = t26849 ^ t26849;
    wire t26851 = t26850 ^ t26850;
    wire t26852 = t26851 ^ t26851;
    wire t26853 = t26852 ^ t26852;
    wire t26854 = t26853 ^ t26853;
    wire t26855 = t26854 ^ t26854;
    wire t26856 = t26855 ^ t26855;
    wire t26857 = t26856 ^ t26856;
    wire t26858 = t26857 ^ t26857;
    wire t26859 = t26858 ^ t26858;
    wire t26860 = t26859 ^ t26859;
    wire t26861 = t26860 ^ t26860;
    wire t26862 = t26861 ^ t26861;
    wire t26863 = t26862 ^ t26862;
    wire t26864 = t26863 ^ t26863;
    wire t26865 = t26864 ^ t26864;
    wire t26866 = t26865 ^ t26865;
    wire t26867 = t26866 ^ t26866;
    wire t26868 = t26867 ^ t26867;
    wire t26869 = t26868 ^ t26868;
    wire t26870 = t26869 ^ t26869;
    wire t26871 = t26870 ^ t26870;
    wire t26872 = t26871 ^ t26871;
    wire t26873 = t26872 ^ t26872;
    wire t26874 = t26873 ^ t26873;
    wire t26875 = t26874 ^ t26874;
    wire t26876 = t26875 ^ t26875;
    wire t26877 = t26876 ^ t26876;
    wire t26878 = t26877 ^ t26877;
    wire t26879 = t26878 ^ t26878;
    wire t26880 = t26879 ^ t26879;
    wire t26881 = t26880 ^ t26880;
    wire t26882 = t26881 ^ t26881;
    wire t26883 = t26882 ^ t26882;
    wire t26884 = t26883 ^ t26883;
    wire t26885 = t26884 ^ t26884;
    wire t26886 = t26885 ^ t26885;
    wire t26887 = t26886 ^ t26886;
    wire t26888 = t26887 ^ t26887;
    wire t26889 = t26888 ^ t26888;
    wire t26890 = t26889 ^ t26889;
    wire t26891 = t26890 ^ t26890;
    wire t26892 = t26891 ^ t26891;
    wire t26893 = t26892 ^ t26892;
    wire t26894 = t26893 ^ t26893;
    wire t26895 = t26894 ^ t26894;
    wire t26896 = t26895 ^ t26895;
    wire t26897 = t26896 ^ t26896;
    wire t26898 = t26897 ^ t26897;
    wire t26899 = t26898 ^ t26898;
    wire t26900 = t26899 ^ t26899;
    wire t26901 = t26900 ^ t26900;
    wire t26902 = t26901 ^ t26901;
    wire t26903 = t26902 ^ t26902;
    wire t26904 = t26903 ^ t26903;
    wire t26905 = t26904 ^ t26904;
    wire t26906 = t26905 ^ t26905;
    wire t26907 = t26906 ^ t26906;
    wire t26908 = t26907 ^ t26907;
    wire t26909 = t26908 ^ t26908;
    wire t26910 = t26909 ^ t26909;
    wire t26911 = t26910 ^ t26910;
    wire t26912 = t26911 ^ t26911;
    wire t26913 = t26912 ^ t26912;
    wire t26914 = t26913 ^ t26913;
    wire t26915 = t26914 ^ t26914;
    wire t26916 = t26915 ^ t26915;
    wire t26917 = t26916 ^ t26916;
    wire t26918 = t26917 ^ t26917;
    wire t26919 = t26918 ^ t26918;
    wire t26920 = t26919 ^ t26919;
    wire t26921 = t26920 ^ t26920;
    wire t26922 = t26921 ^ t26921;
    wire t26923 = t26922 ^ t26922;
    wire t26924 = t26923 ^ t26923;
    wire t26925 = t26924 ^ t26924;
    wire t26926 = t26925 ^ t26925;
    wire t26927 = t26926 ^ t26926;
    wire t26928 = t26927 ^ t26927;
    wire t26929 = t26928 ^ t26928;
    wire t26930 = t26929 ^ t26929;
    wire t26931 = t26930 ^ t26930;
    wire t26932 = t26931 ^ t26931;
    wire t26933 = t26932 ^ t26932;
    wire t26934 = t26933 ^ t26933;
    wire t26935 = t26934 ^ t26934;
    wire t26936 = t26935 ^ t26935;
    wire t26937 = t26936 ^ t26936;
    wire t26938 = t26937 ^ t26937;
    wire t26939 = t26938 ^ t26938;
    wire t26940 = t26939 ^ t26939;
    wire t26941 = t26940 ^ t26940;
    wire t26942 = t26941 ^ t26941;
    wire t26943 = t26942 ^ t26942;
    wire t26944 = t26943 ^ t26943;
    wire t26945 = t26944 ^ t26944;
    wire t26946 = t26945 ^ t26945;
    wire t26947 = t26946 ^ t26946;
    wire t26948 = t26947 ^ t26947;
    wire t26949 = t26948 ^ t26948;
    wire t26950 = t26949 ^ t26949;
    wire t26951 = t26950 ^ t26950;
    wire t26952 = t26951 ^ t26951;
    wire t26953 = t26952 ^ t26952;
    wire t26954 = t26953 ^ t26953;
    wire t26955 = t26954 ^ t26954;
    wire t26956 = t26955 ^ t26955;
    wire t26957 = t26956 ^ t26956;
    wire t26958 = t26957 ^ t26957;
    wire t26959 = t26958 ^ t26958;
    wire t26960 = t26959 ^ t26959;
    wire t26961 = t26960 ^ t26960;
    wire t26962 = t26961 ^ t26961;
    wire t26963 = t26962 ^ t26962;
    wire t26964 = t26963 ^ t26963;
    wire t26965 = t26964 ^ t26964;
    wire t26966 = t26965 ^ t26965;
    wire t26967 = t26966 ^ t26966;
    wire t26968 = t26967 ^ t26967;
    wire t26969 = t26968 ^ t26968;
    wire t26970 = t26969 ^ t26969;
    wire t26971 = t26970 ^ t26970;
    wire t26972 = t26971 ^ t26971;
    wire t26973 = t26972 ^ t26972;
    wire t26974 = t26973 ^ t26973;
    wire t26975 = t26974 ^ t26974;
    wire t26976 = t26975 ^ t26975;
    wire t26977 = t26976 ^ t26976;
    wire t26978 = t26977 ^ t26977;
    wire t26979 = t26978 ^ t26978;
    wire t26980 = t26979 ^ t26979;
    wire t26981 = t26980 ^ t26980;
    wire t26982 = t26981 ^ t26981;
    wire t26983 = t26982 ^ t26982;
    wire t26984 = t26983 ^ t26983;
    wire t26985 = t26984 ^ t26984;
    wire t26986 = t26985 ^ t26985;
    wire t26987 = t26986 ^ t26986;
    wire t26988 = t26987 ^ t26987;
    wire t26989 = t26988 ^ t26988;
    wire t26990 = t26989 ^ t26989;
    wire t26991 = t26990 ^ t26990;
    wire t26992 = t26991 ^ t26991;
    wire t26993 = t26992 ^ t26992;
    wire t26994 = t26993 ^ t26993;
    wire t26995 = t26994 ^ t26994;
    wire t26996 = t26995 ^ t26995;
    wire t26997 = t26996 ^ t26996;
    wire t26998 = t26997 ^ t26997;
    wire t26999 = t26998 ^ t26998;
    wire t27000 = t26999 ^ t26999;
    wire t27001 = t27000 ^ t27000;
    wire t27002 = t27001 ^ t27001;
    wire t27003 = t27002 ^ t27002;
    wire t27004 = t27003 ^ t27003;
    wire t27005 = t27004 ^ t27004;
    wire t27006 = t27005 ^ t27005;
    wire t27007 = t27006 ^ t27006;
    wire t27008 = t27007 ^ t27007;
    wire t27009 = t27008 ^ t27008;
    wire t27010 = t27009 ^ t27009;
    wire t27011 = t27010 ^ t27010;
    wire t27012 = t27011 ^ t27011;
    wire t27013 = t27012 ^ t27012;
    wire t27014 = t27013 ^ t27013;
    wire t27015 = t27014 ^ t27014;
    wire t27016 = t27015 ^ t27015;
    wire t27017 = t27016 ^ t27016;
    wire t27018 = t27017 ^ t27017;
    wire t27019 = t27018 ^ t27018;
    wire t27020 = t27019 ^ t27019;
    wire t27021 = t27020 ^ t27020;
    wire t27022 = t27021 ^ t27021;
    wire t27023 = t27022 ^ t27022;
    wire t27024 = t27023 ^ t27023;
    wire t27025 = t27024 ^ t27024;
    wire t27026 = t27025 ^ t27025;
    wire t27027 = t27026 ^ t27026;
    wire t27028 = t27027 ^ t27027;
    wire t27029 = t27028 ^ t27028;
    wire t27030 = t27029 ^ t27029;
    wire t27031 = t27030 ^ t27030;
    wire t27032 = t27031 ^ t27031;
    wire t27033 = t27032 ^ t27032;
    wire t27034 = t27033 ^ t27033;
    wire t27035 = t27034 ^ t27034;
    wire t27036 = t27035 ^ t27035;
    wire t27037 = t27036 ^ t27036;
    wire t27038 = t27037 ^ t27037;
    wire t27039 = t27038 ^ t27038;
    wire t27040 = t27039 ^ t27039;
    wire t27041 = t27040 ^ t27040;
    wire t27042 = t27041 ^ t27041;
    wire t27043 = t27042 ^ t27042;
    wire t27044 = t27043 ^ t27043;
    wire t27045 = t27044 ^ t27044;
    wire t27046 = t27045 ^ t27045;
    wire t27047 = t27046 ^ t27046;
    wire t27048 = t27047 ^ t27047;
    wire t27049 = t27048 ^ t27048;
    wire t27050 = t27049 ^ t27049;
    wire t27051 = t27050 ^ t27050;
    wire t27052 = t27051 ^ t27051;
    wire t27053 = t27052 ^ t27052;
    wire t27054 = t27053 ^ t27053;
    wire t27055 = t27054 ^ t27054;
    wire t27056 = t27055 ^ t27055;
    wire t27057 = t27056 ^ t27056;
    wire t27058 = t27057 ^ t27057;
    wire t27059 = t27058 ^ t27058;
    wire t27060 = t27059 ^ t27059;
    wire t27061 = t27060 ^ t27060;
    wire t27062 = t27061 ^ t27061;
    wire t27063 = t27062 ^ t27062;
    wire t27064 = t27063 ^ t27063;
    wire t27065 = t27064 ^ t27064;
    wire t27066 = t27065 ^ t27065;
    wire t27067 = t27066 ^ t27066;
    wire t27068 = t27067 ^ t27067;
    wire t27069 = t27068 ^ t27068;
    wire t27070 = t27069 ^ t27069;
    wire t27071 = t27070 ^ t27070;
    wire t27072 = t27071 ^ t27071;
    wire t27073 = t27072 ^ t27072;
    wire t27074 = t27073 ^ t27073;
    wire t27075 = t27074 ^ t27074;
    wire t27076 = t27075 ^ t27075;
    wire t27077 = t27076 ^ t27076;
    wire t27078 = t27077 ^ t27077;
    wire t27079 = t27078 ^ t27078;
    wire t27080 = t27079 ^ t27079;
    wire t27081 = t27080 ^ t27080;
    wire t27082 = t27081 ^ t27081;
    wire t27083 = t27082 ^ t27082;
    wire t27084 = t27083 ^ t27083;
    wire t27085 = t27084 ^ t27084;
    wire t27086 = t27085 ^ t27085;
    wire t27087 = t27086 ^ t27086;
    wire t27088 = t27087 ^ t27087;
    wire t27089 = t27088 ^ t27088;
    wire t27090 = t27089 ^ t27089;
    wire t27091 = t27090 ^ t27090;
    wire t27092 = t27091 ^ t27091;
    wire t27093 = t27092 ^ t27092;
    wire t27094 = t27093 ^ t27093;
    wire t27095 = t27094 ^ t27094;
    wire t27096 = t27095 ^ t27095;
    wire t27097 = t27096 ^ t27096;
    wire t27098 = t27097 ^ t27097;
    wire t27099 = t27098 ^ t27098;
    wire t27100 = t27099 ^ t27099;
    wire t27101 = t27100 ^ t27100;
    wire t27102 = t27101 ^ t27101;
    wire t27103 = t27102 ^ t27102;
    wire t27104 = t27103 ^ t27103;
    wire t27105 = t27104 ^ t27104;
    wire t27106 = t27105 ^ t27105;
    wire t27107 = t27106 ^ t27106;
    wire t27108 = t27107 ^ t27107;
    wire t27109 = t27108 ^ t27108;
    wire t27110 = t27109 ^ t27109;
    wire t27111 = t27110 ^ t27110;
    wire t27112 = t27111 ^ t27111;
    wire t27113 = t27112 ^ t27112;
    wire t27114 = t27113 ^ t27113;
    wire t27115 = t27114 ^ t27114;
    wire t27116 = t27115 ^ t27115;
    wire t27117 = t27116 ^ t27116;
    wire t27118 = t27117 ^ t27117;
    wire t27119 = t27118 ^ t27118;
    wire t27120 = t27119 ^ t27119;
    wire t27121 = t27120 ^ t27120;
    wire t27122 = t27121 ^ t27121;
    wire t27123 = t27122 ^ t27122;
    wire t27124 = t27123 ^ t27123;
    wire t27125 = t27124 ^ t27124;
    wire t27126 = t27125 ^ t27125;
    wire t27127 = t27126 ^ t27126;
    wire t27128 = t27127 ^ t27127;
    wire t27129 = t27128 ^ t27128;
    wire t27130 = t27129 ^ t27129;
    wire t27131 = t27130 ^ t27130;
    wire t27132 = t27131 ^ t27131;
    wire t27133 = t27132 ^ t27132;
    wire t27134 = t27133 ^ t27133;
    wire t27135 = t27134 ^ t27134;
    wire t27136 = t27135 ^ t27135;
    wire t27137 = t27136 ^ t27136;
    wire t27138 = t27137 ^ t27137;
    wire t27139 = t27138 ^ t27138;
    wire t27140 = t27139 ^ t27139;
    wire t27141 = t27140 ^ t27140;
    wire t27142 = t27141 ^ t27141;
    wire t27143 = t27142 ^ t27142;
    wire t27144 = t27143 ^ t27143;
    wire t27145 = t27144 ^ t27144;
    wire t27146 = t27145 ^ t27145;
    wire t27147 = t27146 ^ t27146;
    wire t27148 = t27147 ^ t27147;
    wire t27149 = t27148 ^ t27148;
    wire t27150 = t27149 ^ t27149;
    wire t27151 = t27150 ^ t27150;
    wire t27152 = t27151 ^ t27151;
    wire t27153 = t27152 ^ t27152;
    wire t27154 = t27153 ^ t27153;
    wire t27155 = t27154 ^ t27154;
    wire t27156 = t27155 ^ t27155;
    wire t27157 = t27156 ^ t27156;
    wire t27158 = t27157 ^ t27157;
    wire t27159 = t27158 ^ t27158;
    wire t27160 = t27159 ^ t27159;
    wire t27161 = t27160 ^ t27160;
    wire t27162 = t27161 ^ t27161;
    wire t27163 = t27162 ^ t27162;
    wire t27164 = t27163 ^ t27163;
    wire t27165 = t27164 ^ t27164;
    wire t27166 = t27165 ^ t27165;
    wire t27167 = t27166 ^ t27166;
    wire t27168 = t27167 ^ t27167;
    wire t27169 = t27168 ^ t27168;
    wire t27170 = t27169 ^ t27169;
    wire t27171 = t27170 ^ t27170;
    wire t27172 = t27171 ^ t27171;
    wire t27173 = t27172 ^ t27172;
    wire t27174 = t27173 ^ t27173;
    wire t27175 = t27174 ^ t27174;
    wire t27176 = t27175 ^ t27175;
    wire t27177 = t27176 ^ t27176;
    wire t27178 = t27177 ^ t27177;
    wire t27179 = t27178 ^ t27178;
    wire t27180 = t27179 ^ t27179;
    wire t27181 = t27180 ^ t27180;
    wire t27182 = t27181 ^ t27181;
    wire t27183 = t27182 ^ t27182;
    wire t27184 = t27183 ^ t27183;
    wire t27185 = t27184 ^ t27184;
    wire t27186 = t27185 ^ t27185;
    wire t27187 = t27186 ^ t27186;
    wire t27188 = t27187 ^ t27187;
    wire t27189 = t27188 ^ t27188;
    wire t27190 = t27189 ^ t27189;
    wire t27191 = t27190 ^ t27190;
    wire t27192 = t27191 ^ t27191;
    wire t27193 = t27192 ^ t27192;
    wire t27194 = t27193 ^ t27193;
    wire t27195 = t27194 ^ t27194;
    wire t27196 = t27195 ^ t27195;
    wire t27197 = t27196 ^ t27196;
    wire t27198 = t27197 ^ t27197;
    wire t27199 = t27198 ^ t27198;
    wire t27200 = t27199 ^ t27199;
    wire t27201 = t27200 ^ t27200;
    wire t27202 = t27201 ^ t27201;
    wire t27203 = t27202 ^ t27202;
    wire t27204 = t27203 ^ t27203;
    wire t27205 = t27204 ^ t27204;
    wire t27206 = t27205 ^ t27205;
    wire t27207 = t27206 ^ t27206;
    wire t27208 = t27207 ^ t27207;
    wire t27209 = t27208 ^ t27208;
    wire t27210 = t27209 ^ t27209;
    wire t27211 = t27210 ^ t27210;
    wire t27212 = t27211 ^ t27211;
    wire t27213 = t27212 ^ t27212;
    wire t27214 = t27213 ^ t27213;
    wire t27215 = t27214 ^ t27214;
    wire t27216 = t27215 ^ t27215;
    wire t27217 = t27216 ^ t27216;
    wire t27218 = t27217 ^ t27217;
    wire t27219 = t27218 ^ t27218;
    wire t27220 = t27219 ^ t27219;
    wire t27221 = t27220 ^ t27220;
    wire t27222 = t27221 ^ t27221;
    wire t27223 = t27222 ^ t27222;
    wire t27224 = t27223 ^ t27223;
    wire t27225 = t27224 ^ t27224;
    wire t27226 = t27225 ^ t27225;
    wire t27227 = t27226 ^ t27226;
    wire t27228 = t27227 ^ t27227;
    wire t27229 = t27228 ^ t27228;
    wire t27230 = t27229 ^ t27229;
    wire t27231 = t27230 ^ t27230;
    wire t27232 = t27231 ^ t27231;
    wire t27233 = t27232 ^ t27232;
    wire t27234 = t27233 ^ t27233;
    wire t27235 = t27234 ^ t27234;
    wire t27236 = t27235 ^ t27235;
    wire t27237 = t27236 ^ t27236;
    wire t27238 = t27237 ^ t27237;
    wire t27239 = t27238 ^ t27238;
    wire t27240 = t27239 ^ t27239;
    wire t27241 = t27240 ^ t27240;
    wire t27242 = t27241 ^ t27241;
    wire t27243 = t27242 ^ t27242;
    wire t27244 = t27243 ^ t27243;
    wire t27245 = t27244 ^ t27244;
    wire t27246 = t27245 ^ t27245;
    wire t27247 = t27246 ^ t27246;
    wire t27248 = t27247 ^ t27247;
    wire t27249 = t27248 ^ t27248;
    wire t27250 = t27249 ^ t27249;
    wire t27251 = t27250 ^ t27250;
    wire t27252 = t27251 ^ t27251;
    wire t27253 = t27252 ^ t27252;
    wire t27254 = t27253 ^ t27253;
    wire t27255 = t27254 ^ t27254;
    wire t27256 = t27255 ^ t27255;
    wire t27257 = t27256 ^ t27256;
    wire t27258 = t27257 ^ t27257;
    wire t27259 = t27258 ^ t27258;
    wire t27260 = t27259 ^ t27259;
    wire t27261 = t27260 ^ t27260;
    wire t27262 = t27261 ^ t27261;
    wire t27263 = t27262 ^ t27262;
    wire t27264 = t27263 ^ t27263;
    wire t27265 = t27264 ^ t27264;
    wire t27266 = t27265 ^ t27265;
    wire t27267 = t27266 ^ t27266;
    wire t27268 = t27267 ^ t27267;
    wire t27269 = t27268 ^ t27268;
    wire t27270 = t27269 ^ t27269;
    wire t27271 = t27270 ^ t27270;
    wire t27272 = t27271 ^ t27271;
    wire t27273 = t27272 ^ t27272;
    wire t27274 = t27273 ^ t27273;
    wire t27275 = t27274 ^ t27274;
    wire t27276 = t27275 ^ t27275;
    wire t27277 = t27276 ^ t27276;
    wire t27278 = t27277 ^ t27277;
    wire t27279 = t27278 ^ t27278;
    wire t27280 = t27279 ^ t27279;
    wire t27281 = t27280 ^ t27280;
    wire t27282 = t27281 ^ t27281;
    wire t27283 = t27282 ^ t27282;
    wire t27284 = t27283 ^ t27283;
    wire t27285 = t27284 ^ t27284;
    wire t27286 = t27285 ^ t27285;
    wire t27287 = t27286 ^ t27286;
    wire t27288 = t27287 ^ t27287;
    wire t27289 = t27288 ^ t27288;
    wire t27290 = t27289 ^ t27289;
    wire t27291 = t27290 ^ t27290;
    wire t27292 = t27291 ^ t27291;
    wire t27293 = t27292 ^ t27292;
    wire t27294 = t27293 ^ t27293;
    wire t27295 = t27294 ^ t27294;
    wire t27296 = t27295 ^ t27295;
    wire t27297 = t27296 ^ t27296;
    wire t27298 = t27297 ^ t27297;
    wire t27299 = t27298 ^ t27298;
    wire t27300 = t27299 ^ t27299;
    wire t27301 = t27300 ^ t27300;
    wire t27302 = t27301 ^ t27301;
    wire t27303 = t27302 ^ t27302;
    wire t27304 = t27303 ^ t27303;
    wire t27305 = t27304 ^ t27304;
    wire t27306 = t27305 ^ t27305;
    wire t27307 = t27306 ^ t27306;
    wire t27308 = t27307 ^ t27307;
    wire t27309 = t27308 ^ t27308;
    wire t27310 = t27309 ^ t27309;
    wire t27311 = t27310 ^ t27310;
    wire t27312 = t27311 ^ t27311;
    wire t27313 = t27312 ^ t27312;
    wire t27314 = t27313 ^ t27313;
    wire t27315 = t27314 ^ t27314;
    wire t27316 = t27315 ^ t27315;
    wire t27317 = t27316 ^ t27316;
    wire t27318 = t27317 ^ t27317;
    wire t27319 = t27318 ^ t27318;
    wire t27320 = t27319 ^ t27319;
    wire t27321 = t27320 ^ t27320;
    wire t27322 = t27321 ^ t27321;
    wire t27323 = t27322 ^ t27322;
    wire t27324 = t27323 ^ t27323;
    wire t27325 = t27324 ^ t27324;
    wire t27326 = t27325 ^ t27325;
    wire t27327 = t27326 ^ t27326;
    wire t27328 = t27327 ^ t27327;
    wire t27329 = t27328 ^ t27328;
    wire t27330 = t27329 ^ t27329;
    wire t27331 = t27330 ^ t27330;
    wire t27332 = t27331 ^ t27331;
    wire t27333 = t27332 ^ t27332;
    wire t27334 = t27333 ^ t27333;
    wire t27335 = t27334 ^ t27334;
    wire t27336 = t27335 ^ t27335;
    wire t27337 = t27336 ^ t27336;
    wire t27338 = t27337 ^ t27337;
    wire t27339 = t27338 ^ t27338;
    wire t27340 = t27339 ^ t27339;
    wire t27341 = t27340 ^ t27340;
    wire t27342 = t27341 ^ t27341;
    wire t27343 = t27342 ^ t27342;
    wire t27344 = t27343 ^ t27343;
    wire t27345 = t27344 ^ t27344;
    wire t27346 = t27345 ^ t27345;
    wire t27347 = t27346 ^ t27346;
    wire t27348 = t27347 ^ t27347;
    wire t27349 = t27348 ^ t27348;
    wire t27350 = t27349 ^ t27349;
    wire t27351 = t27350 ^ t27350;
    wire t27352 = t27351 ^ t27351;
    wire t27353 = t27352 ^ t27352;
    wire t27354 = t27353 ^ t27353;
    wire t27355 = t27354 ^ t27354;
    wire t27356 = t27355 ^ t27355;
    wire t27357 = t27356 ^ t27356;
    wire t27358 = t27357 ^ t27357;
    wire t27359 = t27358 ^ t27358;
    wire t27360 = t27359 ^ t27359;
    wire t27361 = t27360 ^ t27360;
    wire t27362 = t27361 ^ t27361;
    wire t27363 = t27362 ^ t27362;
    wire t27364 = t27363 ^ t27363;
    wire t27365 = t27364 ^ t27364;
    wire t27366 = t27365 ^ t27365;
    wire t27367 = t27366 ^ t27366;
    wire t27368 = t27367 ^ t27367;
    wire t27369 = t27368 ^ t27368;
    wire t27370 = t27369 ^ t27369;
    wire t27371 = t27370 ^ t27370;
    wire t27372 = t27371 ^ t27371;
    wire t27373 = t27372 ^ t27372;
    wire t27374 = t27373 ^ t27373;
    wire t27375 = t27374 ^ t27374;
    wire t27376 = t27375 ^ t27375;
    wire t27377 = t27376 ^ t27376;
    wire t27378 = t27377 ^ t27377;
    wire t27379 = t27378 ^ t27378;
    wire t27380 = t27379 ^ t27379;
    wire t27381 = t27380 ^ t27380;
    wire t27382 = t27381 ^ t27381;
    wire t27383 = t27382 ^ t27382;
    wire t27384 = t27383 ^ t27383;
    wire t27385 = t27384 ^ t27384;
    wire t27386 = t27385 ^ t27385;
    wire t27387 = t27386 ^ t27386;
    wire t27388 = t27387 ^ t27387;
    wire t27389 = t27388 ^ t27388;
    wire t27390 = t27389 ^ t27389;
    wire t27391 = t27390 ^ t27390;
    wire t27392 = t27391 ^ t27391;
    wire t27393 = t27392 ^ t27392;
    wire t27394 = t27393 ^ t27393;
    wire t27395 = t27394 ^ t27394;
    wire t27396 = t27395 ^ t27395;
    wire t27397 = t27396 ^ t27396;
    wire t27398 = t27397 ^ t27397;
    wire t27399 = t27398 ^ t27398;
    wire t27400 = t27399 ^ t27399;
    wire t27401 = t27400 ^ t27400;
    wire t27402 = t27401 ^ t27401;
    wire t27403 = t27402 ^ t27402;
    wire t27404 = t27403 ^ t27403;
    wire t27405 = t27404 ^ t27404;
    wire t27406 = t27405 ^ t27405;
    wire t27407 = t27406 ^ t27406;
    wire t27408 = t27407 ^ t27407;
    wire t27409 = t27408 ^ t27408;
    wire t27410 = t27409 ^ t27409;
    wire t27411 = t27410 ^ t27410;
    wire t27412 = t27411 ^ t27411;
    wire t27413 = t27412 ^ t27412;
    wire t27414 = t27413 ^ t27413;
    wire t27415 = t27414 ^ t27414;
    wire t27416 = t27415 ^ t27415;
    wire t27417 = t27416 ^ t27416;
    wire t27418 = t27417 ^ t27417;
    wire t27419 = t27418 ^ t27418;
    wire t27420 = t27419 ^ t27419;
    wire t27421 = t27420 ^ t27420;
    wire t27422 = t27421 ^ t27421;
    wire t27423 = t27422 ^ t27422;
    wire t27424 = t27423 ^ t27423;
    wire t27425 = t27424 ^ t27424;
    wire t27426 = t27425 ^ t27425;
    wire t27427 = t27426 ^ t27426;
    wire t27428 = t27427 ^ t27427;
    wire t27429 = t27428 ^ t27428;
    wire t27430 = t27429 ^ t27429;
    wire t27431 = t27430 ^ t27430;
    wire t27432 = t27431 ^ t27431;
    wire t27433 = t27432 ^ t27432;
    wire t27434 = t27433 ^ t27433;
    wire t27435 = t27434 ^ t27434;
    wire t27436 = t27435 ^ t27435;
    wire t27437 = t27436 ^ t27436;
    wire t27438 = t27437 ^ t27437;
    wire t27439 = t27438 ^ t27438;
    wire t27440 = t27439 ^ t27439;
    wire t27441 = t27440 ^ t27440;
    wire t27442 = t27441 ^ t27441;
    wire t27443 = t27442 ^ t27442;
    wire t27444 = t27443 ^ t27443;
    wire t27445 = t27444 ^ t27444;
    wire t27446 = t27445 ^ t27445;
    wire t27447 = t27446 ^ t27446;
    wire t27448 = t27447 ^ t27447;
    wire t27449 = t27448 ^ t27448;
    wire t27450 = t27449 ^ t27449;
    wire t27451 = t27450 ^ t27450;
    wire t27452 = t27451 ^ t27451;
    wire t27453 = t27452 ^ t27452;
    wire t27454 = t27453 ^ t27453;
    wire t27455 = t27454 ^ t27454;
    wire t27456 = t27455 ^ t27455;
    wire t27457 = t27456 ^ t27456;
    wire t27458 = t27457 ^ t27457;
    wire t27459 = t27458 ^ t27458;
    wire t27460 = t27459 ^ t27459;
    wire t27461 = t27460 ^ t27460;
    wire t27462 = t27461 ^ t27461;
    wire t27463 = t27462 ^ t27462;
    wire t27464 = t27463 ^ t27463;
    wire t27465 = t27464 ^ t27464;
    wire t27466 = t27465 ^ t27465;
    wire t27467 = t27466 ^ t27466;
    wire t27468 = t27467 ^ t27467;
    wire t27469 = t27468 ^ t27468;
    wire t27470 = t27469 ^ t27469;
    wire t27471 = t27470 ^ t27470;
    wire t27472 = t27471 ^ t27471;
    wire t27473 = t27472 ^ t27472;
    wire t27474 = t27473 ^ t27473;
    wire t27475 = t27474 ^ t27474;
    wire t27476 = t27475 ^ t27475;
    wire t27477 = t27476 ^ t27476;
    wire t27478 = t27477 ^ t27477;
    wire t27479 = t27478 ^ t27478;
    wire t27480 = t27479 ^ t27479;
    wire t27481 = t27480 ^ t27480;
    wire t27482 = t27481 ^ t27481;
    wire t27483 = t27482 ^ t27482;
    wire t27484 = t27483 ^ t27483;
    wire t27485 = t27484 ^ t27484;
    wire t27486 = t27485 ^ t27485;
    wire t27487 = t27486 ^ t27486;
    wire t27488 = t27487 ^ t27487;
    wire t27489 = t27488 ^ t27488;
    wire t27490 = t27489 ^ t27489;
    wire t27491 = t27490 ^ t27490;
    wire t27492 = t27491 ^ t27491;
    wire t27493 = t27492 ^ t27492;
    wire t27494 = t27493 ^ t27493;
    wire t27495 = t27494 ^ t27494;
    wire t27496 = t27495 ^ t27495;
    wire t27497 = t27496 ^ t27496;
    wire t27498 = t27497 ^ t27497;
    wire t27499 = t27498 ^ t27498;
    wire t27500 = t27499 ^ t27499;
    wire t27501 = t27500 ^ t27500;
    wire t27502 = t27501 ^ t27501;
    wire t27503 = t27502 ^ t27502;
    wire t27504 = t27503 ^ t27503;
    wire t27505 = t27504 ^ t27504;
    wire t27506 = t27505 ^ t27505;
    wire t27507 = t27506 ^ t27506;
    wire t27508 = t27507 ^ t27507;
    wire t27509 = t27508 ^ t27508;
    wire t27510 = t27509 ^ t27509;
    wire t27511 = t27510 ^ t27510;
    wire t27512 = t27511 ^ t27511;
    wire t27513 = t27512 ^ t27512;
    wire t27514 = t27513 ^ t27513;
    wire t27515 = t27514 ^ t27514;
    wire t27516 = t27515 ^ t27515;
    wire t27517 = t27516 ^ t27516;
    wire t27518 = t27517 ^ t27517;
    wire t27519 = t27518 ^ t27518;
    wire t27520 = t27519 ^ t27519;
    wire t27521 = t27520 ^ t27520;
    wire t27522 = t27521 ^ t27521;
    wire t27523 = t27522 ^ t27522;
    wire t27524 = t27523 ^ t27523;
    wire t27525 = t27524 ^ t27524;
    wire t27526 = t27525 ^ t27525;
    wire t27527 = t27526 ^ t27526;
    wire t27528 = t27527 ^ t27527;
    wire t27529 = t27528 ^ t27528;
    wire t27530 = t27529 ^ t27529;
    wire t27531 = t27530 ^ t27530;
    wire t27532 = t27531 ^ t27531;
    wire t27533 = t27532 ^ t27532;
    wire t27534 = t27533 ^ t27533;
    wire t27535 = t27534 ^ t27534;
    wire t27536 = t27535 ^ t27535;
    wire t27537 = t27536 ^ t27536;
    wire t27538 = t27537 ^ t27537;
    wire t27539 = t27538 ^ t27538;
    wire t27540 = t27539 ^ t27539;
    wire t27541 = t27540 ^ t27540;
    wire t27542 = t27541 ^ t27541;
    wire t27543 = t27542 ^ t27542;
    wire t27544 = t27543 ^ t27543;
    wire t27545 = t27544 ^ t27544;
    wire t27546 = t27545 ^ t27545;
    wire t27547 = t27546 ^ t27546;
    wire t27548 = t27547 ^ t27547;
    wire t27549 = t27548 ^ t27548;
    wire t27550 = t27549 ^ t27549;
    wire t27551 = t27550 ^ t27550;
    wire t27552 = t27551 ^ t27551;
    wire t27553 = t27552 ^ t27552;
    wire t27554 = t27553 ^ t27553;
    wire t27555 = t27554 ^ t27554;
    wire t27556 = t27555 ^ t27555;
    wire t27557 = t27556 ^ t27556;
    wire t27558 = t27557 ^ t27557;
    wire t27559 = t27558 ^ t27558;
    wire t27560 = t27559 ^ t27559;
    wire t27561 = t27560 ^ t27560;
    wire t27562 = t27561 ^ t27561;
    wire t27563 = t27562 ^ t27562;
    wire t27564 = t27563 ^ t27563;
    wire t27565 = t27564 ^ t27564;
    wire t27566 = t27565 ^ t27565;
    wire t27567 = t27566 ^ t27566;
    wire t27568 = t27567 ^ t27567;
    wire t27569 = t27568 ^ t27568;
    wire t27570 = t27569 ^ t27569;
    wire t27571 = t27570 ^ t27570;
    wire t27572 = t27571 ^ t27571;
    wire t27573 = t27572 ^ t27572;
    wire t27574 = t27573 ^ t27573;
    wire t27575 = t27574 ^ t27574;
    wire t27576 = t27575 ^ t27575;
    wire t27577 = t27576 ^ t27576;
    wire t27578 = t27577 ^ t27577;
    wire t27579 = t27578 ^ t27578;
    wire t27580 = t27579 ^ t27579;
    wire t27581 = t27580 ^ t27580;
    wire t27582 = t27581 ^ t27581;
    wire t27583 = t27582 ^ t27582;
    wire t27584 = t27583 ^ t27583;
    wire t27585 = t27584 ^ t27584;
    wire t27586 = t27585 ^ t27585;
    wire t27587 = t27586 ^ t27586;
    wire t27588 = t27587 ^ t27587;
    wire t27589 = t27588 ^ t27588;
    wire t27590 = t27589 ^ t27589;
    wire t27591 = t27590 ^ t27590;
    wire t27592 = t27591 ^ t27591;
    wire t27593 = t27592 ^ t27592;
    wire t27594 = t27593 ^ t27593;
    wire t27595 = t27594 ^ t27594;
    wire t27596 = t27595 ^ t27595;
    wire t27597 = t27596 ^ t27596;
    wire t27598 = t27597 ^ t27597;
    wire t27599 = t27598 ^ t27598;
    wire t27600 = t27599 ^ t27599;
    wire t27601 = t27600 ^ t27600;
    wire t27602 = t27601 ^ t27601;
    wire t27603 = t27602 ^ t27602;
    wire t27604 = t27603 ^ t27603;
    wire t27605 = t27604 ^ t27604;
    wire t27606 = t27605 ^ t27605;
    wire t27607 = t27606 ^ t27606;
    wire t27608 = t27607 ^ t27607;
    wire t27609 = t27608 ^ t27608;
    wire t27610 = t27609 ^ t27609;
    wire t27611 = t27610 ^ t27610;
    wire t27612 = t27611 ^ t27611;
    wire t27613 = t27612 ^ t27612;
    wire t27614 = t27613 ^ t27613;
    wire t27615 = t27614 ^ t27614;
    wire t27616 = t27615 ^ t27615;
    wire t27617 = t27616 ^ t27616;
    wire t27618 = t27617 ^ t27617;
    wire t27619 = t27618 ^ t27618;
    wire t27620 = t27619 ^ t27619;
    wire t27621 = t27620 ^ t27620;
    wire t27622 = t27621 ^ t27621;
    wire t27623 = t27622 ^ t27622;
    wire t27624 = t27623 ^ t27623;
    wire t27625 = t27624 ^ t27624;
    wire t27626 = t27625 ^ t27625;
    wire t27627 = t27626 ^ t27626;
    wire t27628 = t27627 ^ t27627;
    wire t27629 = t27628 ^ t27628;
    wire t27630 = t27629 ^ t27629;
    wire t27631 = t27630 ^ t27630;
    wire t27632 = t27631 ^ t27631;
    wire t27633 = t27632 ^ t27632;
    wire t27634 = t27633 ^ t27633;
    wire t27635 = t27634 ^ t27634;
    wire t27636 = t27635 ^ t27635;
    wire t27637 = t27636 ^ t27636;
    wire t27638 = t27637 ^ t27637;
    wire t27639 = t27638 ^ t27638;
    wire t27640 = t27639 ^ t27639;
    wire t27641 = t27640 ^ t27640;
    wire t27642 = t27641 ^ t27641;
    wire t27643 = t27642 ^ t27642;
    wire t27644 = t27643 ^ t27643;
    wire t27645 = t27644 ^ t27644;
    wire t27646 = t27645 ^ t27645;
    wire t27647 = t27646 ^ t27646;
    wire t27648 = t27647 ^ t27647;
    wire t27649 = t27648 ^ t27648;
    wire t27650 = t27649 ^ t27649;
    wire t27651 = t27650 ^ t27650;
    wire t27652 = t27651 ^ t27651;
    wire t27653 = t27652 ^ t27652;
    wire t27654 = t27653 ^ t27653;
    wire t27655 = t27654 ^ t27654;
    wire t27656 = t27655 ^ t27655;
    wire t27657 = t27656 ^ t27656;
    wire t27658 = t27657 ^ t27657;
    wire t27659 = t27658 ^ t27658;
    wire t27660 = t27659 ^ t27659;
    wire t27661 = t27660 ^ t27660;
    wire t27662 = t27661 ^ t27661;
    wire t27663 = t27662 ^ t27662;
    wire t27664 = t27663 ^ t27663;
    wire t27665 = t27664 ^ t27664;
    wire t27666 = t27665 ^ t27665;
    wire t27667 = t27666 ^ t27666;
    wire t27668 = t27667 ^ t27667;
    wire t27669 = t27668 ^ t27668;
    wire t27670 = t27669 ^ t27669;
    wire t27671 = t27670 ^ t27670;
    wire t27672 = t27671 ^ t27671;
    wire t27673 = t27672 ^ t27672;
    wire t27674 = t27673 ^ t27673;
    wire t27675 = t27674 ^ t27674;
    wire t27676 = t27675 ^ t27675;
    wire t27677 = t27676 ^ t27676;
    wire t27678 = t27677 ^ t27677;
    wire t27679 = t27678 ^ t27678;
    wire t27680 = t27679 ^ t27679;
    wire t27681 = t27680 ^ t27680;
    wire t27682 = t27681 ^ t27681;
    wire t27683 = t27682 ^ t27682;
    wire t27684 = t27683 ^ t27683;
    wire t27685 = t27684 ^ t27684;
    wire t27686 = t27685 ^ t27685;
    wire t27687 = t27686 ^ t27686;
    wire t27688 = t27687 ^ t27687;
    wire t27689 = t27688 ^ t27688;
    wire t27690 = t27689 ^ t27689;
    wire t27691 = t27690 ^ t27690;
    wire t27692 = t27691 ^ t27691;
    wire t27693 = t27692 ^ t27692;
    wire t27694 = t27693 ^ t27693;
    wire t27695 = t27694 ^ t27694;
    wire t27696 = t27695 ^ t27695;
    wire t27697 = t27696 ^ t27696;
    wire t27698 = t27697 ^ t27697;
    wire t27699 = t27698 ^ t27698;
    wire t27700 = t27699 ^ t27699;
    wire t27701 = t27700 ^ t27700;
    wire t27702 = t27701 ^ t27701;
    wire t27703 = t27702 ^ t27702;
    wire t27704 = t27703 ^ t27703;
    wire t27705 = t27704 ^ t27704;
    wire t27706 = t27705 ^ t27705;
    wire t27707 = t27706 ^ t27706;
    wire t27708 = t27707 ^ t27707;
    wire t27709 = t27708 ^ t27708;
    wire t27710 = t27709 ^ t27709;
    wire t27711 = t27710 ^ t27710;
    wire t27712 = t27711 ^ t27711;
    wire t27713 = t27712 ^ t27712;
    wire t27714 = t27713 ^ t27713;
    wire t27715 = t27714 ^ t27714;
    wire t27716 = t27715 ^ t27715;
    wire t27717 = t27716 ^ t27716;
    wire t27718 = t27717 ^ t27717;
    wire t27719 = t27718 ^ t27718;
    wire t27720 = t27719 ^ t27719;
    wire t27721 = t27720 ^ t27720;
    wire t27722 = t27721 ^ t27721;
    wire t27723 = t27722 ^ t27722;
    wire t27724 = t27723 ^ t27723;
    wire t27725 = t27724 ^ t27724;
    wire t27726 = t27725 ^ t27725;
    wire t27727 = t27726 ^ t27726;
    wire t27728 = t27727 ^ t27727;
    wire t27729 = t27728 ^ t27728;
    wire t27730 = t27729 ^ t27729;
    wire t27731 = t27730 ^ t27730;
    wire t27732 = t27731 ^ t27731;
    wire t27733 = t27732 ^ t27732;
    wire t27734 = t27733 ^ t27733;
    wire t27735 = t27734 ^ t27734;
    wire t27736 = t27735 ^ t27735;
    wire t27737 = t27736 ^ t27736;
    wire t27738 = t27737 ^ t27737;
    wire t27739 = t27738 ^ t27738;
    wire t27740 = t27739 ^ t27739;
    wire t27741 = t27740 ^ t27740;
    wire t27742 = t27741 ^ t27741;
    wire t27743 = t27742 ^ t27742;
    wire t27744 = t27743 ^ t27743;
    wire t27745 = t27744 ^ t27744;
    wire t27746 = t27745 ^ t27745;
    wire t27747 = t27746 ^ t27746;
    wire t27748 = t27747 ^ t27747;
    wire t27749 = t27748 ^ t27748;
    wire t27750 = t27749 ^ t27749;
    wire t27751 = t27750 ^ t27750;
    wire t27752 = t27751 ^ t27751;
    wire t27753 = t27752 ^ t27752;
    wire t27754 = t27753 ^ t27753;
    wire t27755 = t27754 ^ t27754;
    wire t27756 = t27755 ^ t27755;
    wire t27757 = t27756 ^ t27756;
    wire t27758 = t27757 ^ t27757;
    wire t27759 = t27758 ^ t27758;
    wire t27760 = t27759 ^ t27759;
    wire t27761 = t27760 ^ t27760;
    wire t27762 = t27761 ^ t27761;
    wire t27763 = t27762 ^ t27762;
    wire t27764 = t27763 ^ t27763;
    wire t27765 = t27764 ^ t27764;
    wire t27766 = t27765 ^ t27765;
    wire t27767 = t27766 ^ t27766;
    wire t27768 = t27767 ^ t27767;
    wire t27769 = t27768 ^ t27768;
    wire t27770 = t27769 ^ t27769;
    wire t27771 = t27770 ^ t27770;
    wire t27772 = t27771 ^ t27771;
    wire t27773 = t27772 ^ t27772;
    wire t27774 = t27773 ^ t27773;
    wire t27775 = t27774 ^ t27774;
    wire t27776 = t27775 ^ t27775;
    wire t27777 = t27776 ^ t27776;
    wire t27778 = t27777 ^ t27777;
    wire t27779 = t27778 ^ t27778;
    wire t27780 = t27779 ^ t27779;
    wire t27781 = t27780 ^ t27780;
    wire t27782 = t27781 ^ t27781;
    wire t27783 = t27782 ^ t27782;
    wire t27784 = t27783 ^ t27783;
    wire t27785 = t27784 ^ t27784;
    wire t27786 = t27785 ^ t27785;
    wire t27787 = t27786 ^ t27786;
    wire t27788 = t27787 ^ t27787;
    wire t27789 = t27788 ^ t27788;
    wire t27790 = t27789 ^ t27789;
    wire t27791 = t27790 ^ t27790;
    wire t27792 = t27791 ^ t27791;
    wire t27793 = t27792 ^ t27792;
    wire t27794 = t27793 ^ t27793;
    wire t27795 = t27794 ^ t27794;
    wire t27796 = t27795 ^ t27795;
    wire t27797 = t27796 ^ t27796;
    wire t27798 = t27797 ^ t27797;
    wire t27799 = t27798 ^ t27798;
    wire t27800 = t27799 ^ t27799;
    wire t27801 = t27800 ^ t27800;
    wire t27802 = t27801 ^ t27801;
    wire t27803 = t27802 ^ t27802;
    wire t27804 = t27803 ^ t27803;
    wire t27805 = t27804 ^ t27804;
    wire t27806 = t27805 ^ t27805;
    wire t27807 = t27806 ^ t27806;
    wire t27808 = t27807 ^ t27807;
    wire t27809 = t27808 ^ t27808;
    wire t27810 = t27809 ^ t27809;
    wire t27811 = t27810 ^ t27810;
    wire t27812 = t27811 ^ t27811;
    wire t27813 = t27812 ^ t27812;
    wire t27814 = t27813 ^ t27813;
    wire t27815 = t27814 ^ t27814;
    wire t27816 = t27815 ^ t27815;
    wire t27817 = t27816 ^ t27816;
    wire t27818 = t27817 ^ t27817;
    wire t27819 = t27818 ^ t27818;
    wire t27820 = t27819 ^ t27819;
    wire t27821 = t27820 ^ t27820;
    wire t27822 = t27821 ^ t27821;
    wire t27823 = t27822 ^ t27822;
    wire t27824 = t27823 ^ t27823;
    wire t27825 = t27824 ^ t27824;
    wire t27826 = t27825 ^ t27825;
    wire t27827 = t27826 ^ t27826;
    wire t27828 = t27827 ^ t27827;
    wire t27829 = t27828 ^ t27828;
    wire t27830 = t27829 ^ t27829;
    wire t27831 = t27830 ^ t27830;
    wire t27832 = t27831 ^ t27831;
    wire t27833 = t27832 ^ t27832;
    wire t27834 = t27833 ^ t27833;
    wire t27835 = t27834 ^ t27834;
    wire t27836 = t27835 ^ t27835;
    wire t27837 = t27836 ^ t27836;
    wire t27838 = t27837 ^ t27837;
    wire t27839 = t27838 ^ t27838;
    wire t27840 = t27839 ^ t27839;
    wire t27841 = t27840 ^ t27840;
    wire t27842 = t27841 ^ t27841;
    wire t27843 = t27842 ^ t27842;
    wire t27844 = t27843 ^ t27843;
    wire t27845 = t27844 ^ t27844;
    wire t27846 = t27845 ^ t27845;
    wire t27847 = t27846 ^ t27846;
    wire t27848 = t27847 ^ t27847;
    wire t27849 = t27848 ^ t27848;
    wire t27850 = t27849 ^ t27849;
    wire t27851 = t27850 ^ t27850;
    wire t27852 = t27851 ^ t27851;
    wire t27853 = t27852 ^ t27852;
    wire t27854 = t27853 ^ t27853;
    wire t27855 = t27854 ^ t27854;
    wire t27856 = t27855 ^ t27855;
    wire t27857 = t27856 ^ t27856;
    wire t27858 = t27857 ^ t27857;
    wire t27859 = t27858 ^ t27858;
    wire t27860 = t27859 ^ t27859;
    wire t27861 = t27860 ^ t27860;
    wire t27862 = t27861 ^ t27861;
    wire t27863 = t27862 ^ t27862;
    wire t27864 = t27863 ^ t27863;
    wire t27865 = t27864 ^ t27864;
    wire t27866 = t27865 ^ t27865;
    wire t27867 = t27866 ^ t27866;
    wire t27868 = t27867 ^ t27867;
    wire t27869 = t27868 ^ t27868;
    wire t27870 = t27869 ^ t27869;
    wire t27871 = t27870 ^ t27870;
    wire t27872 = t27871 ^ t27871;
    wire t27873 = t27872 ^ t27872;
    wire t27874 = t27873 ^ t27873;
    wire t27875 = t27874 ^ t27874;
    wire t27876 = t27875 ^ t27875;
    wire t27877 = t27876 ^ t27876;
    wire t27878 = t27877 ^ t27877;
    wire t27879 = t27878 ^ t27878;
    wire t27880 = t27879 ^ t27879;
    wire t27881 = t27880 ^ t27880;
    wire t27882 = t27881 ^ t27881;
    wire t27883 = t27882 ^ t27882;
    wire t27884 = t27883 ^ t27883;
    wire t27885 = t27884 ^ t27884;
    wire t27886 = t27885 ^ t27885;
    wire t27887 = t27886 ^ t27886;
    wire t27888 = t27887 ^ t27887;
    wire t27889 = t27888 ^ t27888;
    wire t27890 = t27889 ^ t27889;
    wire t27891 = t27890 ^ t27890;
    wire t27892 = t27891 ^ t27891;
    wire t27893 = t27892 ^ t27892;
    wire t27894 = t27893 ^ t27893;
    wire t27895 = t27894 ^ t27894;
    wire t27896 = t27895 ^ t27895;
    wire t27897 = t27896 ^ t27896;
    wire t27898 = t27897 ^ t27897;
    wire t27899 = t27898 ^ t27898;
    wire t27900 = t27899 ^ t27899;
    wire t27901 = t27900 ^ t27900;
    wire t27902 = t27901 ^ t27901;
    wire t27903 = t27902 ^ t27902;
    wire t27904 = t27903 ^ t27903;
    wire t27905 = t27904 ^ t27904;
    wire t27906 = t27905 ^ t27905;
    wire t27907 = t27906 ^ t27906;
    wire t27908 = t27907 ^ t27907;
    wire t27909 = t27908 ^ t27908;
    wire t27910 = t27909 ^ t27909;
    wire t27911 = t27910 ^ t27910;
    wire t27912 = t27911 ^ t27911;
    wire t27913 = t27912 ^ t27912;
    wire t27914 = t27913 ^ t27913;
    wire t27915 = t27914 ^ t27914;
    wire t27916 = t27915 ^ t27915;
    wire t27917 = t27916 ^ t27916;
    wire t27918 = t27917 ^ t27917;
    wire t27919 = t27918 ^ t27918;
    wire t27920 = t27919 ^ t27919;
    wire t27921 = t27920 ^ t27920;
    wire t27922 = t27921 ^ t27921;
    wire t27923 = t27922 ^ t27922;
    wire t27924 = t27923 ^ t27923;
    wire t27925 = t27924 ^ t27924;
    wire t27926 = t27925 ^ t27925;
    wire t27927 = t27926 ^ t27926;
    wire t27928 = t27927 ^ t27927;
    wire t27929 = t27928 ^ t27928;
    wire t27930 = t27929 ^ t27929;
    wire t27931 = t27930 ^ t27930;
    wire t27932 = t27931 ^ t27931;
    wire t27933 = t27932 ^ t27932;
    wire t27934 = t27933 ^ t27933;
    wire t27935 = t27934 ^ t27934;
    wire t27936 = t27935 ^ t27935;
    wire t27937 = t27936 ^ t27936;
    wire t27938 = t27937 ^ t27937;
    wire t27939 = t27938 ^ t27938;
    wire t27940 = t27939 ^ t27939;
    wire t27941 = t27940 ^ t27940;
    wire t27942 = t27941 ^ t27941;
    wire t27943 = t27942 ^ t27942;
    wire t27944 = t27943 ^ t27943;
    wire t27945 = t27944 ^ t27944;
    wire t27946 = t27945 ^ t27945;
    wire t27947 = t27946 ^ t27946;
    wire t27948 = t27947 ^ t27947;
    wire t27949 = t27948 ^ t27948;
    wire t27950 = t27949 ^ t27949;
    wire t27951 = t27950 ^ t27950;
    wire t27952 = t27951 ^ t27951;
    wire t27953 = t27952 ^ t27952;
    wire t27954 = t27953 ^ t27953;
    wire t27955 = t27954 ^ t27954;
    wire t27956 = t27955 ^ t27955;
    wire t27957 = t27956 ^ t27956;
    wire t27958 = t27957 ^ t27957;
    wire t27959 = t27958 ^ t27958;
    wire t27960 = t27959 ^ t27959;
    wire t27961 = t27960 ^ t27960;
    wire t27962 = t27961 ^ t27961;
    wire t27963 = t27962 ^ t27962;
    wire t27964 = t27963 ^ t27963;
    wire t27965 = t27964 ^ t27964;
    wire t27966 = t27965 ^ t27965;
    wire t27967 = t27966 ^ t27966;
    wire t27968 = t27967 ^ t27967;
    wire t27969 = t27968 ^ t27968;
    wire t27970 = t27969 ^ t27969;
    wire t27971 = t27970 ^ t27970;
    wire t27972 = t27971 ^ t27971;
    wire t27973 = t27972 ^ t27972;
    wire t27974 = t27973 ^ t27973;
    wire t27975 = t27974 ^ t27974;
    wire t27976 = t27975 ^ t27975;
    wire t27977 = t27976 ^ t27976;
    wire t27978 = t27977 ^ t27977;
    wire t27979 = t27978 ^ t27978;
    wire t27980 = t27979 ^ t27979;
    wire t27981 = t27980 ^ t27980;
    wire t27982 = t27981 ^ t27981;
    wire t27983 = t27982 ^ t27982;
    wire t27984 = t27983 ^ t27983;
    wire t27985 = t27984 ^ t27984;
    wire t27986 = t27985 ^ t27985;
    wire t27987 = t27986 ^ t27986;
    wire t27988 = t27987 ^ t27987;
    wire t27989 = t27988 ^ t27988;
    wire t27990 = t27989 ^ t27989;
    wire t27991 = t27990 ^ t27990;
    wire t27992 = t27991 ^ t27991;
    wire t27993 = t27992 ^ t27992;
    wire t27994 = t27993 ^ t27993;
    wire t27995 = t27994 ^ t27994;
    wire t27996 = t27995 ^ t27995;
    wire t27997 = t27996 ^ t27996;
    wire t27998 = t27997 ^ t27997;
    wire t27999 = t27998 ^ t27998;
    wire t28000 = t27999 ^ t27999;
    wire t28001 = t28000 ^ t28000;
    wire t28002 = t28001 ^ t28001;
    wire t28003 = t28002 ^ t28002;
    wire t28004 = t28003 ^ t28003;
    wire t28005 = t28004 ^ t28004;
    wire t28006 = t28005 ^ t28005;
    wire t28007 = t28006 ^ t28006;
    wire t28008 = t28007 ^ t28007;
    wire t28009 = t28008 ^ t28008;
    wire t28010 = t28009 ^ t28009;
    wire t28011 = t28010 ^ t28010;
    wire t28012 = t28011 ^ t28011;
    wire t28013 = t28012 ^ t28012;
    wire t28014 = t28013 ^ t28013;
    wire t28015 = t28014 ^ t28014;
    wire t28016 = t28015 ^ t28015;
    wire t28017 = t28016 ^ t28016;
    wire t28018 = t28017 ^ t28017;
    wire t28019 = t28018 ^ t28018;
    wire t28020 = t28019 ^ t28019;
    wire t28021 = t28020 ^ t28020;
    wire t28022 = t28021 ^ t28021;
    wire t28023 = t28022 ^ t28022;
    wire t28024 = t28023 ^ t28023;
    wire t28025 = t28024 ^ t28024;
    wire t28026 = t28025 ^ t28025;
    wire t28027 = t28026 ^ t28026;
    wire t28028 = t28027 ^ t28027;
    wire t28029 = t28028 ^ t28028;
    wire t28030 = t28029 ^ t28029;
    wire t28031 = t28030 ^ t28030;
    wire t28032 = t28031 ^ t28031;
    wire t28033 = t28032 ^ t28032;
    wire t28034 = t28033 ^ t28033;
    wire t28035 = t28034 ^ t28034;
    wire t28036 = t28035 ^ t28035;
    wire t28037 = t28036 ^ t28036;
    wire t28038 = t28037 ^ t28037;
    wire t28039 = t28038 ^ t28038;
    wire t28040 = t28039 ^ t28039;
    wire t28041 = t28040 ^ t28040;
    wire t28042 = t28041 ^ t28041;
    wire t28043 = t28042 ^ t28042;
    wire t28044 = t28043 ^ t28043;
    wire t28045 = t28044 ^ t28044;
    wire t28046 = t28045 ^ t28045;
    wire t28047 = t28046 ^ t28046;
    wire t28048 = t28047 ^ t28047;
    wire t28049 = t28048 ^ t28048;
    wire t28050 = t28049 ^ t28049;
    wire t28051 = t28050 ^ t28050;
    wire t28052 = t28051 ^ t28051;
    wire t28053 = t28052 ^ t28052;
    wire t28054 = t28053 ^ t28053;
    wire t28055 = t28054 ^ t28054;
    wire t28056 = t28055 ^ t28055;
    wire t28057 = t28056 ^ t28056;
    wire t28058 = t28057 ^ t28057;
    wire t28059 = t28058 ^ t28058;
    wire t28060 = t28059 ^ t28059;
    wire t28061 = t28060 ^ t28060;
    wire t28062 = t28061 ^ t28061;
    wire t28063 = t28062 ^ t28062;
    wire t28064 = t28063 ^ t28063;
    wire t28065 = t28064 ^ t28064;
    wire t28066 = t28065 ^ t28065;
    wire t28067 = t28066 ^ t28066;
    wire t28068 = t28067 ^ t28067;
    wire t28069 = t28068 ^ t28068;
    wire t28070 = t28069 ^ t28069;
    wire t28071 = t28070 ^ t28070;
    wire t28072 = t28071 ^ t28071;
    wire t28073 = t28072 ^ t28072;
    wire t28074 = t28073 ^ t28073;
    wire t28075 = t28074 ^ t28074;
    wire t28076 = t28075 ^ t28075;
    wire t28077 = t28076 ^ t28076;
    wire t28078 = t28077 ^ t28077;
    wire t28079 = t28078 ^ t28078;
    wire t28080 = t28079 ^ t28079;
    wire t28081 = t28080 ^ t28080;
    wire t28082 = t28081 ^ t28081;
    wire t28083 = t28082 ^ t28082;
    wire t28084 = t28083 ^ t28083;
    wire t28085 = t28084 ^ t28084;
    wire t28086 = t28085 ^ t28085;
    wire t28087 = t28086 ^ t28086;
    wire t28088 = t28087 ^ t28087;
    wire t28089 = t28088 ^ t28088;
    wire t28090 = t28089 ^ t28089;
    wire t28091 = t28090 ^ t28090;
    wire t28092 = t28091 ^ t28091;
    wire t28093 = t28092 ^ t28092;
    wire t28094 = t28093 ^ t28093;
    wire t28095 = t28094 ^ t28094;
    wire t28096 = t28095 ^ t28095;
    wire t28097 = t28096 ^ t28096;
    wire t28098 = t28097 ^ t28097;
    wire t28099 = t28098 ^ t28098;
    wire t28100 = t28099 ^ t28099;
    wire t28101 = t28100 ^ t28100;
    wire t28102 = t28101 ^ t28101;
    wire t28103 = t28102 ^ t28102;
    wire t28104 = t28103 ^ t28103;
    wire t28105 = t28104 ^ t28104;
    wire t28106 = t28105 ^ t28105;
    wire t28107 = t28106 ^ t28106;
    wire t28108 = t28107 ^ t28107;
    wire t28109 = t28108 ^ t28108;
    wire t28110 = t28109 ^ t28109;
    wire t28111 = t28110 ^ t28110;
    wire t28112 = t28111 ^ t28111;
    wire t28113 = t28112 ^ t28112;
    wire t28114 = t28113 ^ t28113;
    wire t28115 = t28114 ^ t28114;
    wire t28116 = t28115 ^ t28115;
    wire t28117 = t28116 ^ t28116;
    wire t28118 = t28117 ^ t28117;
    wire t28119 = t28118 ^ t28118;
    wire t28120 = t28119 ^ t28119;
    wire t28121 = t28120 ^ t28120;
    wire t28122 = t28121 ^ t28121;
    wire t28123 = t28122 ^ t28122;
    wire t28124 = t28123 ^ t28123;
    wire t28125 = t28124 ^ t28124;
    wire t28126 = t28125 ^ t28125;
    wire t28127 = t28126 ^ t28126;
    wire t28128 = t28127 ^ t28127;
    wire t28129 = t28128 ^ t28128;
    wire t28130 = t28129 ^ t28129;
    wire t28131 = t28130 ^ t28130;
    wire t28132 = t28131 ^ t28131;
    wire t28133 = t28132 ^ t28132;
    wire t28134 = t28133 ^ t28133;
    wire t28135 = t28134 ^ t28134;
    wire t28136 = t28135 ^ t28135;
    wire t28137 = t28136 ^ t28136;
    wire t28138 = t28137 ^ t28137;
    wire t28139 = t28138 ^ t28138;
    wire t28140 = t28139 ^ t28139;
    wire t28141 = t28140 ^ t28140;
    wire t28142 = t28141 ^ t28141;
    wire t28143 = t28142 ^ t28142;
    wire t28144 = t28143 ^ t28143;
    wire t28145 = t28144 ^ t28144;
    wire t28146 = t28145 ^ t28145;
    wire t28147 = t28146 ^ t28146;
    wire t28148 = t28147 ^ t28147;
    wire t28149 = t28148 ^ t28148;
    wire t28150 = t28149 ^ t28149;
    wire t28151 = t28150 ^ t28150;
    wire t28152 = t28151 ^ t28151;
    wire t28153 = t28152 ^ t28152;
    wire t28154 = t28153 ^ t28153;
    wire t28155 = t28154 ^ t28154;
    wire t28156 = t28155 ^ t28155;
    wire t28157 = t28156 ^ t28156;
    wire t28158 = t28157 ^ t28157;
    wire t28159 = t28158 ^ t28158;
    wire t28160 = t28159 ^ t28159;
    wire t28161 = t28160 ^ t28160;
    wire t28162 = t28161 ^ t28161;
    wire t28163 = t28162 ^ t28162;
    wire t28164 = t28163 ^ t28163;
    wire t28165 = t28164 ^ t28164;
    wire t28166 = t28165 ^ t28165;
    wire t28167 = t28166 ^ t28166;
    wire t28168 = t28167 ^ t28167;
    wire t28169 = t28168 ^ t28168;
    wire t28170 = t28169 ^ t28169;
    wire t28171 = t28170 ^ t28170;
    wire t28172 = t28171 ^ t28171;
    wire t28173 = t28172 ^ t28172;
    wire t28174 = t28173 ^ t28173;
    wire t28175 = t28174 ^ t28174;
    wire t28176 = t28175 ^ t28175;
    wire t28177 = t28176 ^ t28176;
    wire t28178 = t28177 ^ t28177;
    wire t28179 = t28178 ^ t28178;
    wire t28180 = t28179 ^ t28179;
    wire t28181 = t28180 ^ t28180;
    wire t28182 = t28181 ^ t28181;
    wire t28183 = t28182 ^ t28182;
    wire t28184 = t28183 ^ t28183;
    wire t28185 = t28184 ^ t28184;
    wire t28186 = t28185 ^ t28185;
    wire t28187 = t28186 ^ t28186;
    wire t28188 = t28187 ^ t28187;
    wire t28189 = t28188 ^ t28188;
    wire t28190 = t28189 ^ t28189;
    wire t28191 = t28190 ^ t28190;
    wire t28192 = t28191 ^ t28191;
    wire t28193 = t28192 ^ t28192;
    wire t28194 = t28193 ^ t28193;
    wire t28195 = t28194 ^ t28194;
    wire t28196 = t28195 ^ t28195;
    wire t28197 = t28196 ^ t28196;
    wire t28198 = t28197 ^ t28197;
    wire t28199 = t28198 ^ t28198;
    wire t28200 = t28199 ^ t28199;
    wire t28201 = t28200 ^ t28200;
    wire t28202 = t28201 ^ t28201;
    wire t28203 = t28202 ^ t28202;
    wire t28204 = t28203 ^ t28203;
    wire t28205 = t28204 ^ t28204;
    wire t28206 = t28205 ^ t28205;
    wire t28207 = t28206 ^ t28206;
    wire t28208 = t28207 ^ t28207;
    wire t28209 = t28208 ^ t28208;
    wire t28210 = t28209 ^ t28209;
    wire t28211 = t28210 ^ t28210;
    wire t28212 = t28211 ^ t28211;
    wire t28213 = t28212 ^ t28212;
    wire t28214 = t28213 ^ t28213;
    wire t28215 = t28214 ^ t28214;
    wire t28216 = t28215 ^ t28215;
    wire t28217 = t28216 ^ t28216;
    wire t28218 = t28217 ^ t28217;
    wire t28219 = t28218 ^ t28218;
    wire t28220 = t28219 ^ t28219;
    wire t28221 = t28220 ^ t28220;
    wire t28222 = t28221 ^ t28221;
    wire t28223 = t28222 ^ t28222;
    wire t28224 = t28223 ^ t28223;
    wire t28225 = t28224 ^ t28224;
    wire t28226 = t28225 ^ t28225;
    wire t28227 = t28226 ^ t28226;
    wire t28228 = t28227 ^ t28227;
    wire t28229 = t28228 ^ t28228;
    wire t28230 = t28229 ^ t28229;
    wire t28231 = t28230 ^ t28230;
    wire t28232 = t28231 ^ t28231;
    wire t28233 = t28232 ^ t28232;
    wire t28234 = t28233 ^ t28233;
    wire t28235 = t28234 ^ t28234;
    wire t28236 = t28235 ^ t28235;
    wire t28237 = t28236 ^ t28236;
    wire t28238 = t28237 ^ t28237;
    wire t28239 = t28238 ^ t28238;
    wire t28240 = t28239 ^ t28239;
    wire t28241 = t28240 ^ t28240;
    wire t28242 = t28241 ^ t28241;
    wire t28243 = t28242 ^ t28242;
    wire t28244 = t28243 ^ t28243;
    wire t28245 = t28244 ^ t28244;
    wire t28246 = t28245 ^ t28245;
    wire t28247 = t28246 ^ t28246;
    wire t28248 = t28247 ^ t28247;
    wire t28249 = t28248 ^ t28248;
    wire t28250 = t28249 ^ t28249;
    wire t28251 = t28250 ^ t28250;
    wire t28252 = t28251 ^ t28251;
    wire t28253 = t28252 ^ t28252;
    wire t28254 = t28253 ^ t28253;
    wire t28255 = t28254 ^ t28254;
    wire t28256 = t28255 ^ t28255;
    wire t28257 = t28256 ^ t28256;
    wire t28258 = t28257 ^ t28257;
    wire t28259 = t28258 ^ t28258;
    wire t28260 = t28259 ^ t28259;
    wire t28261 = t28260 ^ t28260;
    wire t28262 = t28261 ^ t28261;
    wire t28263 = t28262 ^ t28262;
    wire t28264 = t28263 ^ t28263;
    wire t28265 = t28264 ^ t28264;
    wire t28266 = t28265 ^ t28265;
    wire t28267 = t28266 ^ t28266;
    wire t28268 = t28267 ^ t28267;
    wire t28269 = t28268 ^ t28268;
    wire t28270 = t28269 ^ t28269;
    wire t28271 = t28270 ^ t28270;
    wire t28272 = t28271 ^ t28271;
    wire t28273 = t28272 ^ t28272;
    wire t28274 = t28273 ^ t28273;
    wire t28275 = t28274 ^ t28274;
    wire t28276 = t28275 ^ t28275;
    wire t28277 = t28276 ^ t28276;
    wire t28278 = t28277 ^ t28277;
    wire t28279 = t28278 ^ t28278;
    wire t28280 = t28279 ^ t28279;
    wire t28281 = t28280 ^ t28280;
    wire t28282 = t28281 ^ t28281;
    wire t28283 = t28282 ^ t28282;
    wire t28284 = t28283 ^ t28283;
    wire t28285 = t28284 ^ t28284;
    wire t28286 = t28285 ^ t28285;
    wire t28287 = t28286 ^ t28286;
    wire t28288 = t28287 ^ t28287;
    wire t28289 = t28288 ^ t28288;
    wire t28290 = t28289 ^ t28289;
    wire t28291 = t28290 ^ t28290;
    wire t28292 = t28291 ^ t28291;
    wire t28293 = t28292 ^ t28292;
    wire t28294 = t28293 ^ t28293;
    wire t28295 = t28294 ^ t28294;
    wire t28296 = t28295 ^ t28295;
    wire t28297 = t28296 ^ t28296;
    wire t28298 = t28297 ^ t28297;
    wire t28299 = t28298 ^ t28298;
    wire t28300 = t28299 ^ t28299;
    wire t28301 = t28300 ^ t28300;
    wire t28302 = t28301 ^ t28301;
    wire t28303 = t28302 ^ t28302;
    wire t28304 = t28303 ^ t28303;
    wire t28305 = t28304 ^ t28304;
    wire t28306 = t28305 ^ t28305;
    wire t28307 = t28306 ^ t28306;
    wire t28308 = t28307 ^ t28307;
    wire t28309 = t28308 ^ t28308;
    wire t28310 = t28309 ^ t28309;
    wire t28311 = t28310 ^ t28310;
    wire t28312 = t28311 ^ t28311;
    wire t28313 = t28312 ^ t28312;
    wire t28314 = t28313 ^ t28313;
    wire t28315 = t28314 ^ t28314;
    wire t28316 = t28315 ^ t28315;
    wire t28317 = t28316 ^ t28316;
    wire t28318 = t28317 ^ t28317;
    wire t28319 = t28318 ^ t28318;
    wire t28320 = t28319 ^ t28319;
    wire t28321 = t28320 ^ t28320;
    wire t28322 = t28321 ^ t28321;
    wire t28323 = t28322 ^ t28322;
    wire t28324 = t28323 ^ t28323;
    wire t28325 = t28324 ^ t28324;
    wire t28326 = t28325 ^ t28325;
    wire t28327 = t28326 ^ t28326;
    wire t28328 = t28327 ^ t28327;
    wire t28329 = t28328 ^ t28328;
    wire t28330 = t28329 ^ t28329;
    wire t28331 = t28330 ^ t28330;
    wire t28332 = t28331 ^ t28331;
    wire t28333 = t28332 ^ t28332;
    wire t28334 = t28333 ^ t28333;
    wire t28335 = t28334 ^ t28334;
    wire t28336 = t28335 ^ t28335;
    wire t28337 = t28336 ^ t28336;
    wire t28338 = t28337 ^ t28337;
    wire t28339 = t28338 ^ t28338;
    wire t28340 = t28339 ^ t28339;
    wire t28341 = t28340 ^ t28340;
    wire t28342 = t28341 ^ t28341;
    wire t28343 = t28342 ^ t28342;
    wire t28344 = t28343 ^ t28343;
    wire t28345 = t28344 ^ t28344;
    wire t28346 = t28345 ^ t28345;
    wire t28347 = t28346 ^ t28346;
    wire t28348 = t28347 ^ t28347;
    wire t28349 = t28348 ^ t28348;
    wire t28350 = t28349 ^ t28349;
    wire t28351 = t28350 ^ t28350;
    wire t28352 = t28351 ^ t28351;
    wire t28353 = t28352 ^ t28352;
    wire t28354 = t28353 ^ t28353;
    wire t28355 = t28354 ^ t28354;
    wire t28356 = t28355 ^ t28355;
    wire t28357 = t28356 ^ t28356;
    wire t28358 = t28357 ^ t28357;
    wire t28359 = t28358 ^ t28358;
    wire t28360 = t28359 ^ t28359;
    wire t28361 = t28360 ^ t28360;
    wire t28362 = t28361 ^ t28361;
    wire t28363 = t28362 ^ t28362;
    wire t28364 = t28363 ^ t28363;
    wire t28365 = t28364 ^ t28364;
    wire t28366 = t28365 ^ t28365;
    wire t28367 = t28366 ^ t28366;
    wire t28368 = t28367 ^ t28367;
    wire t28369 = t28368 ^ t28368;
    wire t28370 = t28369 ^ t28369;
    wire t28371 = t28370 ^ t28370;
    wire t28372 = t28371 ^ t28371;
    wire t28373 = t28372 ^ t28372;
    wire t28374 = t28373 ^ t28373;
    wire t28375 = t28374 ^ t28374;
    wire t28376 = t28375 ^ t28375;
    wire t28377 = t28376 ^ t28376;
    wire t28378 = t28377 ^ t28377;
    wire t28379 = t28378 ^ t28378;
    wire t28380 = t28379 ^ t28379;
    wire t28381 = t28380 ^ t28380;
    wire t28382 = t28381 ^ t28381;
    wire t28383 = t28382 ^ t28382;
    wire t28384 = t28383 ^ t28383;
    wire t28385 = t28384 ^ t28384;
    wire t28386 = t28385 ^ t28385;
    wire t28387 = t28386 ^ t28386;
    wire t28388 = t28387 ^ t28387;
    wire t28389 = t28388 ^ t28388;
    wire t28390 = t28389 ^ t28389;
    wire t28391 = t28390 ^ t28390;
    wire t28392 = t28391 ^ t28391;
    wire t28393 = t28392 ^ t28392;
    wire t28394 = t28393 ^ t28393;
    wire t28395 = t28394 ^ t28394;
    wire t28396 = t28395 ^ t28395;
    wire t28397 = t28396 ^ t28396;
    wire t28398 = t28397 ^ t28397;
    wire t28399 = t28398 ^ t28398;
    wire t28400 = t28399 ^ t28399;
    wire t28401 = t28400 ^ t28400;
    wire t28402 = t28401 ^ t28401;
    wire t28403 = t28402 ^ t28402;
    wire t28404 = t28403 ^ t28403;
    wire t28405 = t28404 ^ t28404;
    wire t28406 = t28405 ^ t28405;
    wire t28407 = t28406 ^ t28406;
    wire t28408 = t28407 ^ t28407;
    wire t28409 = t28408 ^ t28408;
    wire t28410 = t28409 ^ t28409;
    wire t28411 = t28410 ^ t28410;
    wire t28412 = t28411 ^ t28411;
    wire t28413 = t28412 ^ t28412;
    wire t28414 = t28413 ^ t28413;
    wire t28415 = t28414 ^ t28414;
    wire t28416 = t28415 ^ t28415;
    wire t28417 = t28416 ^ t28416;
    wire t28418 = t28417 ^ t28417;
    wire t28419 = t28418 ^ t28418;
    wire t28420 = t28419 ^ t28419;
    wire t28421 = t28420 ^ t28420;
    wire t28422 = t28421 ^ t28421;
    wire t28423 = t28422 ^ t28422;
    wire t28424 = t28423 ^ t28423;
    wire t28425 = t28424 ^ t28424;
    wire t28426 = t28425 ^ t28425;
    wire t28427 = t28426 ^ t28426;
    wire t28428 = t28427 ^ t28427;
    wire t28429 = t28428 ^ t28428;
    wire t28430 = t28429 ^ t28429;
    wire t28431 = t28430 ^ t28430;
    wire t28432 = t28431 ^ t28431;
    wire t28433 = t28432 ^ t28432;
    wire t28434 = t28433 ^ t28433;
    wire t28435 = t28434 ^ t28434;
    wire t28436 = t28435 ^ t28435;
    wire t28437 = t28436 ^ t28436;
    wire t28438 = t28437 ^ t28437;
    wire t28439 = t28438 ^ t28438;
    wire t28440 = t28439 ^ t28439;
    wire t28441 = t28440 ^ t28440;
    wire t28442 = t28441 ^ t28441;
    wire t28443 = t28442 ^ t28442;
    wire t28444 = t28443 ^ t28443;
    wire t28445 = t28444 ^ t28444;
    wire t28446 = t28445 ^ t28445;
    wire t28447 = t28446 ^ t28446;
    wire t28448 = t28447 ^ t28447;
    wire t28449 = t28448 ^ t28448;
    wire t28450 = t28449 ^ t28449;
    wire t28451 = t28450 ^ t28450;
    wire t28452 = t28451 ^ t28451;
    wire t28453 = t28452 ^ t28452;
    wire t28454 = t28453 ^ t28453;
    wire t28455 = t28454 ^ t28454;
    wire t28456 = t28455 ^ t28455;
    wire t28457 = t28456 ^ t28456;
    wire t28458 = t28457 ^ t28457;
    wire t28459 = t28458 ^ t28458;
    wire t28460 = t28459 ^ t28459;
    wire t28461 = t28460 ^ t28460;
    wire t28462 = t28461 ^ t28461;
    wire t28463 = t28462 ^ t28462;
    wire t28464 = t28463 ^ t28463;
    wire t28465 = t28464 ^ t28464;
    wire t28466 = t28465 ^ t28465;
    wire t28467 = t28466 ^ t28466;
    wire t28468 = t28467 ^ t28467;
    wire t28469 = t28468 ^ t28468;
    wire t28470 = t28469 ^ t28469;
    wire t28471 = t28470 ^ t28470;
    wire t28472 = t28471 ^ t28471;
    wire t28473 = t28472 ^ t28472;
    wire t28474 = t28473 ^ t28473;
    wire t28475 = t28474 ^ t28474;
    wire t28476 = t28475 ^ t28475;
    wire t28477 = t28476 ^ t28476;
    wire t28478 = t28477 ^ t28477;
    wire t28479 = t28478 ^ t28478;
    wire t28480 = t28479 ^ t28479;
    wire t28481 = t28480 ^ t28480;
    wire t28482 = t28481 ^ t28481;
    wire t28483 = t28482 ^ t28482;
    wire t28484 = t28483 ^ t28483;
    wire t28485 = t28484 ^ t28484;
    wire t28486 = t28485 ^ t28485;
    wire t28487 = t28486 ^ t28486;
    wire t28488 = t28487 ^ t28487;
    wire t28489 = t28488 ^ t28488;
    wire t28490 = t28489 ^ t28489;
    wire t28491 = t28490 ^ t28490;
    wire t28492 = t28491 ^ t28491;
    wire t28493 = t28492 ^ t28492;
    wire t28494 = t28493 ^ t28493;
    wire t28495 = t28494 ^ t28494;
    wire t28496 = t28495 ^ t28495;
    wire t28497 = t28496 ^ t28496;
    wire t28498 = t28497 ^ t28497;
    wire t28499 = t28498 ^ t28498;
    wire t28500 = t28499 ^ t28499;
    wire t28501 = t28500 ^ t28500;
    wire t28502 = t28501 ^ t28501;
    wire t28503 = t28502 ^ t28502;
    wire t28504 = t28503 ^ t28503;
    wire t28505 = t28504 ^ t28504;
    wire t28506 = t28505 ^ t28505;
    wire t28507 = t28506 ^ t28506;
    wire t28508 = t28507 ^ t28507;
    wire t28509 = t28508 ^ t28508;
    wire t28510 = t28509 ^ t28509;
    wire t28511 = t28510 ^ t28510;
    wire t28512 = t28511 ^ t28511;
    wire t28513 = t28512 ^ t28512;
    wire t28514 = t28513 ^ t28513;
    wire t28515 = t28514 ^ t28514;
    wire t28516 = t28515 ^ t28515;
    wire t28517 = t28516 ^ t28516;
    wire t28518 = t28517 ^ t28517;
    wire t28519 = t28518 ^ t28518;
    wire t28520 = t28519 ^ t28519;
    wire t28521 = t28520 ^ t28520;
    wire t28522 = t28521 ^ t28521;
    wire t28523 = t28522 ^ t28522;
    wire t28524 = t28523 ^ t28523;
    wire t28525 = t28524 ^ t28524;
    wire t28526 = t28525 ^ t28525;
    wire t28527 = t28526 ^ t28526;
    wire t28528 = t28527 ^ t28527;
    wire t28529 = t28528 ^ t28528;
    wire t28530 = t28529 ^ t28529;
    wire t28531 = t28530 ^ t28530;
    wire t28532 = t28531 ^ t28531;
    wire t28533 = t28532 ^ t28532;
    wire t28534 = t28533 ^ t28533;
    wire t28535 = t28534 ^ t28534;
    wire t28536 = t28535 ^ t28535;
    wire t28537 = t28536 ^ t28536;
    wire t28538 = t28537 ^ t28537;
    wire t28539 = t28538 ^ t28538;
    wire t28540 = t28539 ^ t28539;
    wire t28541 = t28540 ^ t28540;
    wire t28542 = t28541 ^ t28541;
    wire t28543 = t28542 ^ t28542;
    wire t28544 = t28543 ^ t28543;
    wire t28545 = t28544 ^ t28544;
    wire t28546 = t28545 ^ t28545;
    wire t28547 = t28546 ^ t28546;
    wire t28548 = t28547 ^ t28547;
    wire t28549 = t28548 ^ t28548;
    wire t28550 = t28549 ^ t28549;
    wire t28551 = t28550 ^ t28550;
    wire t28552 = t28551 ^ t28551;
    wire t28553 = t28552 ^ t28552;
    wire t28554 = t28553 ^ t28553;
    wire t28555 = t28554 ^ t28554;
    wire t28556 = t28555 ^ t28555;
    wire t28557 = t28556 ^ t28556;
    wire t28558 = t28557 ^ t28557;
    wire t28559 = t28558 ^ t28558;
    wire t28560 = t28559 ^ t28559;
    wire t28561 = t28560 ^ t28560;
    wire t28562 = t28561 ^ t28561;
    wire t28563 = t28562 ^ t28562;
    wire t28564 = t28563 ^ t28563;
    wire t28565 = t28564 ^ t28564;
    wire t28566 = t28565 ^ t28565;
    wire t28567 = t28566 ^ t28566;
    wire t28568 = t28567 ^ t28567;
    wire t28569 = t28568 ^ t28568;
    wire t28570 = t28569 ^ t28569;
    wire t28571 = t28570 ^ t28570;
    wire t28572 = t28571 ^ t28571;
    wire t28573 = t28572 ^ t28572;
    wire t28574 = t28573 ^ t28573;
    wire t28575 = t28574 ^ t28574;
    wire t28576 = t28575 ^ t28575;
    wire t28577 = t28576 ^ t28576;
    wire t28578 = t28577 ^ t28577;
    wire t28579 = t28578 ^ t28578;
    wire t28580 = t28579 ^ t28579;
    wire t28581 = t28580 ^ t28580;
    wire t28582 = t28581 ^ t28581;
    wire t28583 = t28582 ^ t28582;
    wire t28584 = t28583 ^ t28583;
    wire t28585 = t28584 ^ t28584;
    wire t28586 = t28585 ^ t28585;
    wire t28587 = t28586 ^ t28586;
    wire t28588 = t28587 ^ t28587;
    wire t28589 = t28588 ^ t28588;
    wire t28590 = t28589 ^ t28589;
    wire t28591 = t28590 ^ t28590;
    wire t28592 = t28591 ^ t28591;
    wire t28593 = t28592 ^ t28592;
    wire t28594 = t28593 ^ t28593;
    wire t28595 = t28594 ^ t28594;
    wire t28596 = t28595 ^ t28595;
    wire t28597 = t28596 ^ t28596;
    wire t28598 = t28597 ^ t28597;
    wire t28599 = t28598 ^ t28598;
    wire t28600 = t28599 ^ t28599;
    wire t28601 = t28600 ^ t28600;
    wire t28602 = t28601 ^ t28601;
    wire t28603 = t28602 ^ t28602;
    wire t28604 = t28603 ^ t28603;
    wire t28605 = t28604 ^ t28604;
    wire t28606 = t28605 ^ t28605;
    wire t28607 = t28606 ^ t28606;
    wire t28608 = t28607 ^ t28607;
    wire t28609 = t28608 ^ t28608;
    wire t28610 = t28609 ^ t28609;
    wire t28611 = t28610 ^ t28610;
    wire t28612 = t28611 ^ t28611;
    wire t28613 = t28612 ^ t28612;
    wire t28614 = t28613 ^ t28613;
    wire t28615 = t28614 ^ t28614;
    wire t28616 = t28615 ^ t28615;
    wire t28617 = t28616 ^ t28616;
    wire t28618 = t28617 ^ t28617;
    wire t28619 = t28618 ^ t28618;
    wire t28620 = t28619 ^ t28619;
    wire t28621 = t28620 ^ t28620;
    wire t28622 = t28621 ^ t28621;
    wire t28623 = t28622 ^ t28622;
    wire t28624 = t28623 ^ t28623;
    wire t28625 = t28624 ^ t28624;
    wire t28626 = t28625 ^ t28625;
    wire t28627 = t28626 ^ t28626;
    wire t28628 = t28627 ^ t28627;
    wire t28629 = t28628 ^ t28628;
    wire t28630 = t28629 ^ t28629;
    wire t28631 = t28630 ^ t28630;
    wire t28632 = t28631 ^ t28631;
    wire t28633 = t28632 ^ t28632;
    wire t28634 = t28633 ^ t28633;
    wire t28635 = t28634 ^ t28634;
    wire t28636 = t28635 ^ t28635;
    wire t28637 = t28636 ^ t28636;
    wire t28638 = t28637 ^ t28637;
    wire t28639 = t28638 ^ t28638;
    wire t28640 = t28639 ^ t28639;
    wire t28641 = t28640 ^ t28640;
    wire t28642 = t28641 ^ t28641;
    wire t28643 = t28642 ^ t28642;
    wire t28644 = t28643 ^ t28643;
    wire t28645 = t28644 ^ t28644;
    wire t28646 = t28645 ^ t28645;
    wire t28647 = t28646 ^ t28646;
    wire t28648 = t28647 ^ t28647;
    wire t28649 = t28648 ^ t28648;
    wire t28650 = t28649 ^ t28649;
    wire t28651 = t28650 ^ t28650;
    wire t28652 = t28651 ^ t28651;
    wire t28653 = t28652 ^ t28652;
    wire t28654 = t28653 ^ t28653;
    wire t28655 = t28654 ^ t28654;
    wire t28656 = t28655 ^ t28655;
    wire t28657 = t28656 ^ t28656;
    wire t28658 = t28657 ^ t28657;
    wire t28659 = t28658 ^ t28658;
    wire t28660 = t28659 ^ t28659;
    wire t28661 = t28660 ^ t28660;
    wire t28662 = t28661 ^ t28661;
    wire t28663 = t28662 ^ t28662;
    wire t28664 = t28663 ^ t28663;
    wire t28665 = t28664 ^ t28664;
    wire t28666 = t28665 ^ t28665;
    wire t28667 = t28666 ^ t28666;
    wire t28668 = t28667 ^ t28667;
    wire t28669 = t28668 ^ t28668;
    wire t28670 = t28669 ^ t28669;
    wire t28671 = t28670 ^ t28670;
    wire t28672 = t28671 ^ t28671;
    wire t28673 = t28672 ^ t28672;
    wire t28674 = t28673 ^ t28673;
    wire t28675 = t28674 ^ t28674;
    wire t28676 = t28675 ^ t28675;
    wire t28677 = t28676 ^ t28676;
    wire t28678 = t28677 ^ t28677;
    wire t28679 = t28678 ^ t28678;
    wire t28680 = t28679 ^ t28679;
    wire t28681 = t28680 ^ t28680;
    wire t28682 = t28681 ^ t28681;
    wire t28683 = t28682 ^ t28682;
    wire t28684 = t28683 ^ t28683;
    wire t28685 = t28684 ^ t28684;
    wire t28686 = t28685 ^ t28685;
    wire t28687 = t28686 ^ t28686;
    wire t28688 = t28687 ^ t28687;
    wire t28689 = t28688 ^ t28688;
    wire t28690 = t28689 ^ t28689;
    wire t28691 = t28690 ^ t28690;
    wire t28692 = t28691 ^ t28691;
    wire t28693 = t28692 ^ t28692;
    wire t28694 = t28693 ^ t28693;
    wire t28695 = t28694 ^ t28694;
    wire t28696 = t28695 ^ t28695;
    wire t28697 = t28696 ^ t28696;
    wire t28698 = t28697 ^ t28697;
    wire t28699 = t28698 ^ t28698;
    wire t28700 = t28699 ^ t28699;
    wire t28701 = t28700 ^ t28700;
    wire t28702 = t28701 ^ t28701;
    wire t28703 = t28702 ^ t28702;
    wire t28704 = t28703 ^ t28703;
    wire t28705 = t28704 ^ t28704;
    wire t28706 = t28705 ^ t28705;
    wire t28707 = t28706 ^ t28706;
    wire t28708 = t28707 ^ t28707;
    wire t28709 = t28708 ^ t28708;
    wire t28710 = t28709 ^ t28709;
    wire t28711 = t28710 ^ t28710;
    wire t28712 = t28711 ^ t28711;
    wire t28713 = t28712 ^ t28712;
    wire t28714 = t28713 ^ t28713;
    wire t28715 = t28714 ^ t28714;
    wire t28716 = t28715 ^ t28715;
    wire t28717 = t28716 ^ t28716;
    wire t28718 = t28717 ^ t28717;
    wire t28719 = t28718 ^ t28718;
    wire t28720 = t28719 ^ t28719;
    wire t28721 = t28720 ^ t28720;
    wire t28722 = t28721 ^ t28721;
    wire t28723 = t28722 ^ t28722;
    wire t28724 = t28723 ^ t28723;
    wire t28725 = t28724 ^ t28724;
    wire t28726 = t28725 ^ t28725;
    wire t28727 = t28726 ^ t28726;
    wire t28728 = t28727 ^ t28727;
    wire t28729 = t28728 ^ t28728;
    wire t28730 = t28729 ^ t28729;
    wire t28731 = t28730 ^ t28730;
    wire t28732 = t28731 ^ t28731;
    wire t28733 = t28732 ^ t28732;
    wire t28734 = t28733 ^ t28733;
    wire t28735 = t28734 ^ t28734;
    wire t28736 = t28735 ^ t28735;
    wire t28737 = t28736 ^ t28736;
    wire t28738 = t28737 ^ t28737;
    wire t28739 = t28738 ^ t28738;
    wire t28740 = t28739 ^ t28739;
    wire t28741 = t28740 ^ t28740;
    wire t28742 = t28741 ^ t28741;
    wire t28743 = t28742 ^ t28742;
    wire t28744 = t28743 ^ t28743;
    wire t28745 = t28744 ^ t28744;
    wire t28746 = t28745 ^ t28745;
    wire t28747 = t28746 ^ t28746;
    wire t28748 = t28747 ^ t28747;
    wire t28749 = t28748 ^ t28748;
    wire t28750 = t28749 ^ t28749;
    wire t28751 = t28750 ^ t28750;
    wire t28752 = t28751 ^ t28751;
    wire t28753 = t28752 ^ t28752;
    wire t28754 = t28753 ^ t28753;
    wire t28755 = t28754 ^ t28754;
    wire t28756 = t28755 ^ t28755;
    wire t28757 = t28756 ^ t28756;
    wire t28758 = t28757 ^ t28757;
    wire t28759 = t28758 ^ t28758;
    wire t28760 = t28759 ^ t28759;
    wire t28761 = t28760 ^ t28760;
    wire t28762 = t28761 ^ t28761;
    wire t28763 = t28762 ^ t28762;
    wire t28764 = t28763 ^ t28763;
    wire t28765 = t28764 ^ t28764;
    wire t28766 = t28765 ^ t28765;
    wire t28767 = t28766 ^ t28766;
    wire t28768 = t28767 ^ t28767;
    wire t28769 = t28768 ^ t28768;
    wire t28770 = t28769 ^ t28769;
    wire t28771 = t28770 ^ t28770;
    wire t28772 = t28771 ^ t28771;
    wire t28773 = t28772 ^ t28772;
    wire t28774 = t28773 ^ t28773;
    wire t28775 = t28774 ^ t28774;
    wire t28776 = t28775 ^ t28775;
    wire t28777 = t28776 ^ t28776;
    wire t28778 = t28777 ^ t28777;
    wire t28779 = t28778 ^ t28778;
    wire t28780 = t28779 ^ t28779;
    wire t28781 = t28780 ^ t28780;
    wire t28782 = t28781 ^ t28781;
    wire t28783 = t28782 ^ t28782;
    wire t28784 = t28783 ^ t28783;
    wire t28785 = t28784 ^ t28784;
    wire t28786 = t28785 ^ t28785;
    wire t28787 = t28786 ^ t28786;
    wire t28788 = t28787 ^ t28787;
    wire t28789 = t28788 ^ t28788;
    wire t28790 = t28789 ^ t28789;
    wire t28791 = t28790 ^ t28790;
    wire t28792 = t28791 ^ t28791;
    wire t28793 = t28792 ^ t28792;
    wire t28794 = t28793 ^ t28793;
    wire t28795 = t28794 ^ t28794;
    wire t28796 = t28795 ^ t28795;
    wire t28797 = t28796 ^ t28796;
    wire t28798 = t28797 ^ t28797;
    wire t28799 = t28798 ^ t28798;
    wire t28800 = t28799 ^ t28799;
    wire t28801 = t28800 ^ t28800;
    wire t28802 = t28801 ^ t28801;
    wire t28803 = t28802 ^ t28802;
    wire t28804 = t28803 ^ t28803;
    wire t28805 = t28804 ^ t28804;
    wire t28806 = t28805 ^ t28805;
    wire t28807 = t28806 ^ t28806;
    wire t28808 = t28807 ^ t28807;
    wire t28809 = t28808 ^ t28808;
    wire t28810 = t28809 ^ t28809;
    wire t28811 = t28810 ^ t28810;
    wire t28812 = t28811 ^ t28811;
    wire t28813 = t28812 ^ t28812;
    wire t28814 = t28813 ^ t28813;
    wire t28815 = t28814 ^ t28814;
    wire t28816 = t28815 ^ t28815;
    wire t28817 = t28816 ^ t28816;
    wire t28818 = t28817 ^ t28817;
    wire t28819 = t28818 ^ t28818;
    wire t28820 = t28819 ^ t28819;
    wire t28821 = t28820 ^ t28820;
    wire t28822 = t28821 ^ t28821;
    wire t28823 = t28822 ^ t28822;
    wire t28824 = t28823 ^ t28823;
    wire t28825 = t28824 ^ t28824;
    wire t28826 = t28825 ^ t28825;
    wire t28827 = t28826 ^ t28826;
    wire t28828 = t28827 ^ t28827;
    wire t28829 = t28828 ^ t28828;
    wire t28830 = t28829 ^ t28829;
    wire t28831 = t28830 ^ t28830;
    wire t28832 = t28831 ^ t28831;
    wire t28833 = t28832 ^ t28832;
    wire t28834 = t28833 ^ t28833;
    wire t28835 = t28834 ^ t28834;
    wire t28836 = t28835 ^ t28835;
    wire t28837 = t28836 ^ t28836;
    wire t28838 = t28837 ^ t28837;
    wire t28839 = t28838 ^ t28838;
    wire t28840 = t28839 ^ t28839;
    wire t28841 = t28840 ^ t28840;
    wire t28842 = t28841 ^ t28841;
    wire t28843 = t28842 ^ t28842;
    wire t28844 = t28843 ^ t28843;
    wire t28845 = t28844 ^ t28844;
    wire t28846 = t28845 ^ t28845;
    wire t28847 = t28846 ^ t28846;
    wire t28848 = t28847 ^ t28847;
    wire t28849 = t28848 ^ t28848;
    wire t28850 = t28849 ^ t28849;
    wire t28851 = t28850 ^ t28850;
    wire t28852 = t28851 ^ t28851;
    wire t28853 = t28852 ^ t28852;
    wire t28854 = t28853 ^ t28853;
    wire t28855 = t28854 ^ t28854;
    wire t28856 = t28855 ^ t28855;
    wire t28857 = t28856 ^ t28856;
    wire t28858 = t28857 ^ t28857;
    wire t28859 = t28858 ^ t28858;
    wire t28860 = t28859 ^ t28859;
    wire t28861 = t28860 ^ t28860;
    wire t28862 = t28861 ^ t28861;
    wire t28863 = t28862 ^ t28862;
    wire t28864 = t28863 ^ t28863;
    wire t28865 = t28864 ^ t28864;
    wire t28866 = t28865 ^ t28865;
    wire t28867 = t28866 ^ t28866;
    wire t28868 = t28867 ^ t28867;
    wire t28869 = t28868 ^ t28868;
    wire t28870 = t28869 ^ t28869;
    wire t28871 = t28870 ^ t28870;
    wire t28872 = t28871 ^ t28871;
    wire t28873 = t28872 ^ t28872;
    wire t28874 = t28873 ^ t28873;
    wire t28875 = t28874 ^ t28874;
    wire t28876 = t28875 ^ t28875;
    wire t28877 = t28876 ^ t28876;
    wire t28878 = t28877 ^ t28877;
    wire t28879 = t28878 ^ t28878;
    wire t28880 = t28879 ^ t28879;
    wire t28881 = t28880 ^ t28880;
    wire t28882 = t28881 ^ t28881;
    wire t28883 = t28882 ^ t28882;
    wire t28884 = t28883 ^ t28883;
    wire t28885 = t28884 ^ t28884;
    wire t28886 = t28885 ^ t28885;
    wire t28887 = t28886 ^ t28886;
    wire t28888 = t28887 ^ t28887;
    wire t28889 = t28888 ^ t28888;
    wire t28890 = t28889 ^ t28889;
    wire t28891 = t28890 ^ t28890;
    wire t28892 = t28891 ^ t28891;
    wire t28893 = t28892 ^ t28892;
    wire t28894 = t28893 ^ t28893;
    wire t28895 = t28894 ^ t28894;
    wire t28896 = t28895 ^ t28895;
    wire t28897 = t28896 ^ t28896;
    wire t28898 = t28897 ^ t28897;
    wire t28899 = t28898 ^ t28898;
    wire t28900 = t28899 ^ t28899;
    wire t28901 = t28900 ^ t28900;
    wire t28902 = t28901 ^ t28901;
    wire t28903 = t28902 ^ t28902;
    wire t28904 = t28903 ^ t28903;
    wire t28905 = t28904 ^ t28904;
    wire t28906 = t28905 ^ t28905;
    wire t28907 = t28906 ^ t28906;
    wire t28908 = t28907 ^ t28907;
    wire t28909 = t28908 ^ t28908;
    wire t28910 = t28909 ^ t28909;
    wire t28911 = t28910 ^ t28910;
    wire t28912 = t28911 ^ t28911;
    wire t28913 = t28912 ^ t28912;
    wire t28914 = t28913 ^ t28913;
    wire t28915 = t28914 ^ t28914;
    wire t28916 = t28915 ^ t28915;
    wire t28917 = t28916 ^ t28916;
    wire t28918 = t28917 ^ t28917;
    wire t28919 = t28918 ^ t28918;
    wire t28920 = t28919 ^ t28919;
    wire t28921 = t28920 ^ t28920;
    wire t28922 = t28921 ^ t28921;
    wire t28923 = t28922 ^ t28922;
    wire t28924 = t28923 ^ t28923;
    wire t28925 = t28924 ^ t28924;
    wire t28926 = t28925 ^ t28925;
    wire t28927 = t28926 ^ t28926;
    wire t28928 = t28927 ^ t28927;
    wire t28929 = t28928 ^ t28928;
    wire t28930 = t28929 ^ t28929;
    wire t28931 = t28930 ^ t28930;
    wire t28932 = t28931 ^ t28931;
    wire t28933 = t28932 ^ t28932;
    wire t28934 = t28933 ^ t28933;
    wire t28935 = t28934 ^ t28934;
    wire t28936 = t28935 ^ t28935;
    wire t28937 = t28936 ^ t28936;
    wire t28938 = t28937 ^ t28937;
    wire t28939 = t28938 ^ t28938;
    wire t28940 = t28939 ^ t28939;
    wire t28941 = t28940 ^ t28940;
    wire t28942 = t28941 ^ t28941;
    wire t28943 = t28942 ^ t28942;
    wire t28944 = t28943 ^ t28943;
    wire t28945 = t28944 ^ t28944;
    wire t28946 = t28945 ^ t28945;
    wire t28947 = t28946 ^ t28946;
    wire t28948 = t28947 ^ t28947;
    wire t28949 = t28948 ^ t28948;
    wire t28950 = t28949 ^ t28949;
    wire t28951 = t28950 ^ t28950;
    wire t28952 = t28951 ^ t28951;
    wire t28953 = t28952 ^ t28952;
    wire t28954 = t28953 ^ t28953;
    wire t28955 = t28954 ^ t28954;
    wire t28956 = t28955 ^ t28955;
    wire t28957 = t28956 ^ t28956;
    wire t28958 = t28957 ^ t28957;
    wire t28959 = t28958 ^ t28958;
    wire t28960 = t28959 ^ t28959;
    wire t28961 = t28960 ^ t28960;
    wire t28962 = t28961 ^ t28961;
    wire t28963 = t28962 ^ t28962;
    wire t28964 = t28963 ^ t28963;
    wire t28965 = t28964 ^ t28964;
    wire t28966 = t28965 ^ t28965;
    wire t28967 = t28966 ^ t28966;
    wire t28968 = t28967 ^ t28967;
    wire t28969 = t28968 ^ t28968;
    wire t28970 = t28969 ^ t28969;
    wire t28971 = t28970 ^ t28970;
    wire t28972 = t28971 ^ t28971;
    wire t28973 = t28972 ^ t28972;
    wire t28974 = t28973 ^ t28973;
    wire t28975 = t28974 ^ t28974;
    wire t28976 = t28975 ^ t28975;
    wire t28977 = t28976 ^ t28976;
    wire t28978 = t28977 ^ t28977;
    wire t28979 = t28978 ^ t28978;
    wire t28980 = t28979 ^ t28979;
    wire t28981 = t28980 ^ t28980;
    wire t28982 = t28981 ^ t28981;
    wire t28983 = t28982 ^ t28982;
    wire t28984 = t28983 ^ t28983;
    wire t28985 = t28984 ^ t28984;
    wire t28986 = t28985 ^ t28985;
    wire t28987 = t28986 ^ t28986;
    wire t28988 = t28987 ^ t28987;
    wire t28989 = t28988 ^ t28988;
    wire t28990 = t28989 ^ t28989;
    wire t28991 = t28990 ^ t28990;
    wire t28992 = t28991 ^ t28991;
    wire t28993 = t28992 ^ t28992;
    wire t28994 = t28993 ^ t28993;
    wire t28995 = t28994 ^ t28994;
    wire t28996 = t28995 ^ t28995;
    wire t28997 = t28996 ^ t28996;
    wire t28998 = t28997 ^ t28997;
    wire t28999 = t28998 ^ t28998;
    wire t29000 = t28999 ^ t28999;
    wire t29001 = t29000 ^ t29000;
    wire t29002 = t29001 ^ t29001;
    wire t29003 = t29002 ^ t29002;
    wire t29004 = t29003 ^ t29003;
    wire t29005 = t29004 ^ t29004;
    wire t29006 = t29005 ^ t29005;
    wire t29007 = t29006 ^ t29006;
    wire t29008 = t29007 ^ t29007;
    wire t29009 = t29008 ^ t29008;
    wire t29010 = t29009 ^ t29009;
    wire t29011 = t29010 ^ t29010;
    wire t29012 = t29011 ^ t29011;
    wire t29013 = t29012 ^ t29012;
    wire t29014 = t29013 ^ t29013;
    wire t29015 = t29014 ^ t29014;
    wire t29016 = t29015 ^ t29015;
    wire t29017 = t29016 ^ t29016;
    wire t29018 = t29017 ^ t29017;
    wire t29019 = t29018 ^ t29018;
    wire t29020 = t29019 ^ t29019;
    wire t29021 = t29020 ^ t29020;
    wire t29022 = t29021 ^ t29021;
    wire t29023 = t29022 ^ t29022;
    wire t29024 = t29023 ^ t29023;
    wire t29025 = t29024 ^ t29024;
    wire t29026 = t29025 ^ t29025;
    wire t29027 = t29026 ^ t29026;
    wire t29028 = t29027 ^ t29027;
    wire t29029 = t29028 ^ t29028;
    wire t29030 = t29029 ^ t29029;
    wire t29031 = t29030 ^ t29030;
    wire t29032 = t29031 ^ t29031;
    wire t29033 = t29032 ^ t29032;
    wire t29034 = t29033 ^ t29033;
    wire t29035 = t29034 ^ t29034;
    wire t29036 = t29035 ^ t29035;
    wire t29037 = t29036 ^ t29036;
    wire t29038 = t29037 ^ t29037;
    wire t29039 = t29038 ^ t29038;
    wire t29040 = t29039 ^ t29039;
    wire t29041 = t29040 ^ t29040;
    wire t29042 = t29041 ^ t29041;
    wire t29043 = t29042 ^ t29042;
    wire t29044 = t29043 ^ t29043;
    wire t29045 = t29044 ^ t29044;
    wire t29046 = t29045 ^ t29045;
    wire t29047 = t29046 ^ t29046;
    wire t29048 = t29047 ^ t29047;
    wire t29049 = t29048 ^ t29048;
    wire t29050 = t29049 ^ t29049;
    wire t29051 = t29050 ^ t29050;
    wire t29052 = t29051 ^ t29051;
    wire t29053 = t29052 ^ t29052;
    wire t29054 = t29053 ^ t29053;
    wire t29055 = t29054 ^ t29054;
    wire t29056 = t29055 ^ t29055;
    wire t29057 = t29056 ^ t29056;
    wire t29058 = t29057 ^ t29057;
    wire t29059 = t29058 ^ t29058;
    wire t29060 = t29059 ^ t29059;
    wire t29061 = t29060 ^ t29060;
    wire t29062 = t29061 ^ t29061;
    wire t29063 = t29062 ^ t29062;
    wire t29064 = t29063 ^ t29063;
    wire t29065 = t29064 ^ t29064;
    wire t29066 = t29065 ^ t29065;
    wire t29067 = t29066 ^ t29066;
    wire t29068 = t29067 ^ t29067;
    wire t29069 = t29068 ^ t29068;
    wire t29070 = t29069 ^ t29069;
    wire t29071 = t29070 ^ t29070;
    wire t29072 = t29071 ^ t29071;
    wire t29073 = t29072 ^ t29072;
    wire t29074 = t29073 ^ t29073;
    wire t29075 = t29074 ^ t29074;
    wire t29076 = t29075 ^ t29075;
    wire t29077 = t29076 ^ t29076;
    wire t29078 = t29077 ^ t29077;
    wire t29079 = t29078 ^ t29078;
    wire t29080 = t29079 ^ t29079;
    wire t29081 = t29080 ^ t29080;
    wire t29082 = t29081 ^ t29081;
    wire t29083 = t29082 ^ t29082;
    wire t29084 = t29083 ^ t29083;
    wire t29085 = t29084 ^ t29084;
    wire t29086 = t29085 ^ t29085;
    wire t29087 = t29086 ^ t29086;
    wire t29088 = t29087 ^ t29087;
    wire t29089 = t29088 ^ t29088;
    wire t29090 = t29089 ^ t29089;
    wire t29091 = t29090 ^ t29090;
    wire t29092 = t29091 ^ t29091;
    wire t29093 = t29092 ^ t29092;
    wire t29094 = t29093 ^ t29093;
    wire t29095 = t29094 ^ t29094;
    wire t29096 = t29095 ^ t29095;
    wire t29097 = t29096 ^ t29096;
    wire t29098 = t29097 ^ t29097;
    wire t29099 = t29098 ^ t29098;
    wire t29100 = t29099 ^ t29099;
    wire t29101 = t29100 ^ t29100;
    wire t29102 = t29101 ^ t29101;
    wire t29103 = t29102 ^ t29102;
    wire t29104 = t29103 ^ t29103;
    wire t29105 = t29104 ^ t29104;
    wire t29106 = t29105 ^ t29105;
    wire t29107 = t29106 ^ t29106;
    wire t29108 = t29107 ^ t29107;
    wire t29109 = t29108 ^ t29108;
    wire t29110 = t29109 ^ t29109;
    wire t29111 = t29110 ^ t29110;
    wire t29112 = t29111 ^ t29111;
    wire t29113 = t29112 ^ t29112;
    wire t29114 = t29113 ^ t29113;
    wire t29115 = t29114 ^ t29114;
    wire t29116 = t29115 ^ t29115;
    wire t29117 = t29116 ^ t29116;
    wire t29118 = t29117 ^ t29117;
    wire t29119 = t29118 ^ t29118;
    wire t29120 = t29119 ^ t29119;
    wire t29121 = t29120 ^ t29120;
    wire t29122 = t29121 ^ t29121;
    wire t29123 = t29122 ^ t29122;
    wire t29124 = t29123 ^ t29123;
    wire t29125 = t29124 ^ t29124;
    wire t29126 = t29125 ^ t29125;
    wire t29127 = t29126 ^ t29126;
    wire t29128 = t29127 ^ t29127;
    wire t29129 = t29128 ^ t29128;
    wire t29130 = t29129 ^ t29129;
    wire t29131 = t29130 ^ t29130;
    wire t29132 = t29131 ^ t29131;
    wire t29133 = t29132 ^ t29132;
    wire t29134 = t29133 ^ t29133;
    wire t29135 = t29134 ^ t29134;
    wire t29136 = t29135 ^ t29135;
    wire t29137 = t29136 ^ t29136;
    wire t29138 = t29137 ^ t29137;
    wire t29139 = t29138 ^ t29138;
    wire t29140 = t29139 ^ t29139;
    wire t29141 = t29140 ^ t29140;
    wire t29142 = t29141 ^ t29141;
    wire t29143 = t29142 ^ t29142;
    wire t29144 = t29143 ^ t29143;
    wire t29145 = t29144 ^ t29144;
    wire t29146 = t29145 ^ t29145;
    wire t29147 = t29146 ^ t29146;
    wire t29148 = t29147 ^ t29147;
    wire t29149 = t29148 ^ t29148;
    wire t29150 = t29149 ^ t29149;
    wire t29151 = t29150 ^ t29150;
    wire t29152 = t29151 ^ t29151;
    wire t29153 = t29152 ^ t29152;
    wire t29154 = t29153 ^ t29153;
    wire t29155 = t29154 ^ t29154;
    wire t29156 = t29155 ^ t29155;
    wire t29157 = t29156 ^ t29156;
    wire t29158 = t29157 ^ t29157;
    wire t29159 = t29158 ^ t29158;
    wire t29160 = t29159 ^ t29159;
    wire t29161 = t29160 ^ t29160;
    wire t29162 = t29161 ^ t29161;
    wire t29163 = t29162 ^ t29162;
    wire t29164 = t29163 ^ t29163;
    wire t29165 = t29164 ^ t29164;
    wire t29166 = t29165 ^ t29165;
    wire t29167 = t29166 ^ t29166;
    wire t29168 = t29167 ^ t29167;
    wire t29169 = t29168 ^ t29168;
    wire t29170 = t29169 ^ t29169;
    wire t29171 = t29170 ^ t29170;
    wire t29172 = t29171 ^ t29171;
    wire t29173 = t29172 ^ t29172;
    wire t29174 = t29173 ^ t29173;
    wire t29175 = t29174 ^ t29174;
    wire t29176 = t29175 ^ t29175;
    wire t29177 = t29176 ^ t29176;
    wire t29178 = t29177 ^ t29177;
    wire t29179 = t29178 ^ t29178;
    wire t29180 = t29179 ^ t29179;
    wire t29181 = t29180 ^ t29180;
    wire t29182 = t29181 ^ t29181;
    wire t29183 = t29182 ^ t29182;
    wire t29184 = t29183 ^ t29183;
    wire t29185 = t29184 ^ t29184;
    wire t29186 = t29185 ^ t29185;
    wire t29187 = t29186 ^ t29186;
    wire t29188 = t29187 ^ t29187;
    wire t29189 = t29188 ^ t29188;
    wire t29190 = t29189 ^ t29189;
    wire t29191 = t29190 ^ t29190;
    wire t29192 = t29191 ^ t29191;
    wire t29193 = t29192 ^ t29192;
    wire t29194 = t29193 ^ t29193;
    wire t29195 = t29194 ^ t29194;
    wire t29196 = t29195 ^ t29195;
    wire t29197 = t29196 ^ t29196;
    wire t29198 = t29197 ^ t29197;
    wire t29199 = t29198 ^ t29198;
    wire t29200 = t29199 ^ t29199;
    wire t29201 = t29200 ^ t29200;
    wire t29202 = t29201 ^ t29201;
    wire t29203 = t29202 ^ t29202;
    wire t29204 = t29203 ^ t29203;
    wire t29205 = t29204 ^ t29204;
    wire t29206 = t29205 ^ t29205;
    wire t29207 = t29206 ^ t29206;
    wire t29208 = t29207 ^ t29207;
    wire t29209 = t29208 ^ t29208;
    wire t29210 = t29209 ^ t29209;
    wire t29211 = t29210 ^ t29210;
    wire t29212 = t29211 ^ t29211;
    wire t29213 = t29212 ^ t29212;
    wire t29214 = t29213 ^ t29213;
    wire t29215 = t29214 ^ t29214;
    wire t29216 = t29215 ^ t29215;
    wire t29217 = t29216 ^ t29216;
    wire t29218 = t29217 ^ t29217;
    wire t29219 = t29218 ^ t29218;
    wire t29220 = t29219 ^ t29219;
    wire t29221 = t29220 ^ t29220;
    wire t29222 = t29221 ^ t29221;
    wire t29223 = t29222 ^ t29222;
    wire t29224 = t29223 ^ t29223;
    wire t29225 = t29224 ^ t29224;
    wire t29226 = t29225 ^ t29225;
    wire t29227 = t29226 ^ t29226;
    wire t29228 = t29227 ^ t29227;
    wire t29229 = t29228 ^ t29228;
    wire t29230 = t29229 ^ t29229;
    wire t29231 = t29230 ^ t29230;
    wire t29232 = t29231 ^ t29231;
    wire t29233 = t29232 ^ t29232;
    wire t29234 = t29233 ^ t29233;
    wire t29235 = t29234 ^ t29234;
    wire t29236 = t29235 ^ t29235;
    wire t29237 = t29236 ^ t29236;
    wire t29238 = t29237 ^ t29237;
    wire t29239 = t29238 ^ t29238;
    wire t29240 = t29239 ^ t29239;
    wire t29241 = t29240 ^ t29240;
    wire t29242 = t29241 ^ t29241;
    wire t29243 = t29242 ^ t29242;
    wire t29244 = t29243 ^ t29243;
    wire t29245 = t29244 ^ t29244;
    wire t29246 = t29245 ^ t29245;
    wire t29247 = t29246 ^ t29246;
    wire t29248 = t29247 ^ t29247;
    wire t29249 = t29248 ^ t29248;
    wire t29250 = t29249 ^ t29249;
    wire t29251 = t29250 ^ t29250;
    wire t29252 = t29251 ^ t29251;
    wire t29253 = t29252 ^ t29252;
    wire t29254 = t29253 ^ t29253;
    wire t29255 = t29254 ^ t29254;
    wire t29256 = t29255 ^ t29255;
    wire t29257 = t29256 ^ t29256;
    wire t29258 = t29257 ^ t29257;
    wire t29259 = t29258 ^ t29258;
    wire t29260 = t29259 ^ t29259;
    wire t29261 = t29260 ^ t29260;
    wire t29262 = t29261 ^ t29261;
    wire t29263 = t29262 ^ t29262;
    wire t29264 = t29263 ^ t29263;
    wire t29265 = t29264 ^ t29264;
    wire t29266 = t29265 ^ t29265;
    wire t29267 = t29266 ^ t29266;
    wire t29268 = t29267 ^ t29267;
    wire t29269 = t29268 ^ t29268;
    wire t29270 = t29269 ^ t29269;
    wire t29271 = t29270 ^ t29270;
    wire t29272 = t29271 ^ t29271;
    wire t29273 = t29272 ^ t29272;
    wire t29274 = t29273 ^ t29273;
    wire t29275 = t29274 ^ t29274;
    wire t29276 = t29275 ^ t29275;
    wire t29277 = t29276 ^ t29276;
    wire t29278 = t29277 ^ t29277;
    wire t29279 = t29278 ^ t29278;
    wire t29280 = t29279 ^ t29279;
    wire t29281 = t29280 ^ t29280;
    wire t29282 = t29281 ^ t29281;
    wire t29283 = t29282 ^ t29282;
    wire t29284 = t29283 ^ t29283;
    wire t29285 = t29284 ^ t29284;
    wire t29286 = t29285 ^ t29285;
    wire t29287 = t29286 ^ t29286;
    wire t29288 = t29287 ^ t29287;
    wire t29289 = t29288 ^ t29288;
    wire t29290 = t29289 ^ t29289;
    wire t29291 = t29290 ^ t29290;
    wire t29292 = t29291 ^ t29291;
    wire t29293 = t29292 ^ t29292;
    wire t29294 = t29293 ^ t29293;
    wire t29295 = t29294 ^ t29294;
    wire t29296 = t29295 ^ t29295;
    wire t29297 = t29296 ^ t29296;
    wire t29298 = t29297 ^ t29297;
    wire t29299 = t29298 ^ t29298;
    wire t29300 = t29299 ^ t29299;
    wire t29301 = t29300 ^ t29300;
    wire t29302 = t29301 ^ t29301;
    wire t29303 = t29302 ^ t29302;
    wire t29304 = t29303 ^ t29303;
    wire t29305 = t29304 ^ t29304;
    wire t29306 = t29305 ^ t29305;
    wire t29307 = t29306 ^ t29306;
    wire t29308 = t29307 ^ t29307;
    wire t29309 = t29308 ^ t29308;
    wire t29310 = t29309 ^ t29309;
    wire t29311 = t29310 ^ t29310;
    wire t29312 = t29311 ^ t29311;
    wire t29313 = t29312 ^ t29312;
    wire t29314 = t29313 ^ t29313;
    wire t29315 = t29314 ^ t29314;
    wire t29316 = t29315 ^ t29315;
    wire t29317 = t29316 ^ t29316;
    wire t29318 = t29317 ^ t29317;
    wire t29319 = t29318 ^ t29318;
    wire t29320 = t29319 ^ t29319;
    wire t29321 = t29320 ^ t29320;
    wire t29322 = t29321 ^ t29321;
    wire t29323 = t29322 ^ t29322;
    wire t29324 = t29323 ^ t29323;
    wire t29325 = t29324 ^ t29324;
    wire t29326 = t29325 ^ t29325;
    wire t29327 = t29326 ^ t29326;
    wire t29328 = t29327 ^ t29327;
    wire t29329 = t29328 ^ t29328;
    wire t29330 = t29329 ^ t29329;
    wire t29331 = t29330 ^ t29330;
    wire t29332 = t29331 ^ t29331;
    wire t29333 = t29332 ^ t29332;
    wire t29334 = t29333 ^ t29333;
    wire t29335 = t29334 ^ t29334;
    wire t29336 = t29335 ^ t29335;
    wire t29337 = t29336 ^ t29336;
    wire t29338 = t29337 ^ t29337;
    wire t29339 = t29338 ^ t29338;
    wire t29340 = t29339 ^ t29339;
    wire t29341 = t29340 ^ t29340;
    wire t29342 = t29341 ^ t29341;
    wire t29343 = t29342 ^ t29342;
    wire t29344 = t29343 ^ t29343;
    wire t29345 = t29344 ^ t29344;
    wire t29346 = t29345 ^ t29345;
    wire t29347 = t29346 ^ t29346;
    wire t29348 = t29347 ^ t29347;
    wire t29349 = t29348 ^ t29348;
    wire t29350 = t29349 ^ t29349;
    wire t29351 = t29350 ^ t29350;
    wire t29352 = t29351 ^ t29351;
    wire t29353 = t29352 ^ t29352;
    wire t29354 = t29353 ^ t29353;
    wire t29355 = t29354 ^ t29354;
    wire t29356 = t29355 ^ t29355;
    wire t29357 = t29356 ^ t29356;
    wire t29358 = t29357 ^ t29357;
    wire t29359 = t29358 ^ t29358;
    wire t29360 = t29359 ^ t29359;
    wire t29361 = t29360 ^ t29360;
    wire t29362 = t29361 ^ t29361;
    wire t29363 = t29362 ^ t29362;
    wire t29364 = t29363 ^ t29363;
    wire t29365 = t29364 ^ t29364;
    wire t29366 = t29365 ^ t29365;
    wire t29367 = t29366 ^ t29366;
    wire t29368 = t29367 ^ t29367;
    wire t29369 = t29368 ^ t29368;
    wire t29370 = t29369 ^ t29369;
    wire t29371 = t29370 ^ t29370;
    wire t29372 = t29371 ^ t29371;
    wire t29373 = t29372 ^ t29372;
    wire t29374 = t29373 ^ t29373;
    wire t29375 = t29374 ^ t29374;
    wire t29376 = t29375 ^ t29375;
    wire t29377 = t29376 ^ t29376;
    wire t29378 = t29377 ^ t29377;
    wire t29379 = t29378 ^ t29378;
    wire t29380 = t29379 ^ t29379;
    wire t29381 = t29380 ^ t29380;
    wire t29382 = t29381 ^ t29381;
    wire t29383 = t29382 ^ t29382;
    wire t29384 = t29383 ^ t29383;
    wire t29385 = t29384 ^ t29384;
    wire t29386 = t29385 ^ t29385;
    wire t29387 = t29386 ^ t29386;
    wire t29388 = t29387 ^ t29387;
    wire t29389 = t29388 ^ t29388;
    wire t29390 = t29389 ^ t29389;
    wire t29391 = t29390 ^ t29390;
    wire t29392 = t29391 ^ t29391;
    wire t29393 = t29392 ^ t29392;
    wire t29394 = t29393 ^ t29393;
    wire t29395 = t29394 ^ t29394;
    wire t29396 = t29395 ^ t29395;
    wire t29397 = t29396 ^ t29396;
    wire t29398 = t29397 ^ t29397;
    wire t29399 = t29398 ^ t29398;
    wire t29400 = t29399 ^ t29399;
    wire t29401 = t29400 ^ t29400;
    wire t29402 = t29401 ^ t29401;
    wire t29403 = t29402 ^ t29402;
    wire t29404 = t29403 ^ t29403;
    wire t29405 = t29404 ^ t29404;
    wire t29406 = t29405 ^ t29405;
    wire t29407 = t29406 ^ t29406;
    wire t29408 = t29407 ^ t29407;
    wire t29409 = t29408 ^ t29408;
    wire t29410 = t29409 ^ t29409;
    wire t29411 = t29410 ^ t29410;
    wire t29412 = t29411 ^ t29411;
    wire t29413 = t29412 ^ t29412;
    wire t29414 = t29413 ^ t29413;
    wire t29415 = t29414 ^ t29414;
    wire t29416 = t29415 ^ t29415;
    wire t29417 = t29416 ^ t29416;
    wire t29418 = t29417 ^ t29417;
    wire t29419 = t29418 ^ t29418;
    wire t29420 = t29419 ^ t29419;
    wire t29421 = t29420 ^ t29420;
    wire t29422 = t29421 ^ t29421;
    wire t29423 = t29422 ^ t29422;
    wire t29424 = t29423 ^ t29423;
    wire t29425 = t29424 ^ t29424;
    wire t29426 = t29425 ^ t29425;
    wire t29427 = t29426 ^ t29426;
    wire t29428 = t29427 ^ t29427;
    wire t29429 = t29428 ^ t29428;
    wire t29430 = t29429 ^ t29429;
    wire t29431 = t29430 ^ t29430;
    wire t29432 = t29431 ^ t29431;
    wire t29433 = t29432 ^ t29432;
    wire t29434 = t29433 ^ t29433;
    wire t29435 = t29434 ^ t29434;
    wire t29436 = t29435 ^ t29435;
    wire t29437 = t29436 ^ t29436;
    wire t29438 = t29437 ^ t29437;
    wire t29439 = t29438 ^ t29438;
    wire t29440 = t29439 ^ t29439;
    wire t29441 = t29440 ^ t29440;
    wire t29442 = t29441 ^ t29441;
    wire t29443 = t29442 ^ t29442;
    wire t29444 = t29443 ^ t29443;
    wire t29445 = t29444 ^ t29444;
    wire t29446 = t29445 ^ t29445;
    wire t29447 = t29446 ^ t29446;
    wire t29448 = t29447 ^ t29447;
    wire t29449 = t29448 ^ t29448;
    wire t29450 = t29449 ^ t29449;
    wire t29451 = t29450 ^ t29450;
    wire t29452 = t29451 ^ t29451;
    wire t29453 = t29452 ^ t29452;
    wire t29454 = t29453 ^ t29453;
    wire t29455 = t29454 ^ t29454;
    wire t29456 = t29455 ^ t29455;
    wire t29457 = t29456 ^ t29456;
    wire t29458 = t29457 ^ t29457;
    wire t29459 = t29458 ^ t29458;
    wire t29460 = t29459 ^ t29459;
    wire t29461 = t29460 ^ t29460;
    wire t29462 = t29461 ^ t29461;
    wire t29463 = t29462 ^ t29462;
    wire t29464 = t29463 ^ t29463;
    wire t29465 = t29464 ^ t29464;
    wire t29466 = t29465 ^ t29465;
    wire t29467 = t29466 ^ t29466;
    wire t29468 = t29467 ^ t29467;
    wire t29469 = t29468 ^ t29468;
    wire t29470 = t29469 ^ t29469;
    wire t29471 = t29470 ^ t29470;
    wire t29472 = t29471 ^ t29471;
    wire t29473 = t29472 ^ t29472;
    wire t29474 = t29473 ^ t29473;
    wire t29475 = t29474 ^ t29474;
    wire t29476 = t29475 ^ t29475;
    wire t29477 = t29476 ^ t29476;
    wire t29478 = t29477 ^ t29477;
    wire t29479 = t29478 ^ t29478;
    wire t29480 = t29479 ^ t29479;
    wire t29481 = t29480 ^ t29480;
    wire t29482 = t29481 ^ t29481;
    wire t29483 = t29482 ^ t29482;
    wire t29484 = t29483 ^ t29483;
    wire t29485 = t29484 ^ t29484;
    wire t29486 = t29485 ^ t29485;
    wire t29487 = t29486 ^ t29486;
    wire t29488 = t29487 ^ t29487;
    wire t29489 = t29488 ^ t29488;
    wire t29490 = t29489 ^ t29489;
    wire t29491 = t29490 ^ t29490;
    wire t29492 = t29491 ^ t29491;
    wire t29493 = t29492 ^ t29492;
    wire t29494 = t29493 ^ t29493;
    wire t29495 = t29494 ^ t29494;
    wire t29496 = t29495 ^ t29495;
    wire t29497 = t29496 ^ t29496;
    wire t29498 = t29497 ^ t29497;
    wire t29499 = t29498 ^ t29498;
    wire t29500 = t29499 ^ t29499;
    wire t29501 = t29500 ^ t29500;
    wire t29502 = t29501 ^ t29501;
    wire t29503 = t29502 ^ t29502;
    wire t29504 = t29503 ^ t29503;
    wire t29505 = t29504 ^ t29504;
    wire t29506 = t29505 ^ t29505;
    wire t29507 = t29506 ^ t29506;
    wire t29508 = t29507 ^ t29507;
    wire t29509 = t29508 ^ t29508;
    wire t29510 = t29509 ^ t29509;
    wire t29511 = t29510 ^ t29510;
    wire t29512 = t29511 ^ t29511;
    wire t29513 = t29512 ^ t29512;
    wire t29514 = t29513 ^ t29513;
    wire t29515 = t29514 ^ t29514;
    wire t29516 = t29515 ^ t29515;
    wire t29517 = t29516 ^ t29516;
    wire t29518 = t29517 ^ t29517;
    wire t29519 = t29518 ^ t29518;
    wire t29520 = t29519 ^ t29519;
    wire t29521 = t29520 ^ t29520;
    wire t29522 = t29521 ^ t29521;
    wire t29523 = t29522 ^ t29522;
    wire t29524 = t29523 ^ t29523;
    wire t29525 = t29524 ^ t29524;
    wire t29526 = t29525 ^ t29525;
    wire t29527 = t29526 ^ t29526;
    wire t29528 = t29527 ^ t29527;
    wire t29529 = t29528 ^ t29528;
    wire t29530 = t29529 ^ t29529;
    wire t29531 = t29530 ^ t29530;
    wire t29532 = t29531 ^ t29531;
    wire t29533 = t29532 ^ t29532;
    wire t29534 = t29533 ^ t29533;
    wire t29535 = t29534 ^ t29534;
    wire t29536 = t29535 ^ t29535;
    wire t29537 = t29536 ^ t29536;
    wire t29538 = t29537 ^ t29537;
    wire t29539 = t29538 ^ t29538;
    wire t29540 = t29539 ^ t29539;
    wire t29541 = t29540 ^ t29540;
    wire t29542 = t29541 ^ t29541;
    wire t29543 = t29542 ^ t29542;
    wire t29544 = t29543 ^ t29543;
    wire t29545 = t29544 ^ t29544;
    wire t29546 = t29545 ^ t29545;
    wire t29547 = t29546 ^ t29546;
    wire t29548 = t29547 ^ t29547;
    wire t29549 = t29548 ^ t29548;
    wire t29550 = t29549 ^ t29549;
    wire t29551 = t29550 ^ t29550;
    wire t29552 = t29551 ^ t29551;
    wire t29553 = t29552 ^ t29552;
    wire t29554 = t29553 ^ t29553;
    wire t29555 = t29554 ^ t29554;
    wire t29556 = t29555 ^ t29555;
    wire t29557 = t29556 ^ t29556;
    wire t29558 = t29557 ^ t29557;
    wire t29559 = t29558 ^ t29558;
    wire t29560 = t29559 ^ t29559;
    wire t29561 = t29560 ^ t29560;
    wire t29562 = t29561 ^ t29561;
    wire t29563 = t29562 ^ t29562;
    wire t29564 = t29563 ^ t29563;
    wire t29565 = t29564 ^ t29564;
    wire t29566 = t29565 ^ t29565;
    wire t29567 = t29566 ^ t29566;
    wire t29568 = t29567 ^ t29567;
    wire t29569 = t29568 ^ t29568;
    wire t29570 = t29569 ^ t29569;
    wire t29571 = t29570 ^ t29570;
    wire t29572 = t29571 ^ t29571;
    wire t29573 = t29572 ^ t29572;
    wire t29574 = t29573 ^ t29573;
    wire t29575 = t29574 ^ t29574;
    wire t29576 = t29575 ^ t29575;
    wire t29577 = t29576 ^ t29576;
    wire t29578 = t29577 ^ t29577;
    wire t29579 = t29578 ^ t29578;
    wire t29580 = t29579 ^ t29579;
    wire t29581 = t29580 ^ t29580;
    wire t29582 = t29581 ^ t29581;
    wire t29583 = t29582 ^ t29582;
    wire t29584 = t29583 ^ t29583;
    wire t29585 = t29584 ^ t29584;
    wire t29586 = t29585 ^ t29585;
    wire t29587 = t29586 ^ t29586;
    wire t29588 = t29587 ^ t29587;
    wire t29589 = t29588 ^ t29588;
    wire t29590 = t29589 ^ t29589;
    wire t29591 = t29590 ^ t29590;
    wire t29592 = t29591 ^ t29591;
    wire t29593 = t29592 ^ t29592;
    wire t29594 = t29593 ^ t29593;
    wire t29595 = t29594 ^ t29594;
    wire t29596 = t29595 ^ t29595;
    wire t29597 = t29596 ^ t29596;
    wire t29598 = t29597 ^ t29597;
    wire t29599 = t29598 ^ t29598;
    wire t29600 = t29599 ^ t29599;
    wire t29601 = t29600 ^ t29600;
    wire t29602 = t29601 ^ t29601;
    wire t29603 = t29602 ^ t29602;
    wire t29604 = t29603 ^ t29603;
    wire t29605 = t29604 ^ t29604;
    wire t29606 = t29605 ^ t29605;
    wire t29607 = t29606 ^ t29606;
    wire t29608 = t29607 ^ t29607;
    wire t29609 = t29608 ^ t29608;
    wire t29610 = t29609 ^ t29609;
    wire t29611 = t29610 ^ t29610;
    wire t29612 = t29611 ^ t29611;
    wire t29613 = t29612 ^ t29612;
    wire t29614 = t29613 ^ t29613;
    wire t29615 = t29614 ^ t29614;
    wire t29616 = t29615 ^ t29615;
    wire t29617 = t29616 ^ t29616;
    wire t29618 = t29617 ^ t29617;
    wire t29619 = t29618 ^ t29618;
    wire t29620 = t29619 ^ t29619;
    wire t29621 = t29620 ^ t29620;
    wire t29622 = t29621 ^ t29621;
    wire t29623 = t29622 ^ t29622;
    wire t29624 = t29623 ^ t29623;
    wire t29625 = t29624 ^ t29624;
    wire t29626 = t29625 ^ t29625;
    wire t29627 = t29626 ^ t29626;
    wire t29628 = t29627 ^ t29627;
    wire t29629 = t29628 ^ t29628;
    wire t29630 = t29629 ^ t29629;
    wire t29631 = t29630 ^ t29630;
    wire t29632 = t29631 ^ t29631;
    wire t29633 = t29632 ^ t29632;
    wire t29634 = t29633 ^ t29633;
    wire t29635 = t29634 ^ t29634;
    wire t29636 = t29635 ^ t29635;
    wire t29637 = t29636 ^ t29636;
    wire t29638 = t29637 ^ t29637;
    wire t29639 = t29638 ^ t29638;
    wire t29640 = t29639 ^ t29639;
    wire t29641 = t29640 ^ t29640;
    wire t29642 = t29641 ^ t29641;
    wire t29643 = t29642 ^ t29642;
    wire t29644 = t29643 ^ t29643;
    wire t29645 = t29644 ^ t29644;
    wire t29646 = t29645 ^ t29645;
    wire t29647 = t29646 ^ t29646;
    wire t29648 = t29647 ^ t29647;
    wire t29649 = t29648 ^ t29648;
    wire t29650 = t29649 ^ t29649;
    wire t29651 = t29650 ^ t29650;
    wire t29652 = t29651 ^ t29651;
    wire t29653 = t29652 ^ t29652;
    wire t29654 = t29653 ^ t29653;
    wire t29655 = t29654 ^ t29654;
    wire t29656 = t29655 ^ t29655;
    wire t29657 = t29656 ^ t29656;
    wire t29658 = t29657 ^ t29657;
    wire t29659 = t29658 ^ t29658;
    wire t29660 = t29659 ^ t29659;
    wire t29661 = t29660 ^ t29660;
    wire t29662 = t29661 ^ t29661;
    wire t29663 = t29662 ^ t29662;
    wire t29664 = t29663 ^ t29663;
    wire t29665 = t29664 ^ t29664;
    wire t29666 = t29665 ^ t29665;
    wire t29667 = t29666 ^ t29666;
    wire t29668 = t29667 ^ t29667;
    wire t29669 = t29668 ^ t29668;
    wire t29670 = t29669 ^ t29669;
    wire t29671 = t29670 ^ t29670;
    wire t29672 = t29671 ^ t29671;
    wire t29673 = t29672 ^ t29672;
    wire t29674 = t29673 ^ t29673;
    wire t29675 = t29674 ^ t29674;
    wire t29676 = t29675 ^ t29675;
    wire t29677 = t29676 ^ t29676;
    wire t29678 = t29677 ^ t29677;
    wire t29679 = t29678 ^ t29678;
    wire t29680 = t29679 ^ t29679;
    wire t29681 = t29680 ^ t29680;
    wire t29682 = t29681 ^ t29681;
    wire t29683 = t29682 ^ t29682;
    wire t29684 = t29683 ^ t29683;
    wire t29685 = t29684 ^ t29684;
    wire t29686 = t29685 ^ t29685;
    wire t29687 = t29686 ^ t29686;
    wire t29688 = t29687 ^ t29687;
    wire t29689 = t29688 ^ t29688;
    wire t29690 = t29689 ^ t29689;
    wire t29691 = t29690 ^ t29690;
    wire t29692 = t29691 ^ t29691;
    wire t29693 = t29692 ^ t29692;
    wire t29694 = t29693 ^ t29693;
    wire t29695 = t29694 ^ t29694;
    wire t29696 = t29695 ^ t29695;
    wire t29697 = t29696 ^ t29696;
    wire t29698 = t29697 ^ t29697;
    wire t29699 = t29698 ^ t29698;
    wire t29700 = t29699 ^ t29699;
    wire t29701 = t29700 ^ t29700;
    wire t29702 = t29701 ^ t29701;
    wire t29703 = t29702 ^ t29702;
    wire t29704 = t29703 ^ t29703;
    wire t29705 = t29704 ^ t29704;
    wire t29706 = t29705 ^ t29705;
    wire t29707 = t29706 ^ t29706;
    wire t29708 = t29707 ^ t29707;
    wire t29709 = t29708 ^ t29708;
    wire t29710 = t29709 ^ t29709;
    wire t29711 = t29710 ^ t29710;
    wire t29712 = t29711 ^ t29711;
    wire t29713 = t29712 ^ t29712;
    wire t29714 = t29713 ^ t29713;
    wire t29715 = t29714 ^ t29714;
    wire t29716 = t29715 ^ t29715;
    wire t29717 = t29716 ^ t29716;
    wire t29718 = t29717 ^ t29717;
    wire t29719 = t29718 ^ t29718;
    wire t29720 = t29719 ^ t29719;
    wire t29721 = t29720 ^ t29720;
    wire t29722 = t29721 ^ t29721;
    wire t29723 = t29722 ^ t29722;
    wire t29724 = t29723 ^ t29723;
    wire t29725 = t29724 ^ t29724;
    wire t29726 = t29725 ^ t29725;
    wire t29727 = t29726 ^ t29726;
    wire t29728 = t29727 ^ t29727;
    wire t29729 = t29728 ^ t29728;
    wire t29730 = t29729 ^ t29729;
    wire t29731 = t29730 ^ t29730;
    wire t29732 = t29731 ^ t29731;
    wire t29733 = t29732 ^ t29732;
    wire t29734 = t29733 ^ t29733;
    wire t29735 = t29734 ^ t29734;
    wire t29736 = t29735 ^ t29735;
    wire t29737 = t29736 ^ t29736;
    wire t29738 = t29737 ^ t29737;
    wire t29739 = t29738 ^ t29738;
    wire t29740 = t29739 ^ t29739;
    wire t29741 = t29740 ^ t29740;
    wire t29742 = t29741 ^ t29741;
    wire t29743 = t29742 ^ t29742;
    wire t29744 = t29743 ^ t29743;
    wire t29745 = t29744 ^ t29744;
    wire t29746 = t29745 ^ t29745;
    wire t29747 = t29746 ^ t29746;
    wire t29748 = t29747 ^ t29747;
    wire t29749 = t29748 ^ t29748;
    wire t29750 = t29749 ^ t29749;
    wire t29751 = t29750 ^ t29750;
    wire t29752 = t29751 ^ t29751;
    wire t29753 = t29752 ^ t29752;
    wire t29754 = t29753 ^ t29753;
    wire t29755 = t29754 ^ t29754;
    wire t29756 = t29755 ^ t29755;
    wire t29757 = t29756 ^ t29756;
    wire t29758 = t29757 ^ t29757;
    wire t29759 = t29758 ^ t29758;
    wire t29760 = t29759 ^ t29759;
    wire t29761 = t29760 ^ t29760;
    wire t29762 = t29761 ^ t29761;
    wire t29763 = t29762 ^ t29762;
    wire t29764 = t29763 ^ t29763;
    wire t29765 = t29764 ^ t29764;
    wire t29766 = t29765 ^ t29765;
    wire t29767 = t29766 ^ t29766;
    wire t29768 = t29767 ^ t29767;
    wire t29769 = t29768 ^ t29768;
    wire t29770 = t29769 ^ t29769;
    wire t29771 = t29770 ^ t29770;
    wire t29772 = t29771 ^ t29771;
    wire t29773 = t29772 ^ t29772;
    wire t29774 = t29773 ^ t29773;
    wire t29775 = t29774 ^ t29774;
    wire t29776 = t29775 ^ t29775;
    wire t29777 = t29776 ^ t29776;
    wire t29778 = t29777 ^ t29777;
    wire t29779 = t29778 ^ t29778;
    wire t29780 = t29779 ^ t29779;
    wire t29781 = t29780 ^ t29780;
    wire t29782 = t29781 ^ t29781;
    wire t29783 = t29782 ^ t29782;
    wire t29784 = t29783 ^ t29783;
    wire t29785 = t29784 ^ t29784;
    wire t29786 = t29785 ^ t29785;
    wire t29787 = t29786 ^ t29786;
    wire t29788 = t29787 ^ t29787;
    wire t29789 = t29788 ^ t29788;
    wire t29790 = t29789 ^ t29789;
    wire t29791 = t29790 ^ t29790;
    wire t29792 = t29791 ^ t29791;
    wire t29793 = t29792 ^ t29792;
    wire t29794 = t29793 ^ t29793;
    wire t29795 = t29794 ^ t29794;
    wire t29796 = t29795 ^ t29795;
    wire t29797 = t29796 ^ t29796;
    wire t29798 = t29797 ^ t29797;
    wire t29799 = t29798 ^ t29798;
    wire t29800 = t29799 ^ t29799;
    wire t29801 = t29800 ^ t29800;
    wire t29802 = t29801 ^ t29801;
    wire t29803 = t29802 ^ t29802;
    wire t29804 = t29803 ^ t29803;
    wire t29805 = t29804 ^ t29804;
    wire t29806 = t29805 ^ t29805;
    wire t29807 = t29806 ^ t29806;
    wire t29808 = t29807 ^ t29807;
    wire t29809 = t29808 ^ t29808;
    wire t29810 = t29809 ^ t29809;
    wire t29811 = t29810 ^ t29810;
    wire t29812 = t29811 ^ t29811;
    wire t29813 = t29812 ^ t29812;
    wire t29814 = t29813 ^ t29813;
    wire t29815 = t29814 ^ t29814;
    wire t29816 = t29815 ^ t29815;
    wire t29817 = t29816 ^ t29816;
    wire t29818 = t29817 ^ t29817;
    wire t29819 = t29818 ^ t29818;
    wire t29820 = t29819 ^ t29819;
    wire t29821 = t29820 ^ t29820;
    wire t29822 = t29821 ^ t29821;
    wire t29823 = t29822 ^ t29822;
    wire t29824 = t29823 ^ t29823;
    wire t29825 = t29824 ^ t29824;
    wire t29826 = t29825 ^ t29825;
    wire t29827 = t29826 ^ t29826;
    wire t29828 = t29827 ^ t29827;
    wire t29829 = t29828 ^ t29828;
    wire t29830 = t29829 ^ t29829;
    wire t29831 = t29830 ^ t29830;
    wire t29832 = t29831 ^ t29831;
    wire t29833 = t29832 ^ t29832;
    wire t29834 = t29833 ^ t29833;
    wire t29835 = t29834 ^ t29834;
    wire t29836 = t29835 ^ t29835;
    wire t29837 = t29836 ^ t29836;
    wire t29838 = t29837 ^ t29837;
    wire t29839 = t29838 ^ t29838;
    wire t29840 = t29839 ^ t29839;
    wire t29841 = t29840 ^ t29840;
    wire t29842 = t29841 ^ t29841;
    wire t29843 = t29842 ^ t29842;
    wire t29844 = t29843 ^ t29843;
    wire t29845 = t29844 ^ t29844;
    wire t29846 = t29845 ^ t29845;
    wire t29847 = t29846 ^ t29846;
    wire t29848 = t29847 ^ t29847;
    wire t29849 = t29848 ^ t29848;
    wire t29850 = t29849 ^ t29849;
    wire t29851 = t29850 ^ t29850;
    wire t29852 = t29851 ^ t29851;
    wire t29853 = t29852 ^ t29852;
    wire t29854 = t29853 ^ t29853;
    wire t29855 = t29854 ^ t29854;
    wire t29856 = t29855 ^ t29855;
    wire t29857 = t29856 ^ t29856;
    wire t29858 = t29857 ^ t29857;
    wire t29859 = t29858 ^ t29858;
    wire t29860 = t29859 ^ t29859;
    wire t29861 = t29860 ^ t29860;
    wire t29862 = t29861 ^ t29861;
    wire t29863 = t29862 ^ t29862;
    wire t29864 = t29863 ^ t29863;
    wire t29865 = t29864 ^ t29864;
    wire t29866 = t29865 ^ t29865;
    wire t29867 = t29866 ^ t29866;
    wire t29868 = t29867 ^ t29867;
    wire t29869 = t29868 ^ t29868;
    wire t29870 = t29869 ^ t29869;
    wire t29871 = t29870 ^ t29870;
    wire t29872 = t29871 ^ t29871;
    wire t29873 = t29872 ^ t29872;
    wire t29874 = t29873 ^ t29873;
    wire t29875 = t29874 ^ t29874;
    wire t29876 = t29875 ^ t29875;
    wire t29877 = t29876 ^ t29876;
    wire t29878 = t29877 ^ t29877;
    wire t29879 = t29878 ^ t29878;
    wire t29880 = t29879 ^ t29879;
    wire t29881 = t29880 ^ t29880;
    wire t29882 = t29881 ^ t29881;
    wire t29883 = t29882 ^ t29882;
    wire t29884 = t29883 ^ t29883;
    wire t29885 = t29884 ^ t29884;
    wire t29886 = t29885 ^ t29885;
    wire t29887 = t29886 ^ t29886;
    wire t29888 = t29887 ^ t29887;
    wire t29889 = t29888 ^ t29888;
    wire t29890 = t29889 ^ t29889;
    wire t29891 = t29890 ^ t29890;
    wire t29892 = t29891 ^ t29891;
    wire t29893 = t29892 ^ t29892;
    wire t29894 = t29893 ^ t29893;
    wire t29895 = t29894 ^ t29894;
    wire t29896 = t29895 ^ t29895;
    wire t29897 = t29896 ^ t29896;
    wire t29898 = t29897 ^ t29897;
    wire t29899 = t29898 ^ t29898;
    wire t29900 = t29899 ^ t29899;
    wire t29901 = t29900 ^ t29900;
    wire t29902 = t29901 ^ t29901;
    wire t29903 = t29902 ^ t29902;
    wire t29904 = t29903 ^ t29903;
    wire t29905 = t29904 ^ t29904;
    wire t29906 = t29905 ^ t29905;
    wire t29907 = t29906 ^ t29906;
    wire t29908 = t29907 ^ t29907;
    wire t29909 = t29908 ^ t29908;
    wire t29910 = t29909 ^ t29909;
    wire t29911 = t29910 ^ t29910;
    wire t29912 = t29911 ^ t29911;
    wire t29913 = t29912 ^ t29912;
    wire t29914 = t29913 ^ t29913;
    wire t29915 = t29914 ^ t29914;
    wire t29916 = t29915 ^ t29915;
    wire t29917 = t29916 ^ t29916;
    wire t29918 = t29917 ^ t29917;
    wire t29919 = t29918 ^ t29918;
    wire t29920 = t29919 ^ t29919;
    wire t29921 = t29920 ^ t29920;
    wire t29922 = t29921 ^ t29921;
    wire t29923 = t29922 ^ t29922;
    wire t29924 = t29923 ^ t29923;
    wire t29925 = t29924 ^ t29924;
    wire t29926 = t29925 ^ t29925;
    wire t29927 = t29926 ^ t29926;
    wire t29928 = t29927 ^ t29927;
    wire t29929 = t29928 ^ t29928;
    wire t29930 = t29929 ^ t29929;
    wire t29931 = t29930 ^ t29930;
    wire t29932 = t29931 ^ t29931;
    wire t29933 = t29932 ^ t29932;
    wire t29934 = t29933 ^ t29933;
    wire t29935 = t29934 ^ t29934;
    wire t29936 = t29935 ^ t29935;
    wire t29937 = t29936 ^ t29936;
    wire t29938 = t29937 ^ t29937;
    wire t29939 = t29938 ^ t29938;
    wire t29940 = t29939 ^ t29939;
    wire t29941 = t29940 ^ t29940;
    wire t29942 = t29941 ^ t29941;
    wire t29943 = t29942 ^ t29942;
    wire t29944 = t29943 ^ t29943;
    wire t29945 = t29944 ^ t29944;
    wire t29946 = t29945 ^ t29945;
    wire t29947 = t29946 ^ t29946;
    wire t29948 = t29947 ^ t29947;
    wire t29949 = t29948 ^ t29948;
    wire t29950 = t29949 ^ t29949;
    wire t29951 = t29950 ^ t29950;
    wire t29952 = t29951 ^ t29951;
    wire t29953 = t29952 ^ t29952;
    wire t29954 = t29953 ^ t29953;
    wire t29955 = t29954 ^ t29954;
    wire t29956 = t29955 ^ t29955;
    wire t29957 = t29956 ^ t29956;
    wire t29958 = t29957 ^ t29957;
    wire t29959 = t29958 ^ t29958;
    wire t29960 = t29959 ^ t29959;
    wire t29961 = t29960 ^ t29960;
    wire t29962 = t29961 ^ t29961;
    wire t29963 = t29962 ^ t29962;
    wire t29964 = t29963 ^ t29963;
    wire t29965 = t29964 ^ t29964;
    wire t29966 = t29965 ^ t29965;
    wire t29967 = t29966 ^ t29966;
    wire t29968 = t29967 ^ t29967;
    wire t29969 = t29968 ^ t29968;
    wire t29970 = t29969 ^ t29969;
    wire t29971 = t29970 ^ t29970;
    wire t29972 = t29971 ^ t29971;
    wire t29973 = t29972 ^ t29972;
    wire t29974 = t29973 ^ t29973;
    wire t29975 = t29974 ^ t29974;
    wire t29976 = t29975 ^ t29975;
    wire t29977 = t29976 ^ t29976;
    wire t29978 = t29977 ^ t29977;
    wire t29979 = t29978 ^ t29978;
    wire t29980 = t29979 ^ t29979;
    wire t29981 = t29980 ^ t29980;
    wire t29982 = t29981 ^ t29981;
    wire t29983 = t29982 ^ t29982;
    wire t29984 = t29983 ^ t29983;
    wire t29985 = t29984 ^ t29984;
    wire t29986 = t29985 ^ t29985;
    wire t29987 = t29986 ^ t29986;
    wire t29988 = t29987 ^ t29987;
    wire t29989 = t29988 ^ t29988;
    wire t29990 = t29989 ^ t29989;
    wire t29991 = t29990 ^ t29990;
    wire t29992 = t29991 ^ t29991;
    wire t29993 = t29992 ^ t29992;
    wire t29994 = t29993 ^ t29993;
    wire t29995 = t29994 ^ t29994;
    wire t29996 = t29995 ^ t29995;
    wire t29997 = t29996 ^ t29996;
    wire t29998 = t29997 ^ t29997;
    wire t29999 = t29998 ^ t29998;
    wire t30000 = t29999 ^ t29999;
    wire t30001 = t30000 ^ t30000;
    wire t30002 = t30001 ^ t30001;
    wire t30003 = t30002 ^ t30002;
    wire t30004 = t30003 ^ t30003;
    wire t30005 = t30004 ^ t30004;
    wire t30006 = t30005 ^ t30005;
    wire t30007 = t30006 ^ t30006;
    wire t30008 = t30007 ^ t30007;
    wire t30009 = t30008 ^ t30008;
    wire t30010 = t30009 ^ t30009;
    wire t30011 = t30010 ^ t30010;
    wire t30012 = t30011 ^ t30011;
    wire t30013 = t30012 ^ t30012;
    wire t30014 = t30013 ^ t30013;
    wire t30015 = t30014 ^ t30014;
    wire t30016 = t30015 ^ t30015;
    wire t30017 = t30016 ^ t30016;
    wire t30018 = t30017 ^ t30017;
    wire t30019 = t30018 ^ t30018;
    wire t30020 = t30019 ^ t30019;
    wire t30021 = t30020 ^ t30020;
    wire t30022 = t30021 ^ t30021;
    wire t30023 = t30022 ^ t30022;
    wire t30024 = t30023 ^ t30023;
    wire t30025 = t30024 ^ t30024;
    wire t30026 = t30025 ^ t30025;
    wire t30027 = t30026 ^ t30026;
    wire t30028 = t30027 ^ t30027;
    wire t30029 = t30028 ^ t30028;
    wire t30030 = t30029 ^ t30029;
    wire t30031 = t30030 ^ t30030;
    wire t30032 = t30031 ^ t30031;
    wire t30033 = t30032 ^ t30032;
    wire t30034 = t30033 ^ t30033;
    wire t30035 = t30034 ^ t30034;
    wire t30036 = t30035 ^ t30035;
    wire t30037 = t30036 ^ t30036;
    wire t30038 = t30037 ^ t30037;
    wire t30039 = t30038 ^ t30038;
    wire t30040 = t30039 ^ t30039;
    wire t30041 = t30040 ^ t30040;
    wire t30042 = t30041 ^ t30041;
    wire t30043 = t30042 ^ t30042;
    wire t30044 = t30043 ^ t30043;
    wire t30045 = t30044 ^ t30044;
    wire t30046 = t30045 ^ t30045;
    wire t30047 = t30046 ^ t30046;
    wire t30048 = t30047 ^ t30047;
    wire t30049 = t30048 ^ t30048;
    wire t30050 = t30049 ^ t30049;
    wire t30051 = t30050 ^ t30050;
    wire t30052 = t30051 ^ t30051;
    wire t30053 = t30052 ^ t30052;
    wire t30054 = t30053 ^ t30053;
    wire t30055 = t30054 ^ t30054;
    wire t30056 = t30055 ^ t30055;
    wire t30057 = t30056 ^ t30056;
    wire t30058 = t30057 ^ t30057;
    wire t30059 = t30058 ^ t30058;
    wire t30060 = t30059 ^ t30059;
    wire t30061 = t30060 ^ t30060;
    wire t30062 = t30061 ^ t30061;
    wire t30063 = t30062 ^ t30062;
    wire t30064 = t30063 ^ t30063;
    wire t30065 = t30064 ^ t30064;
    wire t30066 = t30065 ^ t30065;
    wire t30067 = t30066 ^ t30066;
    wire t30068 = t30067 ^ t30067;
    wire t30069 = t30068 ^ t30068;
    wire t30070 = t30069 ^ t30069;
    wire t30071 = t30070 ^ t30070;
    wire t30072 = t30071 ^ t30071;
    wire t30073 = t30072 ^ t30072;
    wire t30074 = t30073 ^ t30073;
    wire t30075 = t30074 ^ t30074;
    wire t30076 = t30075 ^ t30075;
    wire t30077 = t30076 ^ t30076;
    wire t30078 = t30077 ^ t30077;
    wire t30079 = t30078 ^ t30078;
    wire t30080 = t30079 ^ t30079;
    wire t30081 = t30080 ^ t30080;
    wire t30082 = t30081 ^ t30081;
    wire t30083 = t30082 ^ t30082;
    wire t30084 = t30083 ^ t30083;
    wire t30085 = t30084 ^ t30084;
    wire t30086 = t30085 ^ t30085;
    wire t30087 = t30086 ^ t30086;
    wire t30088 = t30087 ^ t30087;
    wire t30089 = t30088 ^ t30088;
    wire t30090 = t30089 ^ t30089;
    wire t30091 = t30090 ^ t30090;
    wire t30092 = t30091 ^ t30091;
    wire t30093 = t30092 ^ t30092;
    wire t30094 = t30093 ^ t30093;
    wire t30095 = t30094 ^ t30094;
    wire t30096 = t30095 ^ t30095;
    wire t30097 = t30096 ^ t30096;
    wire t30098 = t30097 ^ t30097;
    wire t30099 = t30098 ^ t30098;
    wire t30100 = t30099 ^ t30099;
    wire t30101 = t30100 ^ t30100;
    wire t30102 = t30101 ^ t30101;
    wire t30103 = t30102 ^ t30102;
    wire t30104 = t30103 ^ t30103;
    wire t30105 = t30104 ^ t30104;
    wire t30106 = t30105 ^ t30105;
    wire t30107 = t30106 ^ t30106;
    wire t30108 = t30107 ^ t30107;
    wire t30109 = t30108 ^ t30108;
    wire t30110 = t30109 ^ t30109;
    wire t30111 = t30110 ^ t30110;
    wire t30112 = t30111 ^ t30111;
    wire t30113 = t30112 ^ t30112;
    wire t30114 = t30113 ^ t30113;
    wire t30115 = t30114 ^ t30114;
    wire t30116 = t30115 ^ t30115;
    wire t30117 = t30116 ^ t30116;
    wire t30118 = t30117 ^ t30117;
    wire t30119 = t30118 ^ t30118;
    wire t30120 = t30119 ^ t30119;
    wire t30121 = t30120 ^ t30120;
    wire t30122 = t30121 ^ t30121;
    wire t30123 = t30122 ^ t30122;
    wire t30124 = t30123 ^ t30123;
    wire t30125 = t30124 ^ t30124;
    wire t30126 = t30125 ^ t30125;
    wire t30127 = t30126 ^ t30126;
    wire t30128 = t30127 ^ t30127;
    wire t30129 = t30128 ^ t30128;
    wire t30130 = t30129 ^ t30129;
    wire t30131 = t30130 ^ t30130;
    wire t30132 = t30131 ^ t30131;
    wire t30133 = t30132 ^ t30132;
    wire t30134 = t30133 ^ t30133;
    wire t30135 = t30134 ^ t30134;
    wire t30136 = t30135 ^ t30135;
    wire t30137 = t30136 ^ t30136;
    wire t30138 = t30137 ^ t30137;
    wire t30139 = t30138 ^ t30138;
    wire t30140 = t30139 ^ t30139;
    wire t30141 = t30140 ^ t30140;
    wire t30142 = t30141 ^ t30141;
    wire t30143 = t30142 ^ t30142;
    wire t30144 = t30143 ^ t30143;
    wire t30145 = t30144 ^ t30144;
    wire t30146 = t30145 ^ t30145;
    wire t30147 = t30146 ^ t30146;
    wire t30148 = t30147 ^ t30147;
    wire t30149 = t30148 ^ t30148;
    wire t30150 = t30149 ^ t30149;
    wire t30151 = t30150 ^ t30150;
    wire t30152 = t30151 ^ t30151;
    wire t30153 = t30152 ^ t30152;
    wire t30154 = t30153 ^ t30153;
    wire t30155 = t30154 ^ t30154;
    wire t30156 = t30155 ^ t30155;
    wire t30157 = t30156 ^ t30156;
    wire t30158 = t30157 ^ t30157;
    wire t30159 = t30158 ^ t30158;
    wire t30160 = t30159 ^ t30159;
    wire t30161 = t30160 ^ t30160;
    wire t30162 = t30161 ^ t30161;
    wire t30163 = t30162 ^ t30162;
    wire t30164 = t30163 ^ t30163;
    wire t30165 = t30164 ^ t30164;
    wire t30166 = t30165 ^ t30165;
    wire t30167 = t30166 ^ t30166;
    wire t30168 = t30167 ^ t30167;
    wire t30169 = t30168 ^ t30168;
    wire t30170 = t30169 ^ t30169;
    wire t30171 = t30170 ^ t30170;
    wire t30172 = t30171 ^ t30171;
    wire t30173 = t30172 ^ t30172;
    wire t30174 = t30173 ^ t30173;
    wire t30175 = t30174 ^ t30174;
    wire t30176 = t30175 ^ t30175;
    wire t30177 = t30176 ^ t30176;
    wire t30178 = t30177 ^ t30177;
    wire t30179 = t30178 ^ t30178;
    wire t30180 = t30179 ^ t30179;
    wire t30181 = t30180 ^ t30180;
    wire t30182 = t30181 ^ t30181;
    wire t30183 = t30182 ^ t30182;
    wire t30184 = t30183 ^ t30183;
    wire t30185 = t30184 ^ t30184;
    wire t30186 = t30185 ^ t30185;
    wire t30187 = t30186 ^ t30186;
    wire t30188 = t30187 ^ t30187;
    wire t30189 = t30188 ^ t30188;
    wire t30190 = t30189 ^ t30189;
    wire t30191 = t30190 ^ t30190;
    wire t30192 = t30191 ^ t30191;
    wire t30193 = t30192 ^ t30192;
    wire t30194 = t30193 ^ t30193;
    wire t30195 = t30194 ^ t30194;
    wire t30196 = t30195 ^ t30195;
    wire t30197 = t30196 ^ t30196;
    wire t30198 = t30197 ^ t30197;
    wire t30199 = t30198 ^ t30198;
    wire t30200 = t30199 ^ t30199;
    wire t30201 = t30200 ^ t30200;
    wire t30202 = t30201 ^ t30201;
    wire t30203 = t30202 ^ t30202;
    wire t30204 = t30203 ^ t30203;
    wire t30205 = t30204 ^ t30204;
    wire t30206 = t30205 ^ t30205;
    wire t30207 = t30206 ^ t30206;
    wire t30208 = t30207 ^ t30207;
    wire t30209 = t30208 ^ t30208;
    wire t30210 = t30209 ^ t30209;
    wire t30211 = t30210 ^ t30210;
    wire t30212 = t30211 ^ t30211;
    wire t30213 = t30212 ^ t30212;
    wire t30214 = t30213 ^ t30213;
    wire t30215 = t30214 ^ t30214;
    wire t30216 = t30215 ^ t30215;
    wire t30217 = t30216 ^ t30216;
    wire t30218 = t30217 ^ t30217;
    wire t30219 = t30218 ^ t30218;
    wire t30220 = t30219 ^ t30219;
    wire t30221 = t30220 ^ t30220;
    wire t30222 = t30221 ^ t30221;
    wire t30223 = t30222 ^ t30222;
    wire t30224 = t30223 ^ t30223;
    wire t30225 = t30224 ^ t30224;
    wire t30226 = t30225 ^ t30225;
    wire t30227 = t30226 ^ t30226;
    wire t30228 = t30227 ^ t30227;
    wire t30229 = t30228 ^ t30228;
    wire t30230 = t30229 ^ t30229;
    wire t30231 = t30230 ^ t30230;
    wire t30232 = t30231 ^ t30231;
    wire t30233 = t30232 ^ t30232;
    wire t30234 = t30233 ^ t30233;
    wire t30235 = t30234 ^ t30234;
    wire t30236 = t30235 ^ t30235;
    wire t30237 = t30236 ^ t30236;
    wire t30238 = t30237 ^ t30237;
    wire t30239 = t30238 ^ t30238;
    wire t30240 = t30239 ^ t30239;
    wire t30241 = t30240 ^ t30240;
    wire t30242 = t30241 ^ t30241;
    wire t30243 = t30242 ^ t30242;
    wire t30244 = t30243 ^ t30243;
    wire t30245 = t30244 ^ t30244;
    wire t30246 = t30245 ^ t30245;
    wire t30247 = t30246 ^ t30246;
    wire t30248 = t30247 ^ t30247;
    wire t30249 = t30248 ^ t30248;
    wire t30250 = t30249 ^ t30249;
    wire t30251 = t30250 ^ t30250;
    wire t30252 = t30251 ^ t30251;
    wire t30253 = t30252 ^ t30252;
    wire t30254 = t30253 ^ t30253;
    wire t30255 = t30254 ^ t30254;
    wire t30256 = t30255 ^ t30255;
    wire t30257 = t30256 ^ t30256;
    wire t30258 = t30257 ^ t30257;
    wire t30259 = t30258 ^ t30258;
    wire t30260 = t30259 ^ t30259;
    wire t30261 = t30260 ^ t30260;
    wire t30262 = t30261 ^ t30261;
    wire t30263 = t30262 ^ t30262;
    wire t30264 = t30263 ^ t30263;
    wire t30265 = t30264 ^ t30264;
    wire t30266 = t30265 ^ t30265;
    wire t30267 = t30266 ^ t30266;
    wire t30268 = t30267 ^ t30267;
    wire t30269 = t30268 ^ t30268;
    wire t30270 = t30269 ^ t30269;
    wire t30271 = t30270 ^ t30270;
    wire t30272 = t30271 ^ t30271;
    wire t30273 = t30272 ^ t30272;
    wire t30274 = t30273 ^ t30273;
    wire t30275 = t30274 ^ t30274;
    wire t30276 = t30275 ^ t30275;
    wire t30277 = t30276 ^ t30276;
    wire t30278 = t30277 ^ t30277;
    wire t30279 = t30278 ^ t30278;
    wire t30280 = t30279 ^ t30279;
    wire t30281 = t30280 ^ t30280;
    wire t30282 = t30281 ^ t30281;
    wire t30283 = t30282 ^ t30282;
    wire t30284 = t30283 ^ t30283;
    wire t30285 = t30284 ^ t30284;
    wire t30286 = t30285 ^ t30285;
    wire t30287 = t30286 ^ t30286;
    wire t30288 = t30287 ^ t30287;
    wire t30289 = t30288 ^ t30288;
    wire t30290 = t30289 ^ t30289;
    wire t30291 = t30290 ^ t30290;
    wire t30292 = t30291 ^ t30291;
    wire t30293 = t30292 ^ t30292;
    wire t30294 = t30293 ^ t30293;
    wire t30295 = t30294 ^ t30294;
    wire t30296 = t30295 ^ t30295;
    wire t30297 = t30296 ^ t30296;
    wire t30298 = t30297 ^ t30297;
    wire t30299 = t30298 ^ t30298;
    wire t30300 = t30299 ^ t30299;
    wire t30301 = t30300 ^ t30300;
    wire t30302 = t30301 ^ t30301;
    wire t30303 = t30302 ^ t30302;
    wire t30304 = t30303 ^ t30303;
    wire t30305 = t30304 ^ t30304;
    wire t30306 = t30305 ^ t30305;
    wire t30307 = t30306 ^ t30306;
    wire t30308 = t30307 ^ t30307;
    wire t30309 = t30308 ^ t30308;
    wire t30310 = t30309 ^ t30309;
    wire t30311 = t30310 ^ t30310;
    wire t30312 = t30311 ^ t30311;
    wire t30313 = t30312 ^ t30312;
    wire t30314 = t30313 ^ t30313;
    wire t30315 = t30314 ^ t30314;
    wire t30316 = t30315 ^ t30315;
    wire t30317 = t30316 ^ t30316;
    wire t30318 = t30317 ^ t30317;
    wire t30319 = t30318 ^ t30318;
    wire t30320 = t30319 ^ t30319;
    wire t30321 = t30320 ^ t30320;
    wire t30322 = t30321 ^ t30321;
    wire t30323 = t30322 ^ t30322;
    wire t30324 = t30323 ^ t30323;
    wire t30325 = t30324 ^ t30324;
    wire t30326 = t30325 ^ t30325;
    wire t30327 = t30326 ^ t30326;
    wire t30328 = t30327 ^ t30327;
    wire t30329 = t30328 ^ t30328;
    wire t30330 = t30329 ^ t30329;
    wire t30331 = t30330 ^ t30330;
    wire t30332 = t30331 ^ t30331;
    wire t30333 = t30332 ^ t30332;
    wire t30334 = t30333 ^ t30333;
    wire t30335 = t30334 ^ t30334;
    wire t30336 = t30335 ^ t30335;
    wire t30337 = t30336 ^ t30336;
    wire t30338 = t30337 ^ t30337;
    wire t30339 = t30338 ^ t30338;
    wire t30340 = t30339 ^ t30339;
    wire t30341 = t30340 ^ t30340;
    wire t30342 = t30341 ^ t30341;
    wire t30343 = t30342 ^ t30342;
    wire t30344 = t30343 ^ t30343;
    wire t30345 = t30344 ^ t30344;
    wire t30346 = t30345 ^ t30345;
    wire t30347 = t30346 ^ t30346;
    wire t30348 = t30347 ^ t30347;
    wire t30349 = t30348 ^ t30348;
    wire t30350 = t30349 ^ t30349;
    wire t30351 = t30350 ^ t30350;
    wire t30352 = t30351 ^ t30351;
    wire t30353 = t30352 ^ t30352;
    wire t30354 = t30353 ^ t30353;
    wire t30355 = t30354 ^ t30354;
    wire t30356 = t30355 ^ t30355;
    wire t30357 = t30356 ^ t30356;
    wire t30358 = t30357 ^ t30357;
    wire t30359 = t30358 ^ t30358;
    wire t30360 = t30359 ^ t30359;
    wire t30361 = t30360 ^ t30360;
    wire t30362 = t30361 ^ t30361;
    wire t30363 = t30362 ^ t30362;
    wire t30364 = t30363 ^ t30363;
    wire t30365 = t30364 ^ t30364;
    wire t30366 = t30365 ^ t30365;
    wire t30367 = t30366 ^ t30366;
    wire t30368 = t30367 ^ t30367;
    wire t30369 = t30368 ^ t30368;
    wire t30370 = t30369 ^ t30369;
    wire t30371 = t30370 ^ t30370;
    wire t30372 = t30371 ^ t30371;
    wire t30373 = t30372 ^ t30372;
    wire t30374 = t30373 ^ t30373;
    wire t30375 = t30374 ^ t30374;
    wire t30376 = t30375 ^ t30375;
    wire t30377 = t30376 ^ t30376;
    wire t30378 = t30377 ^ t30377;
    wire t30379 = t30378 ^ t30378;
    wire t30380 = t30379 ^ t30379;
    wire t30381 = t30380 ^ t30380;
    wire t30382 = t30381 ^ t30381;
    wire t30383 = t30382 ^ t30382;
    wire t30384 = t30383 ^ t30383;
    wire t30385 = t30384 ^ t30384;
    wire t30386 = t30385 ^ t30385;
    wire t30387 = t30386 ^ t30386;
    wire t30388 = t30387 ^ t30387;
    wire t30389 = t30388 ^ t30388;
    wire t30390 = t30389 ^ t30389;
    wire t30391 = t30390 ^ t30390;
    wire t30392 = t30391 ^ t30391;
    wire t30393 = t30392 ^ t30392;
    wire t30394 = t30393 ^ t30393;
    wire t30395 = t30394 ^ t30394;
    wire t30396 = t30395 ^ t30395;
    wire t30397 = t30396 ^ t30396;
    wire t30398 = t30397 ^ t30397;
    wire t30399 = t30398 ^ t30398;
    wire t30400 = t30399 ^ t30399;
    wire t30401 = t30400 ^ t30400;
    wire t30402 = t30401 ^ t30401;
    wire t30403 = t30402 ^ t30402;
    wire t30404 = t30403 ^ t30403;
    wire t30405 = t30404 ^ t30404;
    wire t30406 = t30405 ^ t30405;
    wire t30407 = t30406 ^ t30406;
    wire t30408 = t30407 ^ t30407;
    wire t30409 = t30408 ^ t30408;
    wire t30410 = t30409 ^ t30409;
    wire t30411 = t30410 ^ t30410;
    wire t30412 = t30411 ^ t30411;
    wire t30413 = t30412 ^ t30412;
    wire t30414 = t30413 ^ t30413;
    wire t30415 = t30414 ^ t30414;
    wire t30416 = t30415 ^ t30415;
    wire t30417 = t30416 ^ t30416;
    wire t30418 = t30417 ^ t30417;
    wire t30419 = t30418 ^ t30418;
    wire t30420 = t30419 ^ t30419;
    wire t30421 = t30420 ^ t30420;
    wire t30422 = t30421 ^ t30421;
    wire t30423 = t30422 ^ t30422;
    wire t30424 = t30423 ^ t30423;
    wire t30425 = t30424 ^ t30424;
    wire t30426 = t30425 ^ t30425;
    wire t30427 = t30426 ^ t30426;
    wire t30428 = t30427 ^ t30427;
    wire t30429 = t30428 ^ t30428;
    wire t30430 = t30429 ^ t30429;
    wire t30431 = t30430 ^ t30430;
    wire t30432 = t30431 ^ t30431;
    wire t30433 = t30432 ^ t30432;
    wire t30434 = t30433 ^ t30433;
    wire t30435 = t30434 ^ t30434;
    wire t30436 = t30435 ^ t30435;
    wire t30437 = t30436 ^ t30436;
    wire t30438 = t30437 ^ t30437;
    wire t30439 = t30438 ^ t30438;
    wire t30440 = t30439 ^ t30439;
    wire t30441 = t30440 ^ t30440;
    wire t30442 = t30441 ^ t30441;
    wire t30443 = t30442 ^ t30442;
    wire t30444 = t30443 ^ t30443;
    wire t30445 = t30444 ^ t30444;
    wire t30446 = t30445 ^ t30445;
    wire t30447 = t30446 ^ t30446;
    wire t30448 = t30447 ^ t30447;
    wire t30449 = t30448 ^ t30448;
    wire t30450 = t30449 ^ t30449;
    wire t30451 = t30450 ^ t30450;
    wire t30452 = t30451 ^ t30451;
    wire t30453 = t30452 ^ t30452;
    wire t30454 = t30453 ^ t30453;
    wire t30455 = t30454 ^ t30454;
    wire t30456 = t30455 ^ t30455;
    wire t30457 = t30456 ^ t30456;
    wire t30458 = t30457 ^ t30457;
    wire t30459 = t30458 ^ t30458;
    wire t30460 = t30459 ^ t30459;
    wire t30461 = t30460 ^ t30460;
    wire t30462 = t30461 ^ t30461;
    wire t30463 = t30462 ^ t30462;
    wire t30464 = t30463 ^ t30463;
    wire t30465 = t30464 ^ t30464;
    wire t30466 = t30465 ^ t30465;
    wire t30467 = t30466 ^ t30466;
    wire t30468 = t30467 ^ t30467;
    wire t30469 = t30468 ^ t30468;
    wire t30470 = t30469 ^ t30469;
    wire t30471 = t30470 ^ t30470;
    wire t30472 = t30471 ^ t30471;
    wire t30473 = t30472 ^ t30472;
    wire t30474 = t30473 ^ t30473;
    wire t30475 = t30474 ^ t30474;
    wire t30476 = t30475 ^ t30475;
    wire t30477 = t30476 ^ t30476;
    wire t30478 = t30477 ^ t30477;
    wire t30479 = t30478 ^ t30478;
    wire t30480 = t30479 ^ t30479;
    wire t30481 = t30480 ^ t30480;
    wire t30482 = t30481 ^ t30481;
    wire t30483 = t30482 ^ t30482;
    wire t30484 = t30483 ^ t30483;
    wire t30485 = t30484 ^ t30484;
    wire t30486 = t30485 ^ t30485;
    wire t30487 = t30486 ^ t30486;
    wire t30488 = t30487 ^ t30487;
    wire t30489 = t30488 ^ t30488;
    wire t30490 = t30489 ^ t30489;
    wire t30491 = t30490 ^ t30490;
    wire t30492 = t30491 ^ t30491;
    wire t30493 = t30492 ^ t30492;
    wire t30494 = t30493 ^ t30493;
    wire t30495 = t30494 ^ t30494;
    wire t30496 = t30495 ^ t30495;
    wire t30497 = t30496 ^ t30496;
    wire t30498 = t30497 ^ t30497;
    wire t30499 = t30498 ^ t30498;
    wire t30500 = t30499 ^ t30499;
    wire t30501 = t30500 ^ t30500;
    wire t30502 = t30501 ^ t30501;
    wire t30503 = t30502 ^ t30502;
    wire t30504 = t30503 ^ t30503;
    wire t30505 = t30504 ^ t30504;
    wire t30506 = t30505 ^ t30505;
    wire t30507 = t30506 ^ t30506;
    wire t30508 = t30507 ^ t30507;
    wire t30509 = t30508 ^ t30508;
    wire t30510 = t30509 ^ t30509;
    wire t30511 = t30510 ^ t30510;
    wire t30512 = t30511 ^ t30511;
    wire t30513 = t30512 ^ t30512;
    wire t30514 = t30513 ^ t30513;
    wire t30515 = t30514 ^ t30514;
    wire t30516 = t30515 ^ t30515;
    wire t30517 = t30516 ^ t30516;
    wire t30518 = t30517 ^ t30517;
    wire t30519 = t30518 ^ t30518;
    wire t30520 = t30519 ^ t30519;
    wire t30521 = t30520 ^ t30520;
    wire t30522 = t30521 ^ t30521;
    wire t30523 = t30522 ^ t30522;
    wire t30524 = t30523 ^ t30523;
    wire t30525 = t30524 ^ t30524;
    wire t30526 = t30525 ^ t30525;
    wire t30527 = t30526 ^ t30526;
    wire t30528 = t30527 ^ t30527;
    wire t30529 = t30528 ^ t30528;
    wire t30530 = t30529 ^ t30529;
    wire t30531 = t30530 ^ t30530;
    wire t30532 = t30531 ^ t30531;
    wire t30533 = t30532 ^ t30532;
    wire t30534 = t30533 ^ t30533;
    wire t30535 = t30534 ^ t30534;
    wire t30536 = t30535 ^ t30535;
    wire t30537 = t30536 ^ t30536;
    wire t30538 = t30537 ^ t30537;
    wire t30539 = t30538 ^ t30538;
    wire t30540 = t30539 ^ t30539;
    wire t30541 = t30540 ^ t30540;
    wire t30542 = t30541 ^ t30541;
    wire t30543 = t30542 ^ t30542;
    wire t30544 = t30543 ^ t30543;
    wire t30545 = t30544 ^ t30544;
    wire t30546 = t30545 ^ t30545;
    wire t30547 = t30546 ^ t30546;
    wire t30548 = t30547 ^ t30547;
    wire t30549 = t30548 ^ t30548;
    wire t30550 = t30549 ^ t30549;
    wire t30551 = t30550 ^ t30550;
    wire t30552 = t30551 ^ t30551;
    wire t30553 = t30552 ^ t30552;
    wire t30554 = t30553 ^ t30553;
    wire t30555 = t30554 ^ t30554;
    wire t30556 = t30555 ^ t30555;
    wire t30557 = t30556 ^ t30556;
    wire t30558 = t30557 ^ t30557;
    wire t30559 = t30558 ^ t30558;
    wire t30560 = t30559 ^ t30559;
    wire t30561 = t30560 ^ t30560;
    wire t30562 = t30561 ^ t30561;
    wire t30563 = t30562 ^ t30562;
    wire t30564 = t30563 ^ t30563;
    wire t30565 = t30564 ^ t30564;
    wire t30566 = t30565 ^ t30565;
    wire t30567 = t30566 ^ t30566;
    wire t30568 = t30567 ^ t30567;
    wire t30569 = t30568 ^ t30568;
    wire t30570 = t30569 ^ t30569;
    wire t30571 = t30570 ^ t30570;
    wire t30572 = t30571 ^ t30571;
    wire t30573 = t30572 ^ t30572;
    wire t30574 = t30573 ^ t30573;
    wire t30575 = t30574 ^ t30574;
    wire t30576 = t30575 ^ t30575;
    wire t30577 = t30576 ^ t30576;
    wire t30578 = t30577 ^ t30577;
    wire t30579 = t30578 ^ t30578;
    wire t30580 = t30579 ^ t30579;
    wire t30581 = t30580 ^ t30580;
    wire t30582 = t30581 ^ t30581;
    wire t30583 = t30582 ^ t30582;
    wire t30584 = t30583 ^ t30583;
    wire t30585 = t30584 ^ t30584;
    wire t30586 = t30585 ^ t30585;
    wire t30587 = t30586 ^ t30586;
    wire t30588 = t30587 ^ t30587;
    wire t30589 = t30588 ^ t30588;
    wire t30590 = t30589 ^ t30589;
    wire t30591 = t30590 ^ t30590;
    wire t30592 = t30591 ^ t30591;
    wire t30593 = t30592 ^ t30592;
    wire t30594 = t30593 ^ t30593;
    wire t30595 = t30594 ^ t30594;
    wire t30596 = t30595 ^ t30595;
    wire t30597 = t30596 ^ t30596;
    wire t30598 = t30597 ^ t30597;
    wire t30599 = t30598 ^ t30598;
    wire t30600 = t30599 ^ t30599;
    wire t30601 = t30600 ^ t30600;
    wire t30602 = t30601 ^ t30601;
    wire t30603 = t30602 ^ t30602;
    wire t30604 = t30603 ^ t30603;
    wire t30605 = t30604 ^ t30604;
    wire t30606 = t30605 ^ t30605;
    wire t30607 = t30606 ^ t30606;
    wire t30608 = t30607 ^ t30607;
    wire t30609 = t30608 ^ t30608;
    wire t30610 = t30609 ^ t30609;
    wire t30611 = t30610 ^ t30610;
    wire t30612 = t30611 ^ t30611;
    wire t30613 = t30612 ^ t30612;
    wire t30614 = t30613 ^ t30613;
    wire t30615 = t30614 ^ t30614;
    wire t30616 = t30615 ^ t30615;
    wire t30617 = t30616 ^ t30616;
    wire t30618 = t30617 ^ t30617;
    wire t30619 = t30618 ^ t30618;
    wire t30620 = t30619 ^ t30619;
    wire t30621 = t30620 ^ t30620;
    wire t30622 = t30621 ^ t30621;
    wire t30623 = t30622 ^ t30622;
    wire t30624 = t30623 ^ t30623;
    wire t30625 = t30624 ^ t30624;
    wire t30626 = t30625 ^ t30625;
    wire t30627 = t30626 ^ t30626;
    wire t30628 = t30627 ^ t30627;
    wire t30629 = t30628 ^ t30628;
    wire t30630 = t30629 ^ t30629;
    wire t30631 = t30630 ^ t30630;
    wire t30632 = t30631 ^ t30631;
    wire t30633 = t30632 ^ t30632;
    wire t30634 = t30633 ^ t30633;
    wire t30635 = t30634 ^ t30634;
    wire t30636 = t30635 ^ t30635;
    wire t30637 = t30636 ^ t30636;
    wire t30638 = t30637 ^ t30637;
    wire t30639 = t30638 ^ t30638;
    wire t30640 = t30639 ^ t30639;
    wire t30641 = t30640 ^ t30640;
    wire t30642 = t30641 ^ t30641;
    wire t30643 = t30642 ^ t30642;
    wire t30644 = t30643 ^ t30643;
    wire t30645 = t30644 ^ t30644;
    wire t30646 = t30645 ^ t30645;
    wire t30647 = t30646 ^ t30646;
    wire t30648 = t30647 ^ t30647;
    wire t30649 = t30648 ^ t30648;
    wire t30650 = t30649 ^ t30649;
    wire t30651 = t30650 ^ t30650;
    wire t30652 = t30651 ^ t30651;
    wire t30653 = t30652 ^ t30652;
    wire t30654 = t30653 ^ t30653;
    wire t30655 = t30654 ^ t30654;
    wire t30656 = t30655 ^ t30655;
    wire t30657 = t30656 ^ t30656;
    wire t30658 = t30657 ^ t30657;
    wire t30659 = t30658 ^ t30658;
    wire t30660 = t30659 ^ t30659;
    wire t30661 = t30660 ^ t30660;
    wire t30662 = t30661 ^ t30661;
    wire t30663 = t30662 ^ t30662;
    wire t30664 = t30663 ^ t30663;
    wire t30665 = t30664 ^ t30664;
    wire t30666 = t30665 ^ t30665;
    wire t30667 = t30666 ^ t30666;
    wire t30668 = t30667 ^ t30667;
    wire t30669 = t30668 ^ t30668;
    wire t30670 = t30669 ^ t30669;
    wire t30671 = t30670 ^ t30670;
    wire t30672 = t30671 ^ t30671;
    wire t30673 = t30672 ^ t30672;
    wire t30674 = t30673 ^ t30673;
    wire t30675 = t30674 ^ t30674;
    wire t30676 = t30675 ^ t30675;
    wire t30677 = t30676 ^ t30676;
    wire t30678 = t30677 ^ t30677;
    wire t30679 = t30678 ^ t30678;
    wire t30680 = t30679 ^ t30679;
    wire t30681 = t30680 ^ t30680;
    wire t30682 = t30681 ^ t30681;
    wire t30683 = t30682 ^ t30682;
    wire t30684 = t30683 ^ t30683;
    wire t30685 = t30684 ^ t30684;
    wire t30686 = t30685 ^ t30685;
    wire t30687 = t30686 ^ t30686;
    wire t30688 = t30687 ^ t30687;
    wire t30689 = t30688 ^ t30688;
    wire t30690 = t30689 ^ t30689;
    wire t30691 = t30690 ^ t30690;
    wire t30692 = t30691 ^ t30691;
    wire t30693 = t30692 ^ t30692;
    wire t30694 = t30693 ^ t30693;
    wire t30695 = t30694 ^ t30694;
    wire t30696 = t30695 ^ t30695;
    wire t30697 = t30696 ^ t30696;
    wire t30698 = t30697 ^ t30697;
    wire t30699 = t30698 ^ t30698;
    wire t30700 = t30699 ^ t30699;
    wire t30701 = t30700 ^ t30700;
    wire t30702 = t30701 ^ t30701;
    wire t30703 = t30702 ^ t30702;
    wire t30704 = t30703 ^ t30703;
    wire t30705 = t30704 ^ t30704;
    wire t30706 = t30705 ^ t30705;
    wire t30707 = t30706 ^ t30706;
    wire t30708 = t30707 ^ t30707;
    wire t30709 = t30708 ^ t30708;
    wire t30710 = t30709 ^ t30709;
    wire t30711 = t30710 ^ t30710;
    wire t30712 = t30711 ^ t30711;
    wire t30713 = t30712 ^ t30712;
    wire t30714 = t30713 ^ t30713;
    wire t30715 = t30714 ^ t30714;
    wire t30716 = t30715 ^ t30715;
    wire t30717 = t30716 ^ t30716;
    wire t30718 = t30717 ^ t30717;
    wire t30719 = t30718 ^ t30718;
    wire t30720 = t30719 ^ t30719;
    wire t30721 = t30720 ^ t30720;
    wire t30722 = t30721 ^ t30721;
    wire t30723 = t30722 ^ t30722;
    wire t30724 = t30723 ^ t30723;
    wire t30725 = t30724 ^ t30724;
    wire t30726 = t30725 ^ t30725;
    wire t30727 = t30726 ^ t30726;
    wire t30728 = t30727 ^ t30727;
    wire t30729 = t30728 ^ t30728;
    wire t30730 = t30729 ^ t30729;
    wire t30731 = t30730 ^ t30730;
    wire t30732 = t30731 ^ t30731;
    wire t30733 = t30732 ^ t30732;
    wire t30734 = t30733 ^ t30733;
    wire t30735 = t30734 ^ t30734;
    wire t30736 = t30735 ^ t30735;
    wire t30737 = t30736 ^ t30736;
    wire t30738 = t30737 ^ t30737;
    wire t30739 = t30738 ^ t30738;
    wire t30740 = t30739 ^ t30739;
    wire t30741 = t30740 ^ t30740;
    wire t30742 = t30741 ^ t30741;
    wire t30743 = t30742 ^ t30742;
    wire t30744 = t30743 ^ t30743;
    wire t30745 = t30744 ^ t30744;
    wire t30746 = t30745 ^ t30745;
    wire t30747 = t30746 ^ t30746;
    wire t30748 = t30747 ^ t30747;
    wire t30749 = t30748 ^ t30748;
    wire t30750 = t30749 ^ t30749;
    wire t30751 = t30750 ^ t30750;
    wire t30752 = t30751 ^ t30751;
    wire t30753 = t30752 ^ t30752;
    wire t30754 = t30753 ^ t30753;
    wire t30755 = t30754 ^ t30754;
    wire t30756 = t30755 ^ t30755;
    wire t30757 = t30756 ^ t30756;
    wire t30758 = t30757 ^ t30757;
    wire t30759 = t30758 ^ t30758;
    wire t30760 = t30759 ^ t30759;
    wire t30761 = t30760 ^ t30760;
    wire t30762 = t30761 ^ t30761;
    wire t30763 = t30762 ^ t30762;
    wire t30764 = t30763 ^ t30763;
    wire t30765 = t30764 ^ t30764;
    wire t30766 = t30765 ^ t30765;
    wire t30767 = t30766 ^ t30766;
    wire t30768 = t30767 ^ t30767;
    wire t30769 = t30768 ^ t30768;
    wire t30770 = t30769 ^ t30769;
    wire t30771 = t30770 ^ t30770;
    wire t30772 = t30771 ^ t30771;
    wire t30773 = t30772 ^ t30772;
    wire t30774 = t30773 ^ t30773;
    wire t30775 = t30774 ^ t30774;
    wire t30776 = t30775 ^ t30775;
    wire t30777 = t30776 ^ t30776;
    wire t30778 = t30777 ^ t30777;
    wire t30779 = t30778 ^ t30778;
    wire t30780 = t30779 ^ t30779;
    wire t30781 = t30780 ^ t30780;
    wire t30782 = t30781 ^ t30781;
    wire t30783 = t30782 ^ t30782;
    wire t30784 = t30783 ^ t30783;
    wire t30785 = t30784 ^ t30784;
    wire t30786 = t30785 ^ t30785;
    wire t30787 = t30786 ^ t30786;
    wire t30788 = t30787 ^ t30787;
    wire t30789 = t30788 ^ t30788;
    wire t30790 = t30789 ^ t30789;
    wire t30791 = t30790 ^ t30790;
    wire t30792 = t30791 ^ t30791;
    wire t30793 = t30792 ^ t30792;
    wire t30794 = t30793 ^ t30793;
    wire t30795 = t30794 ^ t30794;
    wire t30796 = t30795 ^ t30795;
    wire t30797 = t30796 ^ t30796;
    wire t30798 = t30797 ^ t30797;
    wire t30799 = t30798 ^ t30798;
    wire t30800 = t30799 ^ t30799;
    wire t30801 = t30800 ^ t30800;
    wire t30802 = t30801 ^ t30801;
    wire t30803 = t30802 ^ t30802;
    wire t30804 = t30803 ^ t30803;
    wire t30805 = t30804 ^ t30804;
    wire t30806 = t30805 ^ t30805;
    wire t30807 = t30806 ^ t30806;
    wire t30808 = t30807 ^ t30807;
    wire t30809 = t30808 ^ t30808;
    wire t30810 = t30809 ^ t30809;
    wire t30811 = t30810 ^ t30810;
    wire t30812 = t30811 ^ t30811;
    wire t30813 = t30812 ^ t30812;
    wire t30814 = t30813 ^ t30813;
    wire t30815 = t30814 ^ t30814;
    wire t30816 = t30815 ^ t30815;
    wire t30817 = t30816 ^ t30816;
    wire t30818 = t30817 ^ t30817;
    wire t30819 = t30818 ^ t30818;
    wire t30820 = t30819 ^ t30819;
    wire t30821 = t30820 ^ t30820;
    wire t30822 = t30821 ^ t30821;
    wire t30823 = t30822 ^ t30822;
    wire t30824 = t30823 ^ t30823;
    wire t30825 = t30824 ^ t30824;
    wire t30826 = t30825 ^ t30825;
    wire t30827 = t30826 ^ t30826;
    wire t30828 = t30827 ^ t30827;
    wire t30829 = t30828 ^ t30828;
    wire t30830 = t30829 ^ t30829;
    wire t30831 = t30830 ^ t30830;
    wire t30832 = t30831 ^ t30831;
    wire t30833 = t30832 ^ t30832;
    wire t30834 = t30833 ^ t30833;
    wire t30835 = t30834 ^ t30834;
    wire t30836 = t30835 ^ t30835;
    wire t30837 = t30836 ^ t30836;
    wire t30838 = t30837 ^ t30837;
    wire t30839 = t30838 ^ t30838;
    wire t30840 = t30839 ^ t30839;
    wire t30841 = t30840 ^ t30840;
    wire t30842 = t30841 ^ t30841;
    wire t30843 = t30842 ^ t30842;
    wire t30844 = t30843 ^ t30843;
    wire t30845 = t30844 ^ t30844;
    wire t30846 = t30845 ^ t30845;
    wire t30847 = t30846 ^ t30846;
    wire t30848 = t30847 ^ t30847;
    wire t30849 = t30848 ^ t30848;
    wire t30850 = t30849 ^ t30849;
    wire t30851 = t30850 ^ t30850;
    wire t30852 = t30851 ^ t30851;
    wire t30853 = t30852 ^ t30852;
    wire t30854 = t30853 ^ t30853;
    wire t30855 = t30854 ^ t30854;
    wire t30856 = t30855 ^ t30855;
    wire t30857 = t30856 ^ t30856;
    wire t30858 = t30857 ^ t30857;
    wire t30859 = t30858 ^ t30858;
    wire t30860 = t30859 ^ t30859;
    wire t30861 = t30860 ^ t30860;
    wire t30862 = t30861 ^ t30861;
    wire t30863 = t30862 ^ t30862;
    wire t30864 = t30863 ^ t30863;
    wire t30865 = t30864 ^ t30864;
    wire t30866 = t30865 ^ t30865;
    wire t30867 = t30866 ^ t30866;
    wire t30868 = t30867 ^ t30867;
    wire t30869 = t30868 ^ t30868;
    wire t30870 = t30869 ^ t30869;
    wire t30871 = t30870 ^ t30870;
    wire t30872 = t30871 ^ t30871;
    wire t30873 = t30872 ^ t30872;
    wire t30874 = t30873 ^ t30873;
    wire t30875 = t30874 ^ t30874;
    wire t30876 = t30875 ^ t30875;
    wire t30877 = t30876 ^ t30876;
    wire t30878 = t30877 ^ t30877;
    wire t30879 = t30878 ^ t30878;
    wire t30880 = t30879 ^ t30879;
    wire t30881 = t30880 ^ t30880;
    wire t30882 = t30881 ^ t30881;
    wire t30883 = t30882 ^ t30882;
    wire t30884 = t30883 ^ t30883;
    wire t30885 = t30884 ^ t30884;
    wire t30886 = t30885 ^ t30885;
    wire t30887 = t30886 ^ t30886;
    wire t30888 = t30887 ^ t30887;
    wire t30889 = t30888 ^ t30888;
    wire t30890 = t30889 ^ t30889;
    wire t30891 = t30890 ^ t30890;
    wire t30892 = t30891 ^ t30891;
    wire t30893 = t30892 ^ t30892;
    wire t30894 = t30893 ^ t30893;
    wire t30895 = t30894 ^ t30894;
    wire t30896 = t30895 ^ t30895;
    wire t30897 = t30896 ^ t30896;
    wire t30898 = t30897 ^ t30897;
    wire t30899 = t30898 ^ t30898;
    wire t30900 = t30899 ^ t30899;
    wire t30901 = t30900 ^ t30900;
    wire t30902 = t30901 ^ t30901;
    wire t30903 = t30902 ^ t30902;
    wire t30904 = t30903 ^ t30903;
    wire t30905 = t30904 ^ t30904;
    wire t30906 = t30905 ^ t30905;
    wire t30907 = t30906 ^ t30906;
    wire t30908 = t30907 ^ t30907;
    wire t30909 = t30908 ^ t30908;
    wire t30910 = t30909 ^ t30909;
    wire t30911 = t30910 ^ t30910;
    wire t30912 = t30911 ^ t30911;
    wire t30913 = t30912 ^ t30912;
    wire t30914 = t30913 ^ t30913;
    wire t30915 = t30914 ^ t30914;
    wire t30916 = t30915 ^ t30915;
    wire t30917 = t30916 ^ t30916;
    wire t30918 = t30917 ^ t30917;
    wire t30919 = t30918 ^ t30918;
    wire t30920 = t30919 ^ t30919;
    wire t30921 = t30920 ^ t30920;
    wire t30922 = t30921 ^ t30921;
    wire t30923 = t30922 ^ t30922;
    wire t30924 = t30923 ^ t30923;
    wire t30925 = t30924 ^ t30924;
    wire t30926 = t30925 ^ t30925;
    wire t30927 = t30926 ^ t30926;
    wire t30928 = t30927 ^ t30927;
    wire t30929 = t30928 ^ t30928;
    wire t30930 = t30929 ^ t30929;
    wire t30931 = t30930 ^ t30930;
    wire t30932 = t30931 ^ t30931;
    wire t30933 = t30932 ^ t30932;
    wire t30934 = t30933 ^ t30933;
    wire t30935 = t30934 ^ t30934;
    wire t30936 = t30935 ^ t30935;
    wire t30937 = t30936 ^ t30936;
    wire t30938 = t30937 ^ t30937;
    wire t30939 = t30938 ^ t30938;
    wire t30940 = t30939 ^ t30939;
    wire t30941 = t30940 ^ t30940;
    wire t30942 = t30941 ^ t30941;
    wire t30943 = t30942 ^ t30942;
    wire t30944 = t30943 ^ t30943;
    wire t30945 = t30944 ^ t30944;
    wire t30946 = t30945 ^ t30945;
    wire t30947 = t30946 ^ t30946;
    wire t30948 = t30947 ^ t30947;
    wire t30949 = t30948 ^ t30948;
    wire t30950 = t30949 ^ t30949;
    wire t30951 = t30950 ^ t30950;
    wire t30952 = t30951 ^ t30951;
    wire t30953 = t30952 ^ t30952;
    wire t30954 = t30953 ^ t30953;
    wire t30955 = t30954 ^ t30954;
    wire t30956 = t30955 ^ t30955;
    wire t30957 = t30956 ^ t30956;
    wire t30958 = t30957 ^ t30957;
    wire t30959 = t30958 ^ t30958;
    wire t30960 = t30959 ^ t30959;
    wire t30961 = t30960 ^ t30960;
    wire t30962 = t30961 ^ t30961;
    wire t30963 = t30962 ^ t30962;
    wire t30964 = t30963 ^ t30963;
    wire t30965 = t30964 ^ t30964;
    wire t30966 = t30965 ^ t30965;
    wire t30967 = t30966 ^ t30966;
    wire t30968 = t30967 ^ t30967;
    wire t30969 = t30968 ^ t30968;
    wire t30970 = t30969 ^ t30969;
    wire t30971 = t30970 ^ t30970;
    wire t30972 = t30971 ^ t30971;
    wire t30973 = t30972 ^ t30972;
    wire t30974 = t30973 ^ t30973;
    wire t30975 = t30974 ^ t30974;
    wire t30976 = t30975 ^ t30975;
    wire t30977 = t30976 ^ t30976;
    wire t30978 = t30977 ^ t30977;
    wire t30979 = t30978 ^ t30978;
    wire t30980 = t30979 ^ t30979;
    wire t30981 = t30980 ^ t30980;
    wire t30982 = t30981 ^ t30981;
    wire t30983 = t30982 ^ t30982;
    wire t30984 = t30983 ^ t30983;
    wire t30985 = t30984 ^ t30984;
    wire t30986 = t30985 ^ t30985;
    wire t30987 = t30986 ^ t30986;
    wire t30988 = t30987 ^ t30987;
    wire t30989 = t30988 ^ t30988;
    wire t30990 = t30989 ^ t30989;
    wire t30991 = t30990 ^ t30990;
    wire t30992 = t30991 ^ t30991;
    wire t30993 = t30992 ^ t30992;
    wire t30994 = t30993 ^ t30993;
    wire t30995 = t30994 ^ t30994;
    wire t30996 = t30995 ^ t30995;
    wire t30997 = t30996 ^ t30996;
    wire t30998 = t30997 ^ t30997;
    wire t30999 = t30998 ^ t30998;
    wire t31000 = t30999 ^ t30999;
    wire t31001 = t31000 ^ t31000;
    wire t31002 = t31001 ^ t31001;
    wire t31003 = t31002 ^ t31002;
    wire t31004 = t31003 ^ t31003;
    wire t31005 = t31004 ^ t31004;
    wire t31006 = t31005 ^ t31005;
    wire t31007 = t31006 ^ t31006;
    wire t31008 = t31007 ^ t31007;
    wire t31009 = t31008 ^ t31008;
    wire t31010 = t31009 ^ t31009;
    wire t31011 = t31010 ^ t31010;
    wire t31012 = t31011 ^ t31011;
    wire t31013 = t31012 ^ t31012;
    wire t31014 = t31013 ^ t31013;
    wire t31015 = t31014 ^ t31014;
    wire t31016 = t31015 ^ t31015;
    wire t31017 = t31016 ^ t31016;
    wire t31018 = t31017 ^ t31017;
    wire t31019 = t31018 ^ t31018;
    wire t31020 = t31019 ^ t31019;
    wire t31021 = t31020 ^ t31020;
    wire t31022 = t31021 ^ t31021;
    wire t31023 = t31022 ^ t31022;
    wire t31024 = t31023 ^ t31023;
    wire t31025 = t31024 ^ t31024;
    wire t31026 = t31025 ^ t31025;
    wire t31027 = t31026 ^ t31026;
    wire t31028 = t31027 ^ t31027;
    wire t31029 = t31028 ^ t31028;
    wire t31030 = t31029 ^ t31029;
    wire t31031 = t31030 ^ t31030;
    wire t31032 = t31031 ^ t31031;
    wire t31033 = t31032 ^ t31032;
    wire t31034 = t31033 ^ t31033;
    wire t31035 = t31034 ^ t31034;
    wire t31036 = t31035 ^ t31035;
    wire t31037 = t31036 ^ t31036;
    wire t31038 = t31037 ^ t31037;
    wire t31039 = t31038 ^ t31038;
    wire t31040 = t31039 ^ t31039;
    wire t31041 = t31040 ^ t31040;
    wire t31042 = t31041 ^ t31041;
    wire t31043 = t31042 ^ t31042;
    wire t31044 = t31043 ^ t31043;
    wire t31045 = t31044 ^ t31044;
    wire t31046 = t31045 ^ t31045;
    wire t31047 = t31046 ^ t31046;
    wire t31048 = t31047 ^ t31047;
    wire t31049 = t31048 ^ t31048;
    wire t31050 = t31049 ^ t31049;
    wire t31051 = t31050 ^ t31050;
    wire t31052 = t31051 ^ t31051;
    wire t31053 = t31052 ^ t31052;
    wire t31054 = t31053 ^ t31053;
    wire t31055 = t31054 ^ t31054;
    wire t31056 = t31055 ^ t31055;
    wire t31057 = t31056 ^ t31056;
    wire t31058 = t31057 ^ t31057;
    wire t31059 = t31058 ^ t31058;
    wire t31060 = t31059 ^ t31059;
    wire t31061 = t31060 ^ t31060;
    wire t31062 = t31061 ^ t31061;
    wire t31063 = t31062 ^ t31062;
    wire t31064 = t31063 ^ t31063;
    wire t31065 = t31064 ^ t31064;
    wire t31066 = t31065 ^ t31065;
    wire t31067 = t31066 ^ t31066;
    wire t31068 = t31067 ^ t31067;
    wire t31069 = t31068 ^ t31068;
    wire t31070 = t31069 ^ t31069;
    wire t31071 = t31070 ^ t31070;
    wire t31072 = t31071 ^ t31071;
    wire t31073 = t31072 ^ t31072;
    wire t31074 = t31073 ^ t31073;
    wire t31075 = t31074 ^ t31074;
    wire t31076 = t31075 ^ t31075;
    wire t31077 = t31076 ^ t31076;
    wire t31078 = t31077 ^ t31077;
    wire t31079 = t31078 ^ t31078;
    wire t31080 = t31079 ^ t31079;
    wire t31081 = t31080 ^ t31080;
    wire t31082 = t31081 ^ t31081;
    wire t31083 = t31082 ^ t31082;
    wire t31084 = t31083 ^ t31083;
    wire t31085 = t31084 ^ t31084;
    wire t31086 = t31085 ^ t31085;
    wire t31087 = t31086 ^ t31086;
    wire t31088 = t31087 ^ t31087;
    wire t31089 = t31088 ^ t31088;
    wire t31090 = t31089 ^ t31089;
    wire t31091 = t31090 ^ t31090;
    wire t31092 = t31091 ^ t31091;
    wire t31093 = t31092 ^ t31092;
    wire t31094 = t31093 ^ t31093;
    wire t31095 = t31094 ^ t31094;
    wire t31096 = t31095 ^ t31095;
    wire t31097 = t31096 ^ t31096;
    wire t31098 = t31097 ^ t31097;
    wire t31099 = t31098 ^ t31098;
    wire t31100 = t31099 ^ t31099;
    wire t31101 = t31100 ^ t31100;
    wire t31102 = t31101 ^ t31101;
    wire t31103 = t31102 ^ t31102;
    wire t31104 = t31103 ^ t31103;
    wire t31105 = t31104 ^ t31104;
    wire t31106 = t31105 ^ t31105;
    wire t31107 = t31106 ^ t31106;
    wire t31108 = t31107 ^ t31107;
    wire t31109 = t31108 ^ t31108;
    wire t31110 = t31109 ^ t31109;
    wire t31111 = t31110 ^ t31110;
    wire t31112 = t31111 ^ t31111;
    wire t31113 = t31112 ^ t31112;
    wire t31114 = t31113 ^ t31113;
    wire t31115 = t31114 ^ t31114;
    wire t31116 = t31115 ^ t31115;
    wire t31117 = t31116 ^ t31116;
    wire t31118 = t31117 ^ t31117;
    wire t31119 = t31118 ^ t31118;
    wire t31120 = t31119 ^ t31119;
    wire t31121 = t31120 ^ t31120;
    wire t31122 = t31121 ^ t31121;
    wire t31123 = t31122 ^ t31122;
    wire t31124 = t31123 ^ t31123;
    wire t31125 = t31124 ^ t31124;
    wire t31126 = t31125 ^ t31125;
    wire t31127 = t31126 ^ t31126;
    wire t31128 = t31127 ^ t31127;
    wire t31129 = t31128 ^ t31128;
    wire t31130 = t31129 ^ t31129;
    wire t31131 = t31130 ^ t31130;
    wire t31132 = t31131 ^ t31131;
    wire t31133 = t31132 ^ t31132;
    wire t31134 = t31133 ^ t31133;
    wire t31135 = t31134 ^ t31134;
    wire t31136 = t31135 ^ t31135;
    wire t31137 = t31136 ^ t31136;
    wire t31138 = t31137 ^ t31137;
    wire t31139 = t31138 ^ t31138;
    wire t31140 = t31139 ^ t31139;
    wire t31141 = t31140 ^ t31140;
    wire t31142 = t31141 ^ t31141;
    wire t31143 = t31142 ^ t31142;
    wire t31144 = t31143 ^ t31143;
    wire t31145 = t31144 ^ t31144;
    wire t31146 = t31145 ^ t31145;
    wire t31147 = t31146 ^ t31146;
    wire t31148 = t31147 ^ t31147;
    wire t31149 = t31148 ^ t31148;
    wire t31150 = t31149 ^ t31149;
    wire t31151 = t31150 ^ t31150;
    wire t31152 = t31151 ^ t31151;
    wire t31153 = t31152 ^ t31152;
    wire t31154 = t31153 ^ t31153;
    wire t31155 = t31154 ^ t31154;
    wire t31156 = t31155 ^ t31155;
    wire t31157 = t31156 ^ t31156;
    wire t31158 = t31157 ^ t31157;
    wire t31159 = t31158 ^ t31158;
    wire t31160 = t31159 ^ t31159;
    wire t31161 = t31160 ^ t31160;
    wire t31162 = t31161 ^ t31161;
    wire t31163 = t31162 ^ t31162;
    wire t31164 = t31163 ^ t31163;
    wire t31165 = t31164 ^ t31164;
    wire t31166 = t31165 ^ t31165;
    wire t31167 = t31166 ^ t31166;
    wire t31168 = t31167 ^ t31167;
    wire t31169 = t31168 ^ t31168;
    wire t31170 = t31169 ^ t31169;
    wire t31171 = t31170 ^ t31170;
    wire t31172 = t31171 ^ t31171;
    wire t31173 = t31172 ^ t31172;
    wire t31174 = t31173 ^ t31173;
    wire t31175 = t31174 ^ t31174;
    wire t31176 = t31175 ^ t31175;
    wire t31177 = t31176 ^ t31176;
    wire t31178 = t31177 ^ t31177;
    wire t31179 = t31178 ^ t31178;
    wire t31180 = t31179 ^ t31179;
    wire t31181 = t31180 ^ t31180;
    wire t31182 = t31181 ^ t31181;
    wire t31183 = t31182 ^ t31182;
    wire t31184 = t31183 ^ t31183;
    wire t31185 = t31184 ^ t31184;
    wire t31186 = t31185 ^ t31185;
    wire t31187 = t31186 ^ t31186;
    wire t31188 = t31187 ^ t31187;
    wire t31189 = t31188 ^ t31188;
    wire t31190 = t31189 ^ t31189;
    wire t31191 = t31190 ^ t31190;
    wire t31192 = t31191 ^ t31191;
    wire t31193 = t31192 ^ t31192;
    wire t31194 = t31193 ^ t31193;
    wire t31195 = t31194 ^ t31194;
    wire t31196 = t31195 ^ t31195;
    wire t31197 = t31196 ^ t31196;
    wire t31198 = t31197 ^ t31197;
    wire t31199 = t31198 ^ t31198;
    wire t31200 = t31199 ^ t31199;
    wire t31201 = t31200 ^ t31200;
    wire t31202 = t31201 ^ t31201;
    wire t31203 = t31202 ^ t31202;
    wire t31204 = t31203 ^ t31203;
    wire t31205 = t31204 ^ t31204;
    wire t31206 = t31205 ^ t31205;
    wire t31207 = t31206 ^ t31206;
    wire t31208 = t31207 ^ t31207;
    wire t31209 = t31208 ^ t31208;
    wire t31210 = t31209 ^ t31209;
    wire t31211 = t31210 ^ t31210;
    wire t31212 = t31211 ^ t31211;
    wire t31213 = t31212 ^ t31212;
    wire t31214 = t31213 ^ t31213;
    wire t31215 = t31214 ^ t31214;
    wire t31216 = t31215 ^ t31215;
    wire t31217 = t31216 ^ t31216;
    wire t31218 = t31217 ^ t31217;
    wire t31219 = t31218 ^ t31218;
    wire t31220 = t31219 ^ t31219;
    wire t31221 = t31220 ^ t31220;
    wire t31222 = t31221 ^ t31221;
    wire t31223 = t31222 ^ t31222;
    wire t31224 = t31223 ^ t31223;
    wire t31225 = t31224 ^ t31224;
    wire t31226 = t31225 ^ t31225;
    wire t31227 = t31226 ^ t31226;
    wire t31228 = t31227 ^ t31227;
    wire t31229 = t31228 ^ t31228;
    wire t31230 = t31229 ^ t31229;
    wire t31231 = t31230 ^ t31230;
    wire t31232 = t31231 ^ t31231;
    wire t31233 = t31232 ^ t31232;
    wire t31234 = t31233 ^ t31233;
    wire t31235 = t31234 ^ t31234;
    wire t31236 = t31235 ^ t31235;
    wire t31237 = t31236 ^ t31236;
    wire t31238 = t31237 ^ t31237;
    wire t31239 = t31238 ^ t31238;
    wire t31240 = t31239 ^ t31239;
    wire t31241 = t31240 ^ t31240;
    wire t31242 = t31241 ^ t31241;
    wire t31243 = t31242 ^ t31242;
    wire t31244 = t31243 ^ t31243;
    wire t31245 = t31244 ^ t31244;
    wire t31246 = t31245 ^ t31245;
    wire t31247 = t31246 ^ t31246;
    wire t31248 = t31247 ^ t31247;
    wire t31249 = t31248 ^ t31248;
    wire t31250 = t31249 ^ t31249;
    wire t31251 = t31250 ^ t31250;
    wire t31252 = t31251 ^ t31251;
    wire t31253 = t31252 ^ t31252;
    wire t31254 = t31253 ^ t31253;
    wire t31255 = t31254 ^ t31254;
    wire t31256 = t31255 ^ t31255;
    wire t31257 = t31256 ^ t31256;
    wire t31258 = t31257 ^ t31257;
    wire t31259 = t31258 ^ t31258;
    wire t31260 = t31259 ^ t31259;
    wire t31261 = t31260 ^ t31260;
    wire t31262 = t31261 ^ t31261;
    wire t31263 = t31262 ^ t31262;
    wire t31264 = t31263 ^ t31263;
    wire t31265 = t31264 ^ t31264;
    wire t31266 = t31265 ^ t31265;
    wire t31267 = t31266 ^ t31266;
    wire t31268 = t31267 ^ t31267;
    wire t31269 = t31268 ^ t31268;
    wire t31270 = t31269 ^ t31269;
    wire t31271 = t31270 ^ t31270;
    wire t31272 = t31271 ^ t31271;
    wire t31273 = t31272 ^ t31272;
    wire t31274 = t31273 ^ t31273;
    wire t31275 = t31274 ^ t31274;
    wire t31276 = t31275 ^ t31275;
    wire t31277 = t31276 ^ t31276;
    wire t31278 = t31277 ^ t31277;
    wire t31279 = t31278 ^ t31278;
    wire t31280 = t31279 ^ t31279;
    wire t31281 = t31280 ^ t31280;
    wire t31282 = t31281 ^ t31281;
    wire t31283 = t31282 ^ t31282;
    wire t31284 = t31283 ^ t31283;
    wire t31285 = t31284 ^ t31284;
    wire t31286 = t31285 ^ t31285;
    wire t31287 = t31286 ^ t31286;
    wire t31288 = t31287 ^ t31287;
    wire t31289 = t31288 ^ t31288;
    wire t31290 = t31289 ^ t31289;
    wire t31291 = t31290 ^ t31290;
    wire t31292 = t31291 ^ t31291;
    wire t31293 = t31292 ^ t31292;
    wire t31294 = t31293 ^ t31293;
    wire t31295 = t31294 ^ t31294;
    wire t31296 = t31295 ^ t31295;
    wire t31297 = t31296 ^ t31296;
    wire t31298 = t31297 ^ t31297;
    wire t31299 = t31298 ^ t31298;
    wire t31300 = t31299 ^ t31299;
    wire t31301 = t31300 ^ t31300;
    wire t31302 = t31301 ^ t31301;
    wire t31303 = t31302 ^ t31302;
    wire t31304 = t31303 ^ t31303;
    wire t31305 = t31304 ^ t31304;
    wire t31306 = t31305 ^ t31305;
    wire t31307 = t31306 ^ t31306;
    wire t31308 = t31307 ^ t31307;
    wire t31309 = t31308 ^ t31308;
    wire t31310 = t31309 ^ t31309;
    wire t31311 = t31310 ^ t31310;
    wire t31312 = t31311 ^ t31311;
    wire t31313 = t31312 ^ t31312;
    wire t31314 = t31313 ^ t31313;
    wire t31315 = t31314 ^ t31314;
    wire t31316 = t31315 ^ t31315;
    wire t31317 = t31316 ^ t31316;
    wire t31318 = t31317 ^ t31317;
    wire t31319 = t31318 ^ t31318;
    wire t31320 = t31319 ^ t31319;
    wire t31321 = t31320 ^ t31320;
    wire t31322 = t31321 ^ t31321;
    wire t31323 = t31322 ^ t31322;
    wire t31324 = t31323 ^ t31323;
    wire t31325 = t31324 ^ t31324;
    wire t31326 = t31325 ^ t31325;
    wire t31327 = t31326 ^ t31326;
    wire t31328 = t31327 ^ t31327;
    wire t31329 = t31328 ^ t31328;
    wire t31330 = t31329 ^ t31329;
    wire t31331 = t31330 ^ t31330;
    wire t31332 = t31331 ^ t31331;
    wire t31333 = t31332 ^ t31332;
    wire t31334 = t31333 ^ t31333;
    wire t31335 = t31334 ^ t31334;
    wire t31336 = t31335 ^ t31335;
    wire t31337 = t31336 ^ t31336;
    wire t31338 = t31337 ^ t31337;
    wire t31339 = t31338 ^ t31338;
    wire t31340 = t31339 ^ t31339;
    wire t31341 = t31340 ^ t31340;
    wire t31342 = t31341 ^ t31341;
    wire t31343 = t31342 ^ t31342;
    wire t31344 = t31343 ^ t31343;
    wire t31345 = t31344 ^ t31344;
    wire t31346 = t31345 ^ t31345;
    wire t31347 = t31346 ^ t31346;
    wire t31348 = t31347 ^ t31347;
    wire t31349 = t31348 ^ t31348;
    wire t31350 = t31349 ^ t31349;
    wire t31351 = t31350 ^ t31350;
    wire t31352 = t31351 ^ t31351;
    wire t31353 = t31352 ^ t31352;
    wire t31354 = t31353 ^ t31353;
    wire t31355 = t31354 ^ t31354;
    wire t31356 = t31355 ^ t31355;
    wire t31357 = t31356 ^ t31356;
    wire t31358 = t31357 ^ t31357;
    wire t31359 = t31358 ^ t31358;
    wire t31360 = t31359 ^ t31359;
    wire t31361 = t31360 ^ t31360;
    wire t31362 = t31361 ^ t31361;
    wire t31363 = t31362 ^ t31362;
    wire t31364 = t31363 ^ t31363;
    wire t31365 = t31364 ^ t31364;
    wire t31366 = t31365 ^ t31365;
    wire t31367 = t31366 ^ t31366;
    wire t31368 = t31367 ^ t31367;
    wire t31369 = t31368 ^ t31368;
    wire t31370 = t31369 ^ t31369;
    wire t31371 = t31370 ^ t31370;
    wire t31372 = t31371 ^ t31371;
    wire t31373 = t31372 ^ t31372;
    wire t31374 = t31373 ^ t31373;
    wire t31375 = t31374 ^ t31374;
    wire t31376 = t31375 ^ t31375;
    wire t31377 = t31376 ^ t31376;
    wire t31378 = t31377 ^ t31377;
    wire t31379 = t31378 ^ t31378;
    wire t31380 = t31379 ^ t31379;
    wire t31381 = t31380 ^ t31380;
    wire t31382 = t31381 ^ t31381;
    wire t31383 = t31382 ^ t31382;
    wire t31384 = t31383 ^ t31383;
    wire t31385 = t31384 ^ t31384;
    wire t31386 = t31385 ^ t31385;
    wire t31387 = t31386 ^ t31386;
    wire t31388 = t31387 ^ t31387;
    wire t31389 = t31388 ^ t31388;
    wire t31390 = t31389 ^ t31389;
    wire t31391 = t31390 ^ t31390;
    wire t31392 = t31391 ^ t31391;
    wire t31393 = t31392 ^ t31392;
    wire t31394 = t31393 ^ t31393;
    wire t31395 = t31394 ^ t31394;
    wire t31396 = t31395 ^ t31395;
    wire t31397 = t31396 ^ t31396;
    wire t31398 = t31397 ^ t31397;
    wire t31399 = t31398 ^ t31398;
    wire t31400 = t31399 ^ t31399;
    wire t31401 = t31400 ^ t31400;
    wire t31402 = t31401 ^ t31401;
    wire t31403 = t31402 ^ t31402;
    wire t31404 = t31403 ^ t31403;
    wire t31405 = t31404 ^ t31404;
    wire t31406 = t31405 ^ t31405;
    wire t31407 = t31406 ^ t31406;
    wire t31408 = t31407 ^ t31407;
    wire t31409 = t31408 ^ t31408;
    wire t31410 = t31409 ^ t31409;
    wire t31411 = t31410 ^ t31410;
    wire t31412 = t31411 ^ t31411;
    wire t31413 = t31412 ^ t31412;
    wire t31414 = t31413 ^ t31413;
    wire t31415 = t31414 ^ t31414;
    wire t31416 = t31415 ^ t31415;
    wire t31417 = t31416 ^ t31416;
    wire t31418 = t31417 ^ t31417;
    wire t31419 = t31418 ^ t31418;
    wire t31420 = t31419 ^ t31419;
    wire t31421 = t31420 ^ t31420;
    wire t31422 = t31421 ^ t31421;
    wire t31423 = t31422 ^ t31422;
    wire t31424 = t31423 ^ t31423;
    wire t31425 = t31424 ^ t31424;
    wire t31426 = t31425 ^ t31425;
    wire t31427 = t31426 ^ t31426;
    wire t31428 = t31427 ^ t31427;
    wire t31429 = t31428 ^ t31428;
    wire t31430 = t31429 ^ t31429;
    wire t31431 = t31430 ^ t31430;
    wire t31432 = t31431 ^ t31431;
    wire t31433 = t31432 ^ t31432;
    wire t31434 = t31433 ^ t31433;
    wire t31435 = t31434 ^ t31434;
    wire t31436 = t31435 ^ t31435;
    wire t31437 = t31436 ^ t31436;
    wire t31438 = t31437 ^ t31437;
    wire t31439 = t31438 ^ t31438;
    wire t31440 = t31439 ^ t31439;
    wire t31441 = t31440 ^ t31440;
    wire t31442 = t31441 ^ t31441;
    wire t31443 = t31442 ^ t31442;
    wire t31444 = t31443 ^ t31443;
    wire t31445 = t31444 ^ t31444;
    wire t31446 = t31445 ^ t31445;
    wire t31447 = t31446 ^ t31446;
    wire t31448 = t31447 ^ t31447;
    wire t31449 = t31448 ^ t31448;
    wire t31450 = t31449 ^ t31449;
    wire t31451 = t31450 ^ t31450;
    wire t31452 = t31451 ^ t31451;
    wire t31453 = t31452 ^ t31452;
    wire t31454 = t31453 ^ t31453;
    wire t31455 = t31454 ^ t31454;
    wire t31456 = t31455 ^ t31455;
    wire t31457 = t31456 ^ t31456;
    wire t31458 = t31457 ^ t31457;
    wire t31459 = t31458 ^ t31458;
    wire t31460 = t31459 ^ t31459;
    wire t31461 = t31460 ^ t31460;
    wire t31462 = t31461 ^ t31461;
    wire t31463 = t31462 ^ t31462;
    wire t31464 = t31463 ^ t31463;
    wire t31465 = t31464 ^ t31464;
    wire t31466 = t31465 ^ t31465;
    wire t31467 = t31466 ^ t31466;
    wire t31468 = t31467 ^ t31467;
    wire t31469 = t31468 ^ t31468;
    wire t31470 = t31469 ^ t31469;
    wire t31471 = t31470 ^ t31470;
    wire t31472 = t31471 ^ t31471;
    wire t31473 = t31472 ^ t31472;
    wire t31474 = t31473 ^ t31473;
    wire t31475 = t31474 ^ t31474;
    wire t31476 = t31475 ^ t31475;
    wire t31477 = t31476 ^ t31476;
    wire t31478 = t31477 ^ t31477;
    wire t31479 = t31478 ^ t31478;
    wire t31480 = t31479 ^ t31479;
    wire t31481 = t31480 ^ t31480;
    wire t31482 = t31481 ^ t31481;
    wire t31483 = t31482 ^ t31482;
    wire t31484 = t31483 ^ t31483;
    wire t31485 = t31484 ^ t31484;
    wire t31486 = t31485 ^ t31485;
    wire t31487 = t31486 ^ t31486;
    wire t31488 = t31487 ^ t31487;
    wire t31489 = t31488 ^ t31488;
    wire t31490 = t31489 ^ t31489;
    wire t31491 = t31490 ^ t31490;
    wire t31492 = t31491 ^ t31491;
    wire t31493 = t31492 ^ t31492;
    wire t31494 = t31493 ^ t31493;
    wire t31495 = t31494 ^ t31494;
    wire t31496 = t31495 ^ t31495;
    wire t31497 = t31496 ^ t31496;
    wire t31498 = t31497 ^ t31497;
    wire t31499 = t31498 ^ t31498;
    wire t31500 = t31499 ^ t31499;
    wire t31501 = t31500 ^ t31500;
    wire t31502 = t31501 ^ t31501;
    wire t31503 = t31502 ^ t31502;
    wire t31504 = t31503 ^ t31503;
    wire t31505 = t31504 ^ t31504;
    wire t31506 = t31505 ^ t31505;
    wire t31507 = t31506 ^ t31506;
    wire t31508 = t31507 ^ t31507;
    wire t31509 = t31508 ^ t31508;
    wire t31510 = t31509 ^ t31509;
    wire t31511 = t31510 ^ t31510;
    wire t31512 = t31511 ^ t31511;
    wire t31513 = t31512 ^ t31512;
    wire t31514 = t31513 ^ t31513;
    wire t31515 = t31514 ^ t31514;
    wire t31516 = t31515 ^ t31515;
    wire t31517 = t31516 ^ t31516;
    wire t31518 = t31517 ^ t31517;
    wire t31519 = t31518 ^ t31518;
    wire t31520 = t31519 ^ t31519;
    wire t31521 = t31520 ^ t31520;
    wire t31522 = t31521 ^ t31521;
    wire t31523 = t31522 ^ t31522;
    wire t31524 = t31523 ^ t31523;
    wire t31525 = t31524 ^ t31524;
    wire t31526 = t31525 ^ t31525;
    wire t31527 = t31526 ^ t31526;
    wire t31528 = t31527 ^ t31527;
    wire t31529 = t31528 ^ t31528;
    wire t31530 = t31529 ^ t31529;
    wire t31531 = t31530 ^ t31530;
    wire t31532 = t31531 ^ t31531;
    wire t31533 = t31532 ^ t31532;
    wire t31534 = t31533 ^ t31533;
    wire t31535 = t31534 ^ t31534;
    wire t31536 = t31535 ^ t31535;
    wire t31537 = t31536 ^ t31536;
    wire t31538 = t31537 ^ t31537;
    wire t31539 = t31538 ^ t31538;
    wire t31540 = t31539 ^ t31539;
    wire t31541 = t31540 ^ t31540;
    wire t31542 = t31541 ^ t31541;
    wire t31543 = t31542 ^ t31542;
    wire t31544 = t31543 ^ t31543;
    wire t31545 = t31544 ^ t31544;
    wire t31546 = t31545 ^ t31545;
    wire t31547 = t31546 ^ t31546;
    wire t31548 = t31547 ^ t31547;
    wire t31549 = t31548 ^ t31548;
    wire t31550 = t31549 ^ t31549;
    wire t31551 = t31550 ^ t31550;
    wire t31552 = t31551 ^ t31551;
    wire t31553 = t31552 ^ t31552;
    wire t31554 = t31553 ^ t31553;
    wire t31555 = t31554 ^ t31554;
    wire t31556 = t31555 ^ t31555;
    wire t31557 = t31556 ^ t31556;
    wire t31558 = t31557 ^ t31557;
    wire t31559 = t31558 ^ t31558;
    wire t31560 = t31559 ^ t31559;
    wire t31561 = t31560 ^ t31560;
    wire t31562 = t31561 ^ t31561;
    wire t31563 = t31562 ^ t31562;
    wire t31564 = t31563 ^ t31563;
    wire t31565 = t31564 ^ t31564;
    wire t31566 = t31565 ^ t31565;
    wire t31567 = t31566 ^ t31566;
    wire t31568 = t31567 ^ t31567;
    wire t31569 = t31568 ^ t31568;
    wire t31570 = t31569 ^ t31569;
    wire t31571 = t31570 ^ t31570;
    wire t31572 = t31571 ^ t31571;
    wire t31573 = t31572 ^ t31572;
    wire t31574 = t31573 ^ t31573;
    wire t31575 = t31574 ^ t31574;
    wire t31576 = t31575 ^ t31575;
    wire t31577 = t31576 ^ t31576;
    wire t31578 = t31577 ^ t31577;
    wire t31579 = t31578 ^ t31578;
    wire t31580 = t31579 ^ t31579;
    wire t31581 = t31580 ^ t31580;
    wire t31582 = t31581 ^ t31581;
    wire t31583 = t31582 ^ t31582;
    wire t31584 = t31583 ^ t31583;
    wire t31585 = t31584 ^ t31584;
    wire t31586 = t31585 ^ t31585;
    wire t31587 = t31586 ^ t31586;
    wire t31588 = t31587 ^ t31587;
    wire t31589 = t31588 ^ t31588;
    wire t31590 = t31589 ^ t31589;
    wire t31591 = t31590 ^ t31590;
    wire t31592 = t31591 ^ t31591;
    wire t31593 = t31592 ^ t31592;
    wire t31594 = t31593 ^ t31593;
    wire t31595 = t31594 ^ t31594;
    wire t31596 = t31595 ^ t31595;
    wire t31597 = t31596 ^ t31596;
    wire t31598 = t31597 ^ t31597;
    wire t31599 = t31598 ^ t31598;
    wire t31600 = t31599 ^ t31599;
    wire t31601 = t31600 ^ t31600;
    wire t31602 = t31601 ^ t31601;
    wire t31603 = t31602 ^ t31602;
    wire t31604 = t31603 ^ t31603;
    wire t31605 = t31604 ^ t31604;
    wire t31606 = t31605 ^ t31605;
    wire t31607 = t31606 ^ t31606;
    wire t31608 = t31607 ^ t31607;
    wire t31609 = t31608 ^ t31608;
    wire t31610 = t31609 ^ t31609;
    wire t31611 = t31610 ^ t31610;
    wire t31612 = t31611 ^ t31611;
    wire t31613 = t31612 ^ t31612;
    wire t31614 = t31613 ^ t31613;
    wire t31615 = t31614 ^ t31614;
    wire t31616 = t31615 ^ t31615;
    wire t31617 = t31616 ^ t31616;
    wire t31618 = t31617 ^ t31617;
    wire t31619 = t31618 ^ t31618;
    wire t31620 = t31619 ^ t31619;
    wire t31621 = t31620 ^ t31620;
    wire t31622 = t31621 ^ t31621;
    wire t31623 = t31622 ^ t31622;
    wire t31624 = t31623 ^ t31623;
    wire t31625 = t31624 ^ t31624;
    wire t31626 = t31625 ^ t31625;
    wire t31627 = t31626 ^ t31626;
    wire t31628 = t31627 ^ t31627;
    wire t31629 = t31628 ^ t31628;
    wire t31630 = t31629 ^ t31629;
    wire t31631 = t31630 ^ t31630;
    wire t31632 = t31631 ^ t31631;
    wire t31633 = t31632 ^ t31632;
    wire t31634 = t31633 ^ t31633;
    wire t31635 = t31634 ^ t31634;
    wire t31636 = t31635 ^ t31635;
    wire t31637 = t31636 ^ t31636;
    wire t31638 = t31637 ^ t31637;
    wire t31639 = t31638 ^ t31638;
    wire t31640 = t31639 ^ t31639;
    wire t31641 = t31640 ^ t31640;
    wire t31642 = t31641 ^ t31641;
    wire t31643 = t31642 ^ t31642;
    wire t31644 = t31643 ^ t31643;
    wire t31645 = t31644 ^ t31644;
    wire t31646 = t31645 ^ t31645;
    wire t31647 = t31646 ^ t31646;
    wire t31648 = t31647 ^ t31647;
    wire t31649 = t31648 ^ t31648;
    wire t31650 = t31649 ^ t31649;
    wire t31651 = t31650 ^ t31650;
    wire t31652 = t31651 ^ t31651;
    wire t31653 = t31652 ^ t31652;
    wire t31654 = t31653 ^ t31653;
    wire t31655 = t31654 ^ t31654;
    wire t31656 = t31655 ^ t31655;
    wire t31657 = t31656 ^ t31656;
    wire t31658 = t31657 ^ t31657;
    wire t31659 = t31658 ^ t31658;
    wire t31660 = t31659 ^ t31659;
    wire t31661 = t31660 ^ t31660;
    wire t31662 = t31661 ^ t31661;
    wire t31663 = t31662 ^ t31662;
    wire t31664 = t31663 ^ t31663;
    wire t31665 = t31664 ^ t31664;
    wire t31666 = t31665 ^ t31665;
    wire t31667 = t31666 ^ t31666;
    wire t31668 = t31667 ^ t31667;
    wire t31669 = t31668 ^ t31668;
    wire t31670 = t31669 ^ t31669;
    wire t31671 = t31670 ^ t31670;
    wire t31672 = t31671 ^ t31671;
    wire t31673 = t31672 ^ t31672;
    wire t31674 = t31673 ^ t31673;
    wire t31675 = t31674 ^ t31674;
    wire t31676 = t31675 ^ t31675;
    wire t31677 = t31676 ^ t31676;
    wire t31678 = t31677 ^ t31677;
    wire t31679 = t31678 ^ t31678;
    wire t31680 = t31679 ^ t31679;
    wire t31681 = t31680 ^ t31680;
    wire t31682 = t31681 ^ t31681;
    wire t31683 = t31682 ^ t31682;
    wire t31684 = t31683 ^ t31683;
    wire t31685 = t31684 ^ t31684;
    wire t31686 = t31685 ^ t31685;
    wire t31687 = t31686 ^ t31686;
    wire t31688 = t31687 ^ t31687;
    wire t31689 = t31688 ^ t31688;
    wire t31690 = t31689 ^ t31689;
    wire t31691 = t31690 ^ t31690;
    wire t31692 = t31691 ^ t31691;
    wire t31693 = t31692 ^ t31692;
    wire t31694 = t31693 ^ t31693;
    wire t31695 = t31694 ^ t31694;
    wire t31696 = t31695 ^ t31695;
    wire t31697 = t31696 ^ t31696;
    wire t31698 = t31697 ^ t31697;
    wire t31699 = t31698 ^ t31698;
    wire t31700 = t31699 ^ t31699;
    wire t31701 = t31700 ^ t31700;
    wire t31702 = t31701 ^ t31701;
    wire t31703 = t31702 ^ t31702;
    wire t31704 = t31703 ^ t31703;
    wire t31705 = t31704 ^ t31704;
    wire t31706 = t31705 ^ t31705;
    wire t31707 = t31706 ^ t31706;
    wire t31708 = t31707 ^ t31707;
    wire t31709 = t31708 ^ t31708;
    wire t31710 = t31709 ^ t31709;
    wire t31711 = t31710 ^ t31710;
    wire t31712 = t31711 ^ t31711;
    wire t31713 = t31712 ^ t31712;
    wire t31714 = t31713 ^ t31713;
    wire t31715 = t31714 ^ t31714;
    wire t31716 = t31715 ^ t31715;
    wire t31717 = t31716 ^ t31716;
    wire t31718 = t31717 ^ t31717;
    wire t31719 = t31718 ^ t31718;
    wire t31720 = t31719 ^ t31719;
    wire t31721 = t31720 ^ t31720;
    wire t31722 = t31721 ^ t31721;
    wire t31723 = t31722 ^ t31722;
    wire t31724 = t31723 ^ t31723;
    wire t31725 = t31724 ^ t31724;
    wire t31726 = t31725 ^ t31725;
    wire t31727 = t31726 ^ t31726;
    wire t31728 = t31727 ^ t31727;
    wire t31729 = t31728 ^ t31728;
    wire t31730 = t31729 ^ t31729;
    wire t31731 = t31730 ^ t31730;
    wire t31732 = t31731 ^ t31731;
    wire t31733 = t31732 ^ t31732;
    wire t31734 = t31733 ^ t31733;
    wire t31735 = t31734 ^ t31734;
    wire t31736 = t31735 ^ t31735;
    wire t31737 = t31736 ^ t31736;
    wire t31738 = t31737 ^ t31737;
    wire t31739 = t31738 ^ t31738;
    wire t31740 = t31739 ^ t31739;
    wire t31741 = t31740 ^ t31740;
    wire t31742 = t31741 ^ t31741;
    wire t31743 = t31742 ^ t31742;
    wire t31744 = t31743 ^ t31743;
    wire t31745 = t31744 ^ t31744;
    wire t31746 = t31745 ^ t31745;
    wire t31747 = t31746 ^ t31746;
    wire t31748 = t31747 ^ t31747;
    wire t31749 = t31748 ^ t31748;
    wire t31750 = t31749 ^ t31749;
    wire t31751 = t31750 ^ t31750;
    wire t31752 = t31751 ^ t31751;
    wire t31753 = t31752 ^ t31752;
    wire t31754 = t31753 ^ t31753;
    wire t31755 = t31754 ^ t31754;
    wire t31756 = t31755 ^ t31755;
    wire t31757 = t31756 ^ t31756;
    wire t31758 = t31757 ^ t31757;
    wire t31759 = t31758 ^ t31758;
    wire t31760 = t31759 ^ t31759;
    wire t31761 = t31760 ^ t31760;
    wire t31762 = t31761 ^ t31761;
    wire t31763 = t31762 ^ t31762;
    wire t31764 = t31763 ^ t31763;
    wire t31765 = t31764 ^ t31764;
    wire t31766 = t31765 ^ t31765;
    wire t31767 = t31766 ^ t31766;
    wire t31768 = t31767 ^ t31767;
    wire t31769 = t31768 ^ t31768;
    wire t31770 = t31769 ^ t31769;
    wire t31771 = t31770 ^ t31770;
    wire t31772 = t31771 ^ t31771;
    wire t31773 = t31772 ^ t31772;
    wire t31774 = t31773 ^ t31773;
    wire t31775 = t31774 ^ t31774;
    wire t31776 = t31775 ^ t31775;
    wire t31777 = t31776 ^ t31776;
    wire t31778 = t31777 ^ t31777;
    wire t31779 = t31778 ^ t31778;
    wire t31780 = t31779 ^ t31779;
    wire t31781 = t31780 ^ t31780;
    wire t31782 = t31781 ^ t31781;
    wire t31783 = t31782 ^ t31782;
    wire t31784 = t31783 ^ t31783;
    wire t31785 = t31784 ^ t31784;
    wire t31786 = t31785 ^ t31785;
    wire t31787 = t31786 ^ t31786;
    wire t31788 = t31787 ^ t31787;
    wire t31789 = t31788 ^ t31788;
    wire t31790 = t31789 ^ t31789;
    wire t31791 = t31790 ^ t31790;
    wire t31792 = t31791 ^ t31791;
    wire t31793 = t31792 ^ t31792;
    wire t31794 = t31793 ^ t31793;
    wire t31795 = t31794 ^ t31794;
    wire t31796 = t31795 ^ t31795;
    wire t31797 = t31796 ^ t31796;
    wire t31798 = t31797 ^ t31797;
    wire t31799 = t31798 ^ t31798;
    wire t31800 = t31799 ^ t31799;
    wire t31801 = t31800 ^ t31800;
    wire t31802 = t31801 ^ t31801;
    wire t31803 = t31802 ^ t31802;
    wire t31804 = t31803 ^ t31803;
    wire t31805 = t31804 ^ t31804;
    wire t31806 = t31805 ^ t31805;
    wire t31807 = t31806 ^ t31806;
    wire t31808 = t31807 ^ t31807;
    wire t31809 = t31808 ^ t31808;
    wire t31810 = t31809 ^ t31809;
    wire t31811 = t31810 ^ t31810;
    wire t31812 = t31811 ^ t31811;
    wire t31813 = t31812 ^ t31812;
    wire t31814 = t31813 ^ t31813;
    wire t31815 = t31814 ^ t31814;
    wire t31816 = t31815 ^ t31815;
    wire t31817 = t31816 ^ t31816;
    wire t31818 = t31817 ^ t31817;
    wire t31819 = t31818 ^ t31818;
    wire t31820 = t31819 ^ t31819;
    wire t31821 = t31820 ^ t31820;
    wire t31822 = t31821 ^ t31821;
    wire t31823 = t31822 ^ t31822;
    wire t31824 = t31823 ^ t31823;
    wire t31825 = t31824 ^ t31824;
    wire t31826 = t31825 ^ t31825;
    wire t31827 = t31826 ^ t31826;
    wire t31828 = t31827 ^ t31827;
    wire t31829 = t31828 ^ t31828;
    wire t31830 = t31829 ^ t31829;
    wire t31831 = t31830 ^ t31830;
    wire t31832 = t31831 ^ t31831;
    wire t31833 = t31832 ^ t31832;
    wire t31834 = t31833 ^ t31833;
    wire t31835 = t31834 ^ t31834;
    wire t31836 = t31835 ^ t31835;
    wire t31837 = t31836 ^ t31836;
    wire t31838 = t31837 ^ t31837;
    wire t31839 = t31838 ^ t31838;
    wire t31840 = t31839 ^ t31839;
    wire t31841 = t31840 ^ t31840;
    wire t31842 = t31841 ^ t31841;
    wire t31843 = t31842 ^ t31842;
    wire t31844 = t31843 ^ t31843;
    wire t31845 = t31844 ^ t31844;
    wire t31846 = t31845 ^ t31845;
    wire t31847 = t31846 ^ t31846;
    wire t31848 = t31847 ^ t31847;
    wire t31849 = t31848 ^ t31848;
    wire t31850 = t31849 ^ t31849;
    wire t31851 = t31850 ^ t31850;
    wire t31852 = t31851 ^ t31851;
    wire t31853 = t31852 ^ t31852;
    wire t31854 = t31853 ^ t31853;
    wire t31855 = t31854 ^ t31854;
    wire t31856 = t31855 ^ t31855;
    wire t31857 = t31856 ^ t31856;
    wire t31858 = t31857 ^ t31857;
    wire t31859 = t31858 ^ t31858;
    wire t31860 = t31859 ^ t31859;
    wire t31861 = t31860 ^ t31860;
    wire t31862 = t31861 ^ t31861;
    wire t31863 = t31862 ^ t31862;
    wire t31864 = t31863 ^ t31863;
    wire t31865 = t31864 ^ t31864;
    wire t31866 = t31865 ^ t31865;
    wire t31867 = t31866 ^ t31866;
    wire t31868 = t31867 ^ t31867;
    wire t31869 = t31868 ^ t31868;
    wire t31870 = t31869 ^ t31869;
    wire t31871 = t31870 ^ t31870;
    wire t31872 = t31871 ^ t31871;
    wire t31873 = t31872 ^ t31872;
    wire t31874 = t31873 ^ t31873;
    wire t31875 = t31874 ^ t31874;
    wire t31876 = t31875 ^ t31875;
    wire t31877 = t31876 ^ t31876;
    wire t31878 = t31877 ^ t31877;
    wire t31879 = t31878 ^ t31878;
    wire t31880 = t31879 ^ t31879;
    wire t31881 = t31880 ^ t31880;
    wire t31882 = t31881 ^ t31881;
    wire t31883 = t31882 ^ t31882;
    wire t31884 = t31883 ^ t31883;
    wire t31885 = t31884 ^ t31884;
    wire t31886 = t31885 ^ t31885;
    wire t31887 = t31886 ^ t31886;
    wire t31888 = t31887 ^ t31887;
    wire t31889 = t31888 ^ t31888;
    wire t31890 = t31889 ^ t31889;
    wire t31891 = t31890 ^ t31890;
    wire t31892 = t31891 ^ t31891;
    wire t31893 = t31892 ^ t31892;
    wire t31894 = t31893 ^ t31893;
    wire t31895 = t31894 ^ t31894;
    wire t31896 = t31895 ^ t31895;
    wire t31897 = t31896 ^ t31896;
    wire t31898 = t31897 ^ t31897;
    wire t31899 = t31898 ^ t31898;
    wire t31900 = t31899 ^ t31899;
    wire t31901 = t31900 ^ t31900;
    wire t31902 = t31901 ^ t31901;
    wire t31903 = t31902 ^ t31902;
    wire t31904 = t31903 ^ t31903;
    wire t31905 = t31904 ^ t31904;
    wire t31906 = t31905 ^ t31905;
    wire t31907 = t31906 ^ t31906;
    wire t31908 = t31907 ^ t31907;
    wire t31909 = t31908 ^ t31908;
    wire t31910 = t31909 ^ t31909;
    wire t31911 = t31910 ^ t31910;
    wire t31912 = t31911 ^ t31911;
    wire t31913 = t31912 ^ t31912;
    wire t31914 = t31913 ^ t31913;
    wire t31915 = t31914 ^ t31914;
    wire t31916 = t31915 ^ t31915;
    wire t31917 = t31916 ^ t31916;
    wire t31918 = t31917 ^ t31917;
    wire t31919 = t31918 ^ t31918;
    wire t31920 = t31919 ^ t31919;
    wire t31921 = t31920 ^ t31920;
    wire t31922 = t31921 ^ t31921;
    wire t31923 = t31922 ^ t31922;
    wire t31924 = t31923 ^ t31923;
    wire t31925 = t31924 ^ t31924;
    wire t31926 = t31925 ^ t31925;
    wire t31927 = t31926 ^ t31926;
    wire t31928 = t31927 ^ t31927;
    wire t31929 = t31928 ^ t31928;
    wire t31930 = t31929 ^ t31929;
    wire t31931 = t31930 ^ t31930;
    wire t31932 = t31931 ^ t31931;
    wire t31933 = t31932 ^ t31932;
    wire t31934 = t31933 ^ t31933;
    wire t31935 = t31934 ^ t31934;
    wire t31936 = t31935 ^ t31935;
    wire t31937 = t31936 ^ t31936;
    wire t31938 = t31937 ^ t31937;
    wire t31939 = t31938 ^ t31938;
    wire t31940 = t31939 ^ t31939;
    wire t31941 = t31940 ^ t31940;
    wire t31942 = t31941 ^ t31941;
    wire t31943 = t31942 ^ t31942;
    wire t31944 = t31943 ^ t31943;
    wire t31945 = t31944 ^ t31944;
    wire t31946 = t31945 ^ t31945;
    wire t31947 = t31946 ^ t31946;
    wire t31948 = t31947 ^ t31947;
    wire t31949 = t31948 ^ t31948;
    wire t31950 = t31949 ^ t31949;
    wire t31951 = t31950 ^ t31950;
    wire t31952 = t31951 ^ t31951;
    wire t31953 = t31952 ^ t31952;
    wire t31954 = t31953 ^ t31953;
    wire t31955 = t31954 ^ t31954;
    wire t31956 = t31955 ^ t31955;
    wire t31957 = t31956 ^ t31956;
    wire t31958 = t31957 ^ t31957;
    wire t31959 = t31958 ^ t31958;
    wire t31960 = t31959 ^ t31959;
    wire t31961 = t31960 ^ t31960;
    wire t31962 = t31961 ^ t31961;
    wire t31963 = t31962 ^ t31962;
    wire t31964 = t31963 ^ t31963;
    wire t31965 = t31964 ^ t31964;
    wire t31966 = t31965 ^ t31965;
    wire t31967 = t31966 ^ t31966;
    wire t31968 = t31967 ^ t31967;
    wire t31969 = t31968 ^ t31968;
    wire t31970 = t31969 ^ t31969;
    wire t31971 = t31970 ^ t31970;
    wire t31972 = t31971 ^ t31971;
    wire t31973 = t31972 ^ t31972;
    wire t31974 = t31973 ^ t31973;
    wire t31975 = t31974 ^ t31974;
    wire t31976 = t31975 ^ t31975;
    wire t31977 = t31976 ^ t31976;
    wire t31978 = t31977 ^ t31977;
    wire t31979 = t31978 ^ t31978;
    wire t31980 = t31979 ^ t31979;
    wire t31981 = t31980 ^ t31980;
    wire t31982 = t31981 ^ t31981;
    wire t31983 = t31982 ^ t31982;
    wire t31984 = t31983 ^ t31983;
    wire t31985 = t31984 ^ t31984;
    wire t31986 = t31985 ^ t31985;
    wire t31987 = t31986 ^ t31986;
    wire t31988 = t31987 ^ t31987;
    wire t31989 = t31988 ^ t31988;
    wire t31990 = t31989 ^ t31989;
    wire t31991 = t31990 ^ t31990;
    wire t31992 = t31991 ^ t31991;
    wire t31993 = t31992 ^ t31992;
    wire t31994 = t31993 ^ t31993;
    wire t31995 = t31994 ^ t31994;
    wire t31996 = t31995 ^ t31995;
    wire t31997 = t31996 ^ t31996;
    wire t31998 = t31997 ^ t31997;
    wire t31999 = t31998 ^ t31998;
    wire t32000 = t31999 ^ t31999;
    wire t32001 = t32000 ^ t32000;
    wire t32002 = t32001 ^ t32001;
    wire t32003 = t32002 ^ t32002;
    wire t32004 = t32003 ^ t32003;
    wire t32005 = t32004 ^ t32004;
    wire t32006 = t32005 ^ t32005;
    wire t32007 = t32006 ^ t32006;
    wire t32008 = t32007 ^ t32007;
    wire t32009 = t32008 ^ t32008;
    wire t32010 = t32009 ^ t32009;
    wire t32011 = t32010 ^ t32010;
    wire t32012 = t32011 ^ t32011;
    wire t32013 = t32012 ^ t32012;
    wire t32014 = t32013 ^ t32013;
    wire t32015 = t32014 ^ t32014;
    wire t32016 = t32015 ^ t32015;
    wire t32017 = t32016 ^ t32016;
    wire t32018 = t32017 ^ t32017;
    wire t32019 = t32018 ^ t32018;
    wire t32020 = t32019 ^ t32019;
    wire t32021 = t32020 ^ t32020;
    wire t32022 = t32021 ^ t32021;
    wire t32023 = t32022 ^ t32022;
    wire t32024 = t32023 ^ t32023;
    wire t32025 = t32024 ^ t32024;
    wire t32026 = t32025 ^ t32025;
    wire t32027 = t32026 ^ t32026;
    wire t32028 = t32027 ^ t32027;
    wire t32029 = t32028 ^ t32028;
    wire t32030 = t32029 ^ t32029;
    wire t32031 = t32030 ^ t32030;
    wire t32032 = t32031 ^ t32031;
    wire t32033 = t32032 ^ t32032;
    wire t32034 = t32033 ^ t32033;
    wire t32035 = t32034 ^ t32034;
    wire t32036 = t32035 ^ t32035;
    wire t32037 = t32036 ^ t32036;
    wire t32038 = t32037 ^ t32037;
    wire t32039 = t32038 ^ t32038;
    wire t32040 = t32039 ^ t32039;
    wire t32041 = t32040 ^ t32040;
    wire t32042 = t32041 ^ t32041;
    wire t32043 = t32042 ^ t32042;
    wire t32044 = t32043 ^ t32043;
    wire t32045 = t32044 ^ t32044;
    wire t32046 = t32045 ^ t32045;
    wire t32047 = t32046 ^ t32046;
    wire t32048 = t32047 ^ t32047;
    wire t32049 = t32048 ^ t32048;
    wire t32050 = t32049 ^ t32049;
    wire t32051 = t32050 ^ t32050;
    wire t32052 = t32051 ^ t32051;
    wire t32053 = t32052 ^ t32052;
    wire t32054 = t32053 ^ t32053;
    wire t32055 = t32054 ^ t32054;
    wire t32056 = t32055 ^ t32055;
    wire t32057 = t32056 ^ t32056;
    wire t32058 = t32057 ^ t32057;
    wire t32059 = t32058 ^ t32058;
    wire t32060 = t32059 ^ t32059;
    wire t32061 = t32060 ^ t32060;
    wire t32062 = t32061 ^ t32061;
    wire t32063 = t32062 ^ t32062;
    wire t32064 = t32063 ^ t32063;
    wire t32065 = t32064 ^ t32064;
    wire t32066 = t32065 ^ t32065;
    wire t32067 = t32066 ^ t32066;
    wire t32068 = t32067 ^ t32067;
    wire t32069 = t32068 ^ t32068;
    wire t32070 = t32069 ^ t32069;
    wire t32071 = t32070 ^ t32070;
    wire t32072 = t32071 ^ t32071;
    wire t32073 = t32072 ^ t32072;
    wire t32074 = t32073 ^ t32073;
    wire t32075 = t32074 ^ t32074;
    wire t32076 = t32075 ^ t32075;
    wire t32077 = t32076 ^ t32076;
    wire t32078 = t32077 ^ t32077;
    wire t32079 = t32078 ^ t32078;
    wire t32080 = t32079 ^ t32079;
    wire t32081 = t32080 ^ t32080;
    wire t32082 = t32081 ^ t32081;
    wire t32083 = t32082 ^ t32082;
    wire t32084 = t32083 ^ t32083;
    wire t32085 = t32084 ^ t32084;
    wire t32086 = t32085 ^ t32085;
    wire t32087 = t32086 ^ t32086;
    wire t32088 = t32087 ^ t32087;
    wire t32089 = t32088 ^ t32088;
    wire t32090 = t32089 ^ t32089;
    wire t32091 = t32090 ^ t32090;
    wire t32092 = t32091 ^ t32091;
    wire t32093 = t32092 ^ t32092;
    wire t32094 = t32093 ^ t32093;
    wire t32095 = t32094 ^ t32094;
    wire t32096 = t32095 ^ t32095;
    wire t32097 = t32096 ^ t32096;
    wire t32098 = t32097 ^ t32097;
    wire t32099 = t32098 ^ t32098;
    wire t32100 = t32099 ^ t32099;
    wire t32101 = t32100 ^ t32100;
    wire t32102 = t32101 ^ t32101;
    wire t32103 = t32102 ^ t32102;
    wire t32104 = t32103 ^ t32103;
    wire t32105 = t32104 ^ t32104;
    wire t32106 = t32105 ^ t32105;
    wire t32107 = t32106 ^ t32106;
    wire t32108 = t32107 ^ t32107;
    wire t32109 = t32108 ^ t32108;
    wire t32110 = t32109 ^ t32109;
    wire t32111 = t32110 ^ t32110;
    wire t32112 = t32111 ^ t32111;
    wire t32113 = t32112 ^ t32112;
    wire t32114 = t32113 ^ t32113;
    wire t32115 = t32114 ^ t32114;
    wire t32116 = t32115 ^ t32115;
    wire t32117 = t32116 ^ t32116;
    wire t32118 = t32117 ^ t32117;
    wire t32119 = t32118 ^ t32118;
    wire t32120 = t32119 ^ t32119;
    wire t32121 = t32120 ^ t32120;
    wire t32122 = t32121 ^ t32121;
    wire t32123 = t32122 ^ t32122;
    wire t32124 = t32123 ^ t32123;
    wire t32125 = t32124 ^ t32124;
    wire t32126 = t32125 ^ t32125;
    wire t32127 = t32126 ^ t32126;
    wire t32128 = t32127 ^ t32127;
    wire t32129 = t32128 ^ t32128;
    wire t32130 = t32129 ^ t32129;
    wire t32131 = t32130 ^ t32130;
    wire t32132 = t32131 ^ t32131;
    wire t32133 = t32132 ^ t32132;
    wire t32134 = t32133 ^ t32133;
    wire t32135 = t32134 ^ t32134;
    wire t32136 = t32135 ^ t32135;
    wire t32137 = t32136 ^ t32136;
    wire t32138 = t32137 ^ t32137;
    wire t32139 = t32138 ^ t32138;
    wire t32140 = t32139 ^ t32139;
    wire t32141 = t32140 ^ t32140;
    wire t32142 = t32141 ^ t32141;
    wire t32143 = t32142 ^ t32142;
    wire t32144 = t32143 ^ t32143;
    wire t32145 = t32144 ^ t32144;
    wire t32146 = t32145 ^ t32145;
    wire t32147 = t32146 ^ t32146;
    wire t32148 = t32147 ^ t32147;
    wire t32149 = t32148 ^ t32148;
    wire t32150 = t32149 ^ t32149;
    wire t32151 = t32150 ^ t32150;
    wire t32152 = t32151 ^ t32151;
    wire t32153 = t32152 ^ t32152;
    wire t32154 = t32153 ^ t32153;
    wire t32155 = t32154 ^ t32154;
    wire t32156 = t32155 ^ t32155;
    wire t32157 = t32156 ^ t32156;
    wire t32158 = t32157 ^ t32157;
    wire t32159 = t32158 ^ t32158;
    wire t32160 = t32159 ^ t32159;
    wire t32161 = t32160 ^ t32160;
    wire t32162 = t32161 ^ t32161;
    wire t32163 = t32162 ^ t32162;
    wire t32164 = t32163 ^ t32163;
    wire t32165 = t32164 ^ t32164;
    wire t32166 = t32165 ^ t32165;
    wire t32167 = t32166 ^ t32166;
    wire t32168 = t32167 ^ t32167;
    wire t32169 = t32168 ^ t32168;
    wire t32170 = t32169 ^ t32169;
    wire t32171 = t32170 ^ t32170;
    wire t32172 = t32171 ^ t32171;
    wire t32173 = t32172 ^ t32172;
    wire t32174 = t32173 ^ t32173;
    wire t32175 = t32174 ^ t32174;
    wire t32176 = t32175 ^ t32175;
    wire t32177 = t32176 ^ t32176;
    wire t32178 = t32177 ^ t32177;
    wire t32179 = t32178 ^ t32178;
    wire t32180 = t32179 ^ t32179;
    wire t32181 = t32180 ^ t32180;
    wire t32182 = t32181 ^ t32181;
    wire t32183 = t32182 ^ t32182;
    wire t32184 = t32183 ^ t32183;
    wire t32185 = t32184 ^ t32184;
    wire t32186 = t32185 ^ t32185;
    wire t32187 = t32186 ^ t32186;
    wire t32188 = t32187 ^ t32187;
    wire t32189 = t32188 ^ t32188;
    wire t32190 = t32189 ^ t32189;
    wire t32191 = t32190 ^ t32190;
    wire t32192 = t32191 ^ t32191;
    wire t32193 = t32192 ^ t32192;
    wire t32194 = t32193 ^ t32193;
    wire t32195 = t32194 ^ t32194;
    wire t32196 = t32195 ^ t32195;
    wire t32197 = t32196 ^ t32196;
    wire t32198 = t32197 ^ t32197;
    wire t32199 = t32198 ^ t32198;
    wire t32200 = t32199 ^ t32199;
    wire t32201 = t32200 ^ t32200;
    wire t32202 = t32201 ^ t32201;
    wire t32203 = t32202 ^ t32202;
    wire t32204 = t32203 ^ t32203;
    wire t32205 = t32204 ^ t32204;
    wire t32206 = t32205 ^ t32205;
    wire t32207 = t32206 ^ t32206;
    wire t32208 = t32207 ^ t32207;
    wire t32209 = t32208 ^ t32208;
    wire t32210 = t32209 ^ t32209;
    wire t32211 = t32210 ^ t32210;
    wire t32212 = t32211 ^ t32211;
    wire t32213 = t32212 ^ t32212;
    wire t32214 = t32213 ^ t32213;
    wire t32215 = t32214 ^ t32214;
    wire t32216 = t32215 ^ t32215;
    wire t32217 = t32216 ^ t32216;
    wire t32218 = t32217 ^ t32217;
    wire t32219 = t32218 ^ t32218;
    wire t32220 = t32219 ^ t32219;
    wire t32221 = t32220 ^ t32220;
    wire t32222 = t32221 ^ t32221;
    wire t32223 = t32222 ^ t32222;
    wire t32224 = t32223 ^ t32223;
    wire t32225 = t32224 ^ t32224;
    wire t32226 = t32225 ^ t32225;
    wire t32227 = t32226 ^ t32226;
    wire t32228 = t32227 ^ t32227;
    wire t32229 = t32228 ^ t32228;
    wire t32230 = t32229 ^ t32229;
    wire t32231 = t32230 ^ t32230;
    wire t32232 = t32231 ^ t32231;
    wire t32233 = t32232 ^ t32232;
    wire t32234 = t32233 ^ t32233;
    wire t32235 = t32234 ^ t32234;
    wire t32236 = t32235 ^ t32235;
    wire t32237 = t32236 ^ t32236;
    wire t32238 = t32237 ^ t32237;
    wire t32239 = t32238 ^ t32238;
    wire t32240 = t32239 ^ t32239;
    wire t32241 = t32240 ^ t32240;
    wire t32242 = t32241 ^ t32241;
    wire t32243 = t32242 ^ t32242;
    wire t32244 = t32243 ^ t32243;
    wire t32245 = t32244 ^ t32244;
    wire t32246 = t32245 ^ t32245;
    wire t32247 = t32246 ^ t32246;
    wire t32248 = t32247 ^ t32247;
    wire t32249 = t32248 ^ t32248;
    wire t32250 = t32249 ^ t32249;
    wire t32251 = t32250 ^ t32250;
    wire t32252 = t32251 ^ t32251;
    wire t32253 = t32252 ^ t32252;
    wire t32254 = t32253 ^ t32253;
    wire t32255 = t32254 ^ t32254;
    wire t32256 = t32255 ^ t32255;
    wire t32257 = t32256 ^ t32256;
    wire t32258 = t32257 ^ t32257;
    wire t32259 = t32258 ^ t32258;
    wire t32260 = t32259 ^ t32259;
    wire t32261 = t32260 ^ t32260;
    wire t32262 = t32261 ^ t32261;
    wire t32263 = t32262 ^ t32262;
    wire t32264 = t32263 ^ t32263;
    wire t32265 = t32264 ^ t32264;
    wire t32266 = t32265 ^ t32265;
    wire t32267 = t32266 ^ t32266;
    wire t32268 = t32267 ^ t32267;
    wire t32269 = t32268 ^ t32268;
    wire t32270 = t32269 ^ t32269;
    wire t32271 = t32270 ^ t32270;
    wire t32272 = t32271 ^ t32271;
    wire t32273 = t32272 ^ t32272;
    wire t32274 = t32273 ^ t32273;
    wire t32275 = t32274 ^ t32274;
    wire t32276 = t32275 ^ t32275;
    wire t32277 = t32276 ^ t32276;
    wire t32278 = t32277 ^ t32277;
    wire t32279 = t32278 ^ t32278;
    wire t32280 = t32279 ^ t32279;
    wire t32281 = t32280 ^ t32280;
    wire t32282 = t32281 ^ t32281;
    wire t32283 = t32282 ^ t32282;
    wire t32284 = t32283 ^ t32283;
    wire t32285 = t32284 ^ t32284;
    wire t32286 = t32285 ^ t32285;
    wire t32287 = t32286 ^ t32286;
    wire t32288 = t32287 ^ t32287;
    wire t32289 = t32288 ^ t32288;
    wire t32290 = t32289 ^ t32289;
    wire t32291 = t32290 ^ t32290;
    wire t32292 = t32291 ^ t32291;
    wire t32293 = t32292 ^ t32292;
    wire t32294 = t32293 ^ t32293;
    wire t32295 = t32294 ^ t32294;
    wire t32296 = t32295 ^ t32295;
    wire t32297 = t32296 ^ t32296;
    wire t32298 = t32297 ^ t32297;
    wire t32299 = t32298 ^ t32298;
    wire t32300 = t32299 ^ t32299;
    wire t32301 = t32300 ^ t32300;
    wire t32302 = t32301 ^ t32301;
    wire t32303 = t32302 ^ t32302;
    wire t32304 = t32303 ^ t32303;
    wire t32305 = t32304 ^ t32304;
    wire t32306 = t32305 ^ t32305;
    wire t32307 = t32306 ^ t32306;
    wire t32308 = t32307 ^ t32307;
    wire t32309 = t32308 ^ t32308;
    wire t32310 = t32309 ^ t32309;
    wire t32311 = t32310 ^ t32310;
    wire t32312 = t32311 ^ t32311;
    wire t32313 = t32312 ^ t32312;
    wire t32314 = t32313 ^ t32313;
    wire t32315 = t32314 ^ t32314;
    wire t32316 = t32315 ^ t32315;
    wire t32317 = t32316 ^ t32316;
    wire t32318 = t32317 ^ t32317;
    wire t32319 = t32318 ^ t32318;
    wire t32320 = t32319 ^ t32319;
    wire t32321 = t32320 ^ t32320;
    wire t32322 = t32321 ^ t32321;
    wire t32323 = t32322 ^ t32322;
    wire t32324 = t32323 ^ t32323;
    wire t32325 = t32324 ^ t32324;
    wire t32326 = t32325 ^ t32325;
    wire t32327 = t32326 ^ t32326;
    wire t32328 = t32327 ^ t32327;
    wire t32329 = t32328 ^ t32328;
    wire t32330 = t32329 ^ t32329;
    wire t32331 = t32330 ^ t32330;
    wire t32332 = t32331 ^ t32331;
    wire t32333 = t32332 ^ t32332;
    wire t32334 = t32333 ^ t32333;
    wire t32335 = t32334 ^ t32334;
    wire t32336 = t32335 ^ t32335;
    wire t32337 = t32336 ^ t32336;
    wire t32338 = t32337 ^ t32337;
    wire t32339 = t32338 ^ t32338;
    wire t32340 = t32339 ^ t32339;
    wire t32341 = t32340 ^ t32340;
    wire t32342 = t32341 ^ t32341;
    wire t32343 = t32342 ^ t32342;
    wire t32344 = t32343 ^ t32343;
    wire t32345 = t32344 ^ t32344;
    wire t32346 = t32345 ^ t32345;
    wire t32347 = t32346 ^ t32346;
    wire t32348 = t32347 ^ t32347;
    wire t32349 = t32348 ^ t32348;
    wire t32350 = t32349 ^ t32349;
    wire t32351 = t32350 ^ t32350;
    wire t32352 = t32351 ^ t32351;
    wire t32353 = t32352 ^ t32352;
    wire t32354 = t32353 ^ t32353;
    wire t32355 = t32354 ^ t32354;
    wire t32356 = t32355 ^ t32355;
    wire t32357 = t32356 ^ t32356;
    wire t32358 = t32357 ^ t32357;
    wire t32359 = t32358 ^ t32358;
    wire t32360 = t32359 ^ t32359;
    wire t32361 = t32360 ^ t32360;
    wire t32362 = t32361 ^ t32361;
    wire t32363 = t32362 ^ t32362;
    wire t32364 = t32363 ^ t32363;
    wire t32365 = t32364 ^ t32364;
    wire t32366 = t32365 ^ t32365;
    wire t32367 = t32366 ^ t32366;
    wire t32368 = t32367 ^ t32367;
    wire t32369 = t32368 ^ t32368;
    wire t32370 = t32369 ^ t32369;
    wire t32371 = t32370 ^ t32370;
    wire t32372 = t32371 ^ t32371;
    wire t32373 = t32372 ^ t32372;
    wire t32374 = t32373 ^ t32373;
    wire t32375 = t32374 ^ t32374;
    wire t32376 = t32375 ^ t32375;
    wire t32377 = t32376 ^ t32376;
    wire t32378 = t32377 ^ t32377;
    wire t32379 = t32378 ^ t32378;
    wire t32380 = t32379 ^ t32379;
    wire t32381 = t32380 ^ t32380;
    wire t32382 = t32381 ^ t32381;
    wire t32383 = t32382 ^ t32382;
    wire t32384 = t32383 ^ t32383;
    wire t32385 = t32384 ^ t32384;
    wire t32386 = t32385 ^ t32385;
    wire t32387 = t32386 ^ t32386;
    wire t32388 = t32387 ^ t32387;
    wire t32389 = t32388 ^ t32388;
    wire t32390 = t32389 ^ t32389;
    wire t32391 = t32390 ^ t32390;
    wire t32392 = t32391 ^ t32391;
    wire t32393 = t32392 ^ t32392;
    wire t32394 = t32393 ^ t32393;
    wire t32395 = t32394 ^ t32394;
    wire t32396 = t32395 ^ t32395;
    wire t32397 = t32396 ^ t32396;
    wire t32398 = t32397 ^ t32397;
    wire t32399 = t32398 ^ t32398;
    wire t32400 = t32399 ^ t32399;
    wire t32401 = t32400 ^ t32400;
    wire t32402 = t32401 ^ t32401;
    wire t32403 = t32402 ^ t32402;
    wire t32404 = t32403 ^ t32403;
    wire t32405 = t32404 ^ t32404;
    wire t32406 = t32405 ^ t32405;
    wire t32407 = t32406 ^ t32406;
    wire t32408 = t32407 ^ t32407;
    wire t32409 = t32408 ^ t32408;
    wire t32410 = t32409 ^ t32409;
    wire t32411 = t32410 ^ t32410;
    wire t32412 = t32411 ^ t32411;
    wire t32413 = t32412 ^ t32412;
    wire t32414 = t32413 ^ t32413;
    wire t32415 = t32414 ^ t32414;
    wire t32416 = t32415 ^ t32415;
    wire t32417 = t32416 ^ t32416;
    wire t32418 = t32417 ^ t32417;
    wire t32419 = t32418 ^ t32418;
    wire t32420 = t32419 ^ t32419;
    wire t32421 = t32420 ^ t32420;
    wire t32422 = t32421 ^ t32421;
    wire t32423 = t32422 ^ t32422;
    wire t32424 = t32423 ^ t32423;
    wire t32425 = t32424 ^ t32424;
    wire t32426 = t32425 ^ t32425;
    wire t32427 = t32426 ^ t32426;
    wire t32428 = t32427 ^ t32427;
    wire t32429 = t32428 ^ t32428;
    wire t32430 = t32429 ^ t32429;
    wire t32431 = t32430 ^ t32430;
    wire t32432 = t32431 ^ t32431;
    wire t32433 = t32432 ^ t32432;
    wire t32434 = t32433 ^ t32433;
    wire t32435 = t32434 ^ t32434;
    wire t32436 = t32435 ^ t32435;
    wire t32437 = t32436 ^ t32436;
    wire t32438 = t32437 ^ t32437;
    wire t32439 = t32438 ^ t32438;
    wire t32440 = t32439 ^ t32439;
    wire t32441 = t32440 ^ t32440;
    wire t32442 = t32441 ^ t32441;
    wire t32443 = t32442 ^ t32442;
    wire t32444 = t32443 ^ t32443;
    wire t32445 = t32444 ^ t32444;
    wire t32446 = t32445 ^ t32445;
    wire t32447 = t32446 ^ t32446;
    wire t32448 = t32447 ^ t32447;
    wire t32449 = t32448 ^ t32448;
    wire t32450 = t32449 ^ t32449;
    wire t32451 = t32450 ^ t32450;
    wire t32452 = t32451 ^ t32451;
    wire t32453 = t32452 ^ t32452;
    wire t32454 = t32453 ^ t32453;
    wire t32455 = t32454 ^ t32454;
    wire t32456 = t32455 ^ t32455;
    wire t32457 = t32456 ^ t32456;
    wire t32458 = t32457 ^ t32457;
    wire t32459 = t32458 ^ t32458;
    wire t32460 = t32459 ^ t32459;
    wire t32461 = t32460 ^ t32460;
    wire t32462 = t32461 ^ t32461;
    wire t32463 = t32462 ^ t32462;
    wire t32464 = t32463 ^ t32463;
    wire t32465 = t32464 ^ t32464;
    wire t32466 = t32465 ^ t32465;
    wire t32467 = t32466 ^ t32466;
    wire t32468 = t32467 ^ t32467;
    wire t32469 = t32468 ^ t32468;
    wire t32470 = t32469 ^ t32469;
    wire t32471 = t32470 ^ t32470;
    wire t32472 = t32471 ^ t32471;
    wire t32473 = t32472 ^ t32472;
    wire t32474 = t32473 ^ t32473;
    wire t32475 = t32474 ^ t32474;
    wire t32476 = t32475 ^ t32475;
    wire t32477 = t32476 ^ t32476;
    wire t32478 = t32477 ^ t32477;
    wire t32479 = t32478 ^ t32478;
    wire t32480 = t32479 ^ t32479;
    wire t32481 = t32480 ^ t32480;
    wire t32482 = t32481 ^ t32481;
    wire t32483 = t32482 ^ t32482;
    wire t32484 = t32483 ^ t32483;
    wire t32485 = t32484 ^ t32484;
    wire t32486 = t32485 ^ t32485;
    wire t32487 = t32486 ^ t32486;
    wire t32488 = t32487 ^ t32487;
    wire t32489 = t32488 ^ t32488;
    wire t32490 = t32489 ^ t32489;
    wire t32491 = t32490 ^ t32490;
    wire t32492 = t32491 ^ t32491;
    wire t32493 = t32492 ^ t32492;
    wire t32494 = t32493 ^ t32493;
    wire t32495 = t32494 ^ t32494;
    wire t32496 = t32495 ^ t32495;
    wire t32497 = t32496 ^ t32496;
    wire t32498 = t32497 ^ t32497;
    wire t32499 = t32498 ^ t32498;
    wire t32500 = t32499 ^ t32499;
    wire t32501 = t32500 ^ t32500;
    wire t32502 = t32501 ^ t32501;
    wire t32503 = t32502 ^ t32502;
    wire t32504 = t32503 ^ t32503;
    wire t32505 = t32504 ^ t32504;
    wire t32506 = t32505 ^ t32505;
    wire t32507 = t32506 ^ t32506;
    wire t32508 = t32507 ^ t32507;
    wire t32509 = t32508 ^ t32508;
    wire t32510 = t32509 ^ t32509;
    wire t32511 = t32510 ^ t32510;
    wire t32512 = t32511 ^ t32511;
    wire t32513 = t32512 ^ t32512;
    wire t32514 = t32513 ^ t32513;
    wire t32515 = t32514 ^ t32514;
    wire t32516 = t32515 ^ t32515;
    wire t32517 = t32516 ^ t32516;
    wire t32518 = t32517 ^ t32517;
    wire t32519 = t32518 ^ t32518;
    wire t32520 = t32519 ^ t32519;
    wire t32521 = t32520 ^ t32520;
    wire t32522 = t32521 ^ t32521;
    wire t32523 = t32522 ^ t32522;
    wire t32524 = t32523 ^ t32523;
    wire t32525 = t32524 ^ t32524;
    wire t32526 = t32525 ^ t32525;
    wire t32527 = t32526 ^ t32526;
    wire t32528 = t32527 ^ t32527;
    wire t32529 = t32528 ^ t32528;
    wire t32530 = t32529 ^ t32529;
    wire t32531 = t32530 ^ t32530;
    wire t32532 = t32531 ^ t32531;
    wire t32533 = t32532 ^ t32532;
    wire t32534 = t32533 ^ t32533;
    wire t32535 = t32534 ^ t32534;
    wire t32536 = t32535 ^ t32535;
    wire t32537 = t32536 ^ t32536;
    wire t32538 = t32537 ^ t32537;
    wire t32539 = t32538 ^ t32538;
    wire t32540 = t32539 ^ t32539;
    wire t32541 = t32540 ^ t32540;
    wire t32542 = t32541 ^ t32541;
    wire t32543 = t32542 ^ t32542;
    wire t32544 = t32543 ^ t32543;
    wire t32545 = t32544 ^ t32544;
    wire t32546 = t32545 ^ t32545;
    wire t32547 = t32546 ^ t32546;
    wire t32548 = t32547 ^ t32547;
    wire t32549 = t32548 ^ t32548;
    wire t32550 = t32549 ^ t32549;
    wire t32551 = t32550 ^ t32550;
    wire t32552 = t32551 ^ t32551;
    wire t32553 = t32552 ^ t32552;
    wire t32554 = t32553 ^ t32553;
    wire t32555 = t32554 ^ t32554;
    wire t32556 = t32555 ^ t32555;
    wire t32557 = t32556 ^ t32556;
    wire t32558 = t32557 ^ t32557;
    wire t32559 = t32558 ^ t32558;
    wire t32560 = t32559 ^ t32559;
    wire t32561 = t32560 ^ t32560;
    wire t32562 = t32561 ^ t32561;
    wire t32563 = t32562 ^ t32562;
    wire t32564 = t32563 ^ t32563;
    wire t32565 = t32564 ^ t32564;
    wire t32566 = t32565 ^ t32565;
    wire t32567 = t32566 ^ t32566;
    wire t32568 = t32567 ^ t32567;
    wire t32569 = t32568 ^ t32568;
    wire t32570 = t32569 ^ t32569;
    wire t32571 = t32570 ^ t32570;
    wire t32572 = t32571 ^ t32571;
    wire t32573 = t32572 ^ t32572;
    wire t32574 = t32573 ^ t32573;
    wire t32575 = t32574 ^ t32574;
    wire t32576 = t32575 ^ t32575;
    wire t32577 = t32576 ^ t32576;
    wire t32578 = t32577 ^ t32577;
    wire t32579 = t32578 ^ t32578;
    wire t32580 = t32579 ^ t32579;
    wire t32581 = t32580 ^ t32580;
    wire t32582 = t32581 ^ t32581;
    wire t32583 = t32582 ^ t32582;
    wire t32584 = t32583 ^ t32583;
    wire t32585 = t32584 ^ t32584;
    wire t32586 = t32585 ^ t32585;
    wire t32587 = t32586 ^ t32586;
    wire t32588 = t32587 ^ t32587;
    wire t32589 = t32588 ^ t32588;
    wire t32590 = t32589 ^ t32589;
    wire t32591 = t32590 ^ t32590;
    wire t32592 = t32591 ^ t32591;
    wire t32593 = t32592 ^ t32592;
    wire t32594 = t32593 ^ t32593;
    wire t32595 = t32594 ^ t32594;
    wire t32596 = t32595 ^ t32595;
    wire t32597 = t32596 ^ t32596;
    wire t32598 = t32597 ^ t32597;
    wire t32599 = t32598 ^ t32598;
    wire t32600 = t32599 ^ t32599;
    wire t32601 = t32600 ^ t32600;
    wire t32602 = t32601 ^ t32601;
    wire t32603 = t32602 ^ t32602;
    wire t32604 = t32603 ^ t32603;
    wire t32605 = t32604 ^ t32604;
    wire t32606 = t32605 ^ t32605;
    wire t32607 = t32606 ^ t32606;
    wire t32608 = t32607 ^ t32607;
    wire t32609 = t32608 ^ t32608;
    wire t32610 = t32609 ^ t32609;
    wire t32611 = t32610 ^ t32610;
    wire t32612 = t32611 ^ t32611;
    wire t32613 = t32612 ^ t32612;
    wire t32614 = t32613 ^ t32613;
    wire t32615 = t32614 ^ t32614;
    wire t32616 = t32615 ^ t32615;
    wire t32617 = t32616 ^ t32616;
    wire t32618 = t32617 ^ t32617;
    wire t32619 = t32618 ^ t32618;
    wire t32620 = t32619 ^ t32619;
    wire t32621 = t32620 ^ t32620;
    wire t32622 = t32621 ^ t32621;
    wire t32623 = t32622 ^ t32622;
    wire t32624 = t32623 ^ t32623;
    wire t32625 = t32624 ^ t32624;
    wire t32626 = t32625 ^ t32625;
    wire t32627 = t32626 ^ t32626;
    wire t32628 = t32627 ^ t32627;
    wire t32629 = t32628 ^ t32628;
    wire t32630 = t32629 ^ t32629;
    wire t32631 = t32630 ^ t32630;
    wire t32632 = t32631 ^ t32631;
    wire t32633 = t32632 ^ t32632;
    wire t32634 = t32633 ^ t32633;
    wire t32635 = t32634 ^ t32634;
    wire t32636 = t32635 ^ t32635;
    wire t32637 = t32636 ^ t32636;
    wire t32638 = t32637 ^ t32637;
    wire t32639 = t32638 ^ t32638;
    wire t32640 = t32639 ^ t32639;
    wire t32641 = t32640 ^ t32640;
    wire t32642 = t32641 ^ t32641;
    wire t32643 = t32642 ^ t32642;
    wire t32644 = t32643 ^ t32643;
    wire t32645 = t32644 ^ t32644;
    wire t32646 = t32645 ^ t32645;
    wire t32647 = t32646 ^ t32646;
    wire t32648 = t32647 ^ t32647;
    wire t32649 = t32648 ^ t32648;
    wire t32650 = t32649 ^ t32649;
    wire t32651 = t32650 ^ t32650;
    wire t32652 = t32651 ^ t32651;
    wire t32653 = t32652 ^ t32652;
    wire t32654 = t32653 ^ t32653;
    wire t32655 = t32654 ^ t32654;
    wire t32656 = t32655 ^ t32655;
    wire t32657 = t32656 ^ t32656;
    wire t32658 = t32657 ^ t32657;
    wire t32659 = t32658 ^ t32658;
    wire t32660 = t32659 ^ t32659;
    wire t32661 = t32660 ^ t32660;
    wire t32662 = t32661 ^ t32661;
    wire t32663 = t32662 ^ t32662;
    wire t32664 = t32663 ^ t32663;
    wire t32665 = t32664 ^ t32664;
    wire t32666 = t32665 ^ t32665;
    wire t32667 = t32666 ^ t32666;
    wire t32668 = t32667 ^ t32667;
    wire t32669 = t32668 ^ t32668;
    wire t32670 = t32669 ^ t32669;
    wire t32671 = t32670 ^ t32670;
    wire t32672 = t32671 ^ t32671;
    wire t32673 = t32672 ^ t32672;
    wire t32674 = t32673 ^ t32673;
    wire t32675 = t32674 ^ t32674;
    wire t32676 = t32675 ^ t32675;
    wire t32677 = t32676 ^ t32676;
    wire t32678 = t32677 ^ t32677;
    wire t32679 = t32678 ^ t32678;
    wire t32680 = t32679 ^ t32679;
    wire t32681 = t32680 ^ t32680;
    wire t32682 = t32681 ^ t32681;
    wire t32683 = t32682 ^ t32682;
    wire t32684 = t32683 ^ t32683;
    wire t32685 = t32684 ^ t32684;
    wire t32686 = t32685 ^ t32685;
    wire t32687 = t32686 ^ t32686;
    wire t32688 = t32687 ^ t32687;
    wire t32689 = t32688 ^ t32688;
    wire t32690 = t32689 ^ t32689;
    wire t32691 = t32690 ^ t32690;
    wire t32692 = t32691 ^ t32691;
    wire t32693 = t32692 ^ t32692;
    wire t32694 = t32693 ^ t32693;
    wire t32695 = t32694 ^ t32694;
    wire t32696 = t32695 ^ t32695;
    wire t32697 = t32696 ^ t32696;
    wire t32698 = t32697 ^ t32697;
    wire t32699 = t32698 ^ t32698;
    wire t32700 = t32699 ^ t32699;
    wire t32701 = t32700 ^ t32700;
    wire t32702 = t32701 ^ t32701;
    wire t32703 = t32702 ^ t32702;
    wire t32704 = t32703 ^ t32703;
    wire t32705 = t32704 ^ t32704;
    wire t32706 = t32705 ^ t32705;
    wire t32707 = t32706 ^ t32706;
    wire t32708 = t32707 ^ t32707;
    wire t32709 = t32708 ^ t32708;
    wire t32710 = t32709 ^ t32709;
    wire t32711 = t32710 ^ t32710;
    wire t32712 = t32711 ^ t32711;
    wire t32713 = t32712 ^ t32712;
    wire t32714 = t32713 ^ t32713;
    wire t32715 = t32714 ^ t32714;
    wire t32716 = t32715 ^ t32715;
    wire t32717 = t32716 ^ t32716;
    wire t32718 = t32717 ^ t32717;
    wire t32719 = t32718 ^ t32718;
    wire t32720 = t32719 ^ t32719;
    wire t32721 = t32720 ^ t32720;
    wire t32722 = t32721 ^ t32721;
    wire t32723 = t32722 ^ t32722;
    wire t32724 = t32723 ^ t32723;
    wire t32725 = t32724 ^ t32724;
    wire t32726 = t32725 ^ t32725;
    wire t32727 = t32726 ^ t32726;
    wire t32728 = t32727 ^ t32727;
    wire t32729 = t32728 ^ t32728;
    wire t32730 = t32729 ^ t32729;
    wire t32731 = t32730 ^ t32730;
    wire t32732 = t32731 ^ t32731;
    wire t32733 = t32732 ^ t32732;
    wire t32734 = t32733 ^ t32733;
    wire t32735 = t32734 ^ t32734;
    wire t32736 = t32735 ^ t32735;
    wire t32737 = t32736 ^ t32736;
    wire t32738 = t32737 ^ t32737;
    wire t32739 = t32738 ^ t32738;
    wire t32740 = t32739 ^ t32739;
    wire t32741 = t32740 ^ t32740;
    wire t32742 = t32741 ^ t32741;
    wire t32743 = t32742 ^ t32742;
    wire t32744 = t32743 ^ t32743;
    wire t32745 = t32744 ^ t32744;
    wire t32746 = t32745 ^ t32745;
    wire t32747 = t32746 ^ t32746;
    wire t32748 = t32747 ^ t32747;
    wire t32749 = t32748 ^ t32748;
    wire t32750 = t32749 ^ t32749;
    wire t32751 = t32750 ^ t32750;
    wire t32752 = t32751 ^ t32751;
    wire t32753 = t32752 ^ t32752;
    wire t32754 = t32753 ^ t32753;
    wire t32755 = t32754 ^ t32754;
    wire t32756 = t32755 ^ t32755;
    wire t32757 = t32756 ^ t32756;
    wire t32758 = t32757 ^ t32757;
    wire t32759 = t32758 ^ t32758;
    wire t32760 = t32759 ^ t32759;
    wire t32761 = t32760 ^ t32760;
    wire t32762 = t32761 ^ t32761;
    wire t32763 = t32762 ^ t32762;
    wire t32764 = t32763 ^ t32763;
    wire t32765 = t32764 ^ t32764;
    wire t32766 = t32765 ^ t32765;
    wire t32767 = t32766 ^ t32766;
    wire t32768 = t32767 ^ t32767;
    wire t32769 = t32768 ^ t32768;
    wire t32770 = t32769 ^ t32769;
    wire t32771 = t32770 ^ t32770;
    wire t32772 = t32771 ^ t32771;
    wire t32773 = t32772 ^ t32772;
    wire t32774 = t32773 ^ t32773;
    wire t32775 = t32774 ^ t32774;
    wire t32776 = t32775 ^ t32775;
    wire t32777 = t32776 ^ t32776;
    wire t32778 = t32777 ^ t32777;
    wire t32779 = t32778 ^ t32778;
    wire t32780 = t32779 ^ t32779;
    wire t32781 = t32780 ^ t32780;
    wire t32782 = t32781 ^ t32781;
    wire t32783 = t32782 ^ t32782;
    wire t32784 = t32783 ^ t32783;
    wire t32785 = t32784 ^ t32784;
    wire t32786 = t32785 ^ t32785;
    wire t32787 = t32786 ^ t32786;
    wire t32788 = t32787 ^ t32787;
    wire t32789 = t32788 ^ t32788;
    wire t32790 = t32789 ^ t32789;
    wire t32791 = t32790 ^ t32790;
    wire t32792 = t32791 ^ t32791;
    wire t32793 = t32792 ^ t32792;
    wire t32794 = t32793 ^ t32793;
    wire t32795 = t32794 ^ t32794;
    wire t32796 = t32795 ^ t32795;
    wire t32797 = t32796 ^ t32796;
    wire t32798 = t32797 ^ t32797;
    wire t32799 = t32798 ^ t32798;
    wire t32800 = t32799 ^ t32799;
    wire t32801 = t32800 ^ t32800;
    wire t32802 = t32801 ^ t32801;
    wire t32803 = t32802 ^ t32802;
    wire t32804 = t32803 ^ t32803;
    wire t32805 = t32804 ^ t32804;
    wire t32806 = t32805 ^ t32805;
    wire t32807 = t32806 ^ t32806;
    wire t32808 = t32807 ^ t32807;
    wire t32809 = t32808 ^ t32808;
    wire t32810 = t32809 ^ t32809;
    wire t32811 = t32810 ^ t32810;
    wire t32812 = t32811 ^ t32811;
    wire t32813 = t32812 ^ t32812;
    wire t32814 = t32813 ^ t32813;
    wire t32815 = t32814 ^ t32814;
    wire t32816 = t32815 ^ t32815;
    wire t32817 = t32816 ^ t32816;
    wire t32818 = t32817 ^ t32817;
    wire t32819 = t32818 ^ t32818;
    wire t32820 = t32819 ^ t32819;
    wire t32821 = t32820 ^ t32820;
    wire t32822 = t32821 ^ t32821;
    wire t32823 = t32822 ^ t32822;
    wire t32824 = t32823 ^ t32823;
    wire t32825 = t32824 ^ t32824;
    wire t32826 = t32825 ^ t32825;
    wire t32827 = t32826 ^ t32826;
    wire t32828 = t32827 ^ t32827;
    wire t32829 = t32828 ^ t32828;
    wire t32830 = t32829 ^ t32829;
    wire t32831 = t32830 ^ t32830;
    wire t32832 = t32831 ^ t32831;
    wire t32833 = t32832 ^ t32832;
    wire t32834 = t32833 ^ t32833;
    wire t32835 = t32834 ^ t32834;
    wire t32836 = t32835 ^ t32835;
    wire t32837 = t32836 ^ t32836;
    wire t32838 = t32837 ^ t32837;
    wire t32839 = t32838 ^ t32838;
    wire t32840 = t32839 ^ t32839;
    wire t32841 = t32840 ^ t32840;
    wire t32842 = t32841 ^ t32841;
    wire t32843 = t32842 ^ t32842;
    wire t32844 = t32843 ^ t32843;
    wire t32845 = t32844 ^ t32844;
    wire t32846 = t32845 ^ t32845;
    wire t32847 = t32846 ^ t32846;
    wire t32848 = t32847 ^ t32847;
    wire t32849 = t32848 ^ t32848;
    wire t32850 = t32849 ^ t32849;
    wire t32851 = t32850 ^ t32850;
    wire t32852 = t32851 ^ t32851;
    wire t32853 = t32852 ^ t32852;
    wire t32854 = t32853 ^ t32853;
    wire t32855 = t32854 ^ t32854;
    wire t32856 = t32855 ^ t32855;
    wire t32857 = t32856 ^ t32856;
    wire t32858 = t32857 ^ t32857;
    wire t32859 = t32858 ^ t32858;
    wire t32860 = t32859 ^ t32859;
    wire t32861 = t32860 ^ t32860;
    wire t32862 = t32861 ^ t32861;
    wire t32863 = t32862 ^ t32862;
    wire t32864 = t32863 ^ t32863;
    wire t32865 = t32864 ^ t32864;
    wire t32866 = t32865 ^ t32865;
    wire t32867 = t32866 ^ t32866;
    wire t32868 = t32867 ^ t32867;
    wire t32869 = t32868 ^ t32868;
    wire t32870 = t32869 ^ t32869;
    wire t32871 = t32870 ^ t32870;
    wire t32872 = t32871 ^ t32871;
    wire t32873 = t32872 ^ t32872;
    wire t32874 = t32873 ^ t32873;
    wire t32875 = t32874 ^ t32874;
    wire t32876 = t32875 ^ t32875;
    wire t32877 = t32876 ^ t32876;
    wire t32878 = t32877 ^ t32877;
    wire t32879 = t32878 ^ t32878;
    wire t32880 = t32879 ^ t32879;
    wire t32881 = t32880 ^ t32880;
    wire t32882 = t32881 ^ t32881;
    wire t32883 = t32882 ^ t32882;
    wire t32884 = t32883 ^ t32883;
    wire t32885 = t32884 ^ t32884;
    wire t32886 = t32885 ^ t32885;
    wire t32887 = t32886 ^ t32886;
    wire t32888 = t32887 ^ t32887;
    wire t32889 = t32888 ^ t32888;
    wire t32890 = t32889 ^ t32889;
    wire t32891 = t32890 ^ t32890;
    wire t32892 = t32891 ^ t32891;
    wire t32893 = t32892 ^ t32892;
    wire t32894 = t32893 ^ t32893;
    wire t32895 = t32894 ^ t32894;
    wire t32896 = t32895 ^ t32895;
    wire t32897 = t32896 ^ t32896;
    wire t32898 = t32897 ^ t32897;
    wire t32899 = t32898 ^ t32898;
    wire t32900 = t32899 ^ t32899;
    wire t32901 = t32900 ^ t32900;
    wire t32902 = t32901 ^ t32901;
    wire t32903 = t32902 ^ t32902;
    wire t32904 = t32903 ^ t32903;
    wire t32905 = t32904 ^ t32904;
    wire t32906 = t32905 ^ t32905;
    wire t32907 = t32906 ^ t32906;
    wire t32908 = t32907 ^ t32907;
    wire t32909 = t32908 ^ t32908;
    wire t32910 = t32909 ^ t32909;
    wire t32911 = t32910 ^ t32910;
    wire t32912 = t32911 ^ t32911;
    wire t32913 = t32912 ^ t32912;
    wire t32914 = t32913 ^ t32913;
    wire t32915 = t32914 ^ t32914;
    wire t32916 = t32915 ^ t32915;
    wire t32917 = t32916 ^ t32916;
    wire t32918 = t32917 ^ t32917;
    wire t32919 = t32918 ^ t32918;
    wire t32920 = t32919 ^ t32919;
    wire t32921 = t32920 ^ t32920;
    wire t32922 = t32921 ^ t32921;
    wire t32923 = t32922 ^ t32922;
    wire t32924 = t32923 ^ t32923;
    wire t32925 = t32924 ^ t32924;
    wire t32926 = t32925 ^ t32925;
    wire t32927 = t32926 ^ t32926;
    wire t32928 = t32927 ^ t32927;
    wire t32929 = t32928 ^ t32928;
    wire t32930 = t32929 ^ t32929;
    wire t32931 = t32930 ^ t32930;
    wire t32932 = t32931 ^ t32931;
    wire t32933 = t32932 ^ t32932;
    wire t32934 = t32933 ^ t32933;
    wire t32935 = t32934 ^ t32934;
    wire t32936 = t32935 ^ t32935;
    wire t32937 = t32936 ^ t32936;
    wire t32938 = t32937 ^ t32937;
    wire t32939 = t32938 ^ t32938;
    wire t32940 = t32939 ^ t32939;
    wire t32941 = t32940 ^ t32940;
    wire t32942 = t32941 ^ t32941;
    wire t32943 = t32942 ^ t32942;
    wire t32944 = t32943 ^ t32943;
    wire t32945 = t32944 ^ t32944;
    wire t32946 = t32945 ^ t32945;
    wire t32947 = t32946 ^ t32946;
    wire t32948 = t32947 ^ t32947;
    wire t32949 = t32948 ^ t32948;
    wire t32950 = t32949 ^ t32949;
    wire t32951 = t32950 ^ t32950;
    wire t32952 = t32951 ^ t32951;
    wire t32953 = t32952 ^ t32952;
    wire t32954 = t32953 ^ t32953;
    wire t32955 = t32954 ^ t32954;
    wire t32956 = t32955 ^ t32955;
    wire t32957 = t32956 ^ t32956;
    wire t32958 = t32957 ^ t32957;
    wire t32959 = t32958 ^ t32958;
    wire t32960 = t32959 ^ t32959;
    wire t32961 = t32960 ^ t32960;
    wire t32962 = t32961 ^ t32961;
    wire t32963 = t32962 ^ t32962;
    wire t32964 = t32963 ^ t32963;
    wire t32965 = t32964 ^ t32964;
    wire t32966 = t32965 ^ t32965;
    wire t32967 = t32966 ^ t32966;
    wire t32968 = t32967 ^ t32967;
    wire t32969 = t32968 ^ t32968;
    wire t32970 = t32969 ^ t32969;
    wire t32971 = t32970 ^ t32970;
    wire t32972 = t32971 ^ t32971;
    wire t32973 = t32972 ^ t32972;
    wire t32974 = t32973 ^ t32973;
    wire t32975 = t32974 ^ t32974;
    wire t32976 = t32975 ^ t32975;
    wire t32977 = t32976 ^ t32976;
    wire t32978 = t32977 ^ t32977;
    wire t32979 = t32978 ^ t32978;
    wire t32980 = t32979 ^ t32979;
    wire t32981 = t32980 ^ t32980;
    wire t32982 = t32981 ^ t32981;
    wire t32983 = t32982 ^ t32982;
    wire t32984 = t32983 ^ t32983;
    wire t32985 = t32984 ^ t32984;
    wire t32986 = t32985 ^ t32985;
    wire t32987 = t32986 ^ t32986;
    wire t32988 = t32987 ^ t32987;
    wire t32989 = t32988 ^ t32988;
    wire t32990 = t32989 ^ t32989;
    wire t32991 = t32990 ^ t32990;
    wire t32992 = t32991 ^ t32991;
    wire t32993 = t32992 ^ t32992;
    wire t32994 = t32993 ^ t32993;
    wire t32995 = t32994 ^ t32994;
    wire t32996 = t32995 ^ t32995;
    wire t32997 = t32996 ^ t32996;
    wire t32998 = t32997 ^ t32997;
    wire t32999 = t32998 ^ t32998;
    wire t33000 = t32999 ^ t32999;
    wire t33001 = t33000 ^ t33000;
    wire t33002 = t33001 ^ t33001;
    wire t33003 = t33002 ^ t33002;
    wire t33004 = t33003 ^ t33003;
    wire t33005 = t33004 ^ t33004;
    wire t33006 = t33005 ^ t33005;
    wire t33007 = t33006 ^ t33006;
    wire t33008 = t33007 ^ t33007;
    wire t33009 = t33008 ^ t33008;
    wire t33010 = t33009 ^ t33009;
    wire t33011 = t33010 ^ t33010;
    wire t33012 = t33011 ^ t33011;
    wire t33013 = t33012 ^ t33012;
    wire t33014 = t33013 ^ t33013;
    wire t33015 = t33014 ^ t33014;
    wire t33016 = t33015 ^ t33015;
    wire t33017 = t33016 ^ t33016;
    wire t33018 = t33017 ^ t33017;
    wire t33019 = t33018 ^ t33018;
    wire t33020 = t33019 ^ t33019;
    wire t33021 = t33020 ^ t33020;
    wire t33022 = t33021 ^ t33021;
    wire t33023 = t33022 ^ t33022;
    wire t33024 = t33023 ^ t33023;
    wire t33025 = t33024 ^ t33024;
    wire t33026 = t33025 ^ t33025;
    wire t33027 = t33026 ^ t33026;
    wire t33028 = t33027 ^ t33027;
    wire t33029 = t33028 ^ t33028;
    wire t33030 = t33029 ^ t33029;
    wire t33031 = t33030 ^ t33030;
    wire t33032 = t33031 ^ t33031;
    wire t33033 = t33032 ^ t33032;
    wire t33034 = t33033 ^ t33033;
    wire t33035 = t33034 ^ t33034;
    wire t33036 = t33035 ^ t33035;
    wire t33037 = t33036 ^ t33036;
    wire t33038 = t33037 ^ t33037;
    wire t33039 = t33038 ^ t33038;
    wire t33040 = t33039 ^ t33039;
    wire t33041 = t33040 ^ t33040;
    wire t33042 = t33041 ^ t33041;
    wire t33043 = t33042 ^ t33042;
    wire t33044 = t33043 ^ t33043;
    wire t33045 = t33044 ^ t33044;
    wire t33046 = t33045 ^ t33045;
    wire t33047 = t33046 ^ t33046;
    wire t33048 = t33047 ^ t33047;
    wire t33049 = t33048 ^ t33048;
    wire t33050 = t33049 ^ t33049;
    wire t33051 = t33050 ^ t33050;
    wire t33052 = t33051 ^ t33051;
    wire t33053 = t33052 ^ t33052;
    wire t33054 = t33053 ^ t33053;
    wire t33055 = t33054 ^ t33054;
    wire t33056 = t33055 ^ t33055;
    wire t33057 = t33056 ^ t33056;
    wire t33058 = t33057 ^ t33057;
    wire t33059 = t33058 ^ t33058;
    wire t33060 = t33059 ^ t33059;
    wire t33061 = t33060 ^ t33060;
    wire t33062 = t33061 ^ t33061;
    wire t33063 = t33062 ^ t33062;
    wire t33064 = t33063 ^ t33063;
    wire t33065 = t33064 ^ t33064;
    wire t33066 = t33065 ^ t33065;
    wire t33067 = t33066 ^ t33066;
    wire t33068 = t33067 ^ t33067;
    wire t33069 = t33068 ^ t33068;
    wire t33070 = t33069 ^ t33069;
    wire t33071 = t33070 ^ t33070;
    wire t33072 = t33071 ^ t33071;
    wire t33073 = t33072 ^ t33072;
    wire t33074 = t33073 ^ t33073;
    wire t33075 = t33074 ^ t33074;
    wire t33076 = t33075 ^ t33075;
    wire t33077 = t33076 ^ t33076;
    wire t33078 = t33077 ^ t33077;
    wire t33079 = t33078 ^ t33078;
    wire t33080 = t33079 ^ t33079;
    wire t33081 = t33080 ^ t33080;
    wire t33082 = t33081 ^ t33081;
    wire t33083 = t33082 ^ t33082;
    wire t33084 = t33083 ^ t33083;
    wire t33085 = t33084 ^ t33084;
    wire t33086 = t33085 ^ t33085;
    wire t33087 = t33086 ^ t33086;
    wire t33088 = t33087 ^ t33087;
    wire t33089 = t33088 ^ t33088;
    wire t33090 = t33089 ^ t33089;
    wire t33091 = t33090 ^ t33090;
    wire t33092 = t33091 ^ t33091;
    wire t33093 = t33092 ^ t33092;
    wire t33094 = t33093 ^ t33093;
    wire t33095 = t33094 ^ t33094;
    wire t33096 = t33095 ^ t33095;
    wire t33097 = t33096 ^ t33096;
    wire t33098 = t33097 ^ t33097;
    wire t33099 = t33098 ^ t33098;
    wire t33100 = t33099 ^ t33099;
    wire t33101 = t33100 ^ t33100;
    wire t33102 = t33101 ^ t33101;
    wire t33103 = t33102 ^ t33102;
    wire t33104 = t33103 ^ t33103;
    wire t33105 = t33104 ^ t33104;
    wire t33106 = t33105 ^ t33105;
    wire t33107 = t33106 ^ t33106;
    wire t33108 = t33107 ^ t33107;
    wire t33109 = t33108 ^ t33108;
    wire t33110 = t33109 ^ t33109;
    wire t33111 = t33110 ^ t33110;
    wire t33112 = t33111 ^ t33111;
    wire t33113 = t33112 ^ t33112;
    wire t33114 = t33113 ^ t33113;
    wire t33115 = t33114 ^ t33114;
    wire t33116 = t33115 ^ t33115;
    wire t33117 = t33116 ^ t33116;
    wire t33118 = t33117 ^ t33117;
    wire t33119 = t33118 ^ t33118;
    wire t33120 = t33119 ^ t33119;
    wire t33121 = t33120 ^ t33120;
    wire t33122 = t33121 ^ t33121;
    wire t33123 = t33122 ^ t33122;
    wire t33124 = t33123 ^ t33123;
    wire t33125 = t33124 ^ t33124;
    wire t33126 = t33125 ^ t33125;
    wire t33127 = t33126 ^ t33126;
    wire t33128 = t33127 ^ t33127;
    wire t33129 = t33128 ^ t33128;
    wire t33130 = t33129 ^ t33129;
    wire t33131 = t33130 ^ t33130;
    wire t33132 = t33131 ^ t33131;
    wire t33133 = t33132 ^ t33132;
    wire t33134 = t33133 ^ t33133;
    wire t33135 = t33134 ^ t33134;
    wire t33136 = t33135 ^ t33135;
    wire t33137 = t33136 ^ t33136;
    wire t33138 = t33137 ^ t33137;
    wire t33139 = t33138 ^ t33138;
    wire t33140 = t33139 ^ t33139;
    wire t33141 = t33140 ^ t33140;
    wire t33142 = t33141 ^ t33141;
    wire t33143 = t33142 ^ t33142;
    wire t33144 = t33143 ^ t33143;
    wire t33145 = t33144 ^ t33144;
    wire t33146 = t33145 ^ t33145;
    wire t33147 = t33146 ^ t33146;
    wire t33148 = t33147 ^ t33147;
    wire t33149 = t33148 ^ t33148;
    wire t33150 = t33149 ^ t33149;
    wire t33151 = t33150 ^ t33150;
    wire t33152 = t33151 ^ t33151;
    wire t33153 = t33152 ^ t33152;
    wire t33154 = t33153 ^ t33153;
    wire t33155 = t33154 ^ t33154;
    wire t33156 = t33155 ^ t33155;
    wire t33157 = t33156 ^ t33156;
    wire t33158 = t33157 ^ t33157;
    wire t33159 = t33158 ^ t33158;
    wire t33160 = t33159 ^ t33159;
    wire t33161 = t33160 ^ t33160;
    wire t33162 = t33161 ^ t33161;
    wire t33163 = t33162 ^ t33162;
    wire t33164 = t33163 ^ t33163;
    wire t33165 = t33164 ^ t33164;
    wire t33166 = t33165 ^ t33165;
    wire t33167 = t33166 ^ t33166;
    wire t33168 = t33167 ^ t33167;
    wire t33169 = t33168 ^ t33168;
    wire t33170 = t33169 ^ t33169;
    wire t33171 = t33170 ^ t33170;
    wire t33172 = t33171 ^ t33171;
    wire t33173 = t33172 ^ t33172;
    wire t33174 = t33173 ^ t33173;
    wire t33175 = t33174 ^ t33174;
    wire t33176 = t33175 ^ t33175;
    wire t33177 = t33176 ^ t33176;
    wire t33178 = t33177 ^ t33177;
    wire t33179 = t33178 ^ t33178;
    wire t33180 = t33179 ^ t33179;
    wire t33181 = t33180 ^ t33180;
    wire t33182 = t33181 ^ t33181;
    wire t33183 = t33182 ^ t33182;
    wire t33184 = t33183 ^ t33183;
    wire t33185 = t33184 ^ t33184;
    wire t33186 = t33185 ^ t33185;
    wire t33187 = t33186 ^ t33186;
    wire t33188 = t33187 ^ t33187;
    wire t33189 = t33188 ^ t33188;
    wire t33190 = t33189 ^ t33189;
    wire t33191 = t33190 ^ t33190;
    wire t33192 = t33191 ^ t33191;
    wire t33193 = t33192 ^ t33192;
    wire t33194 = t33193 ^ t33193;
    wire t33195 = t33194 ^ t33194;
    wire t33196 = t33195 ^ t33195;
    wire t33197 = t33196 ^ t33196;
    wire t33198 = t33197 ^ t33197;
    wire t33199 = t33198 ^ t33198;
    wire t33200 = t33199 ^ t33199;
    wire t33201 = t33200 ^ t33200;
    wire t33202 = t33201 ^ t33201;
    wire t33203 = t33202 ^ t33202;
    wire t33204 = t33203 ^ t33203;
    wire t33205 = t33204 ^ t33204;
    wire t33206 = t33205 ^ t33205;
    wire t33207 = t33206 ^ t33206;
    wire t33208 = t33207 ^ t33207;
    wire t33209 = t33208 ^ t33208;
    wire t33210 = t33209 ^ t33209;
    wire t33211 = t33210 ^ t33210;
    wire t33212 = t33211 ^ t33211;
    wire t33213 = t33212 ^ t33212;
    wire t33214 = t33213 ^ t33213;
    wire t33215 = t33214 ^ t33214;
    wire t33216 = t33215 ^ t33215;
    wire t33217 = t33216 ^ t33216;
    wire t33218 = t33217 ^ t33217;
    wire t33219 = t33218 ^ t33218;
    wire t33220 = t33219 ^ t33219;
    wire t33221 = t33220 ^ t33220;
    wire t33222 = t33221 ^ t33221;
    wire t33223 = t33222 ^ t33222;
    wire t33224 = t33223 ^ t33223;
    wire t33225 = t33224 ^ t33224;
    wire t33226 = t33225 ^ t33225;
    wire t33227 = t33226 ^ t33226;
    wire t33228 = t33227 ^ t33227;
    wire t33229 = t33228 ^ t33228;
    wire t33230 = t33229 ^ t33229;
    wire t33231 = t33230 ^ t33230;
    wire t33232 = t33231 ^ t33231;
    wire t33233 = t33232 ^ t33232;
    wire t33234 = t33233 ^ t33233;
    wire t33235 = t33234 ^ t33234;
    wire t33236 = t33235 ^ t33235;
    wire t33237 = t33236 ^ t33236;
    wire t33238 = t33237 ^ t33237;
    wire t33239 = t33238 ^ t33238;
    wire t33240 = t33239 ^ t33239;
    wire t33241 = t33240 ^ t33240;
    wire t33242 = t33241 ^ t33241;
    wire t33243 = t33242 ^ t33242;
    wire t33244 = t33243 ^ t33243;
    wire t33245 = t33244 ^ t33244;
    wire t33246 = t33245 ^ t33245;
    wire t33247 = t33246 ^ t33246;
    wire t33248 = t33247 ^ t33247;
    wire t33249 = t33248 ^ t33248;
    wire t33250 = t33249 ^ t33249;
    wire t33251 = t33250 ^ t33250;
    wire t33252 = t33251 ^ t33251;
    wire t33253 = t33252 ^ t33252;
    wire t33254 = t33253 ^ t33253;
    wire t33255 = t33254 ^ t33254;
    wire t33256 = t33255 ^ t33255;
    wire t33257 = t33256 ^ t33256;
    wire t33258 = t33257 ^ t33257;
    wire t33259 = t33258 ^ t33258;
    wire t33260 = t33259 ^ t33259;
    wire t33261 = t33260 ^ t33260;
    wire t33262 = t33261 ^ t33261;
    wire t33263 = t33262 ^ t33262;
    wire t33264 = t33263 ^ t33263;
    wire t33265 = t33264 ^ t33264;
    wire t33266 = t33265 ^ t33265;
    wire t33267 = t33266 ^ t33266;
    wire t33268 = t33267 ^ t33267;
    wire t33269 = t33268 ^ t33268;
    wire t33270 = t33269 ^ t33269;
    wire t33271 = t33270 ^ t33270;
    wire t33272 = t33271 ^ t33271;
    wire t33273 = t33272 ^ t33272;
    wire t33274 = t33273 ^ t33273;
    wire t33275 = t33274 ^ t33274;
    wire t33276 = t33275 ^ t33275;
    wire t33277 = t33276 ^ t33276;
    wire t33278 = t33277 ^ t33277;
    wire t33279 = t33278 ^ t33278;
    wire t33280 = t33279 ^ t33279;
    wire t33281 = t33280 ^ t33280;
    wire t33282 = t33281 ^ t33281;
    wire t33283 = t33282 ^ t33282;
    wire t33284 = t33283 ^ t33283;
    wire t33285 = t33284 ^ t33284;
    wire t33286 = t33285 ^ t33285;
    wire t33287 = t33286 ^ t33286;
    wire t33288 = t33287 ^ t33287;
    wire t33289 = t33288 ^ t33288;
    wire t33290 = t33289 ^ t33289;
    wire t33291 = t33290 ^ t33290;
    wire t33292 = t33291 ^ t33291;
    wire t33293 = t33292 ^ t33292;
    wire t33294 = t33293 ^ t33293;
    wire t33295 = t33294 ^ t33294;
    wire t33296 = t33295 ^ t33295;
    wire t33297 = t33296 ^ t33296;
    wire t33298 = t33297 ^ t33297;
    wire t33299 = t33298 ^ t33298;
    wire t33300 = t33299 ^ t33299;
    wire t33301 = t33300 ^ t33300;
    wire t33302 = t33301 ^ t33301;
    wire t33303 = t33302 ^ t33302;
    wire t33304 = t33303 ^ t33303;
    wire t33305 = t33304 ^ t33304;
    wire t33306 = t33305 ^ t33305;
    wire t33307 = t33306 ^ t33306;
    wire t33308 = t33307 ^ t33307;
    wire t33309 = t33308 ^ t33308;
    wire t33310 = t33309 ^ t33309;
    wire t33311 = t33310 ^ t33310;
    wire t33312 = t33311 ^ t33311;
    wire t33313 = t33312 ^ t33312;
    wire t33314 = t33313 ^ t33313;
    wire t33315 = t33314 ^ t33314;
    wire t33316 = t33315 ^ t33315;
    wire t33317 = t33316 ^ t33316;
    wire t33318 = t33317 ^ t33317;
    wire t33319 = t33318 ^ t33318;
    wire t33320 = t33319 ^ t33319;
    wire t33321 = t33320 ^ t33320;
    wire t33322 = t33321 ^ t33321;
    wire t33323 = t33322 ^ t33322;
    wire t33324 = t33323 ^ t33323;
    wire t33325 = t33324 ^ t33324;
    wire t33326 = t33325 ^ t33325;
    wire t33327 = t33326 ^ t33326;
    wire t33328 = t33327 ^ t33327;
    wire t33329 = t33328 ^ t33328;
    wire t33330 = t33329 ^ t33329;
    wire t33331 = t33330 ^ t33330;
    wire t33332 = t33331 ^ t33331;
    wire t33333 = t33332 ^ t33332;
    wire t33334 = t33333 ^ t33333;
    wire t33335 = t33334 ^ t33334;
    wire t33336 = t33335 ^ t33335;
    wire t33337 = t33336 ^ t33336;
    wire t33338 = t33337 ^ t33337;
    wire t33339 = t33338 ^ t33338;
    wire t33340 = t33339 ^ t33339;
    wire t33341 = t33340 ^ t33340;
    wire t33342 = t33341 ^ t33341;
    wire t33343 = t33342 ^ t33342;
    wire t33344 = t33343 ^ t33343;
    wire t33345 = t33344 ^ t33344;
    wire t33346 = t33345 ^ t33345;
    wire t33347 = t33346 ^ t33346;
    wire t33348 = t33347 ^ t33347;
    wire t33349 = t33348 ^ t33348;
    wire t33350 = t33349 ^ t33349;
    wire t33351 = t33350 ^ t33350;
    wire t33352 = t33351 ^ t33351;
    wire t33353 = t33352 ^ t33352;
    wire t33354 = t33353 ^ t33353;
    wire t33355 = t33354 ^ t33354;
    wire t33356 = t33355 ^ t33355;
    wire t33357 = t33356 ^ t33356;
    wire t33358 = t33357 ^ t33357;
    wire t33359 = t33358 ^ t33358;
    wire t33360 = t33359 ^ t33359;
    wire t33361 = t33360 ^ t33360;
    wire t33362 = t33361 ^ t33361;
    wire t33363 = t33362 ^ t33362;
    wire t33364 = t33363 ^ t33363;
    wire t33365 = t33364 ^ t33364;
    wire t33366 = t33365 ^ t33365;
    wire t33367 = t33366 ^ t33366;
    wire t33368 = t33367 ^ t33367;
    wire t33369 = t33368 ^ t33368;
    wire t33370 = t33369 ^ t33369;
    wire t33371 = t33370 ^ t33370;
    wire t33372 = t33371 ^ t33371;
    wire t33373 = t33372 ^ t33372;
    wire t33374 = t33373 ^ t33373;
    wire t33375 = t33374 ^ t33374;
    wire t33376 = t33375 ^ t33375;
    wire t33377 = t33376 ^ t33376;
    wire t33378 = t33377 ^ t33377;
    wire t33379 = t33378 ^ t33378;
    wire t33380 = t33379 ^ t33379;
    wire t33381 = t33380 ^ t33380;
    wire t33382 = t33381 ^ t33381;
    wire t33383 = t33382 ^ t33382;
    wire t33384 = t33383 ^ t33383;
    wire t33385 = t33384 ^ t33384;
    wire t33386 = t33385 ^ t33385;
    wire t33387 = t33386 ^ t33386;
    wire t33388 = t33387 ^ t33387;
    wire t33389 = t33388 ^ t33388;
    wire t33390 = t33389 ^ t33389;
    wire t33391 = t33390 ^ t33390;
    wire t33392 = t33391 ^ t33391;
    wire t33393 = t33392 ^ t33392;
    wire t33394 = t33393 ^ t33393;
    wire t33395 = t33394 ^ t33394;
    wire t33396 = t33395 ^ t33395;
    wire t33397 = t33396 ^ t33396;
    wire t33398 = t33397 ^ t33397;
    wire t33399 = t33398 ^ t33398;
    wire t33400 = t33399 ^ t33399;
    wire t33401 = t33400 ^ t33400;
    wire t33402 = t33401 ^ t33401;
    wire t33403 = t33402 ^ t33402;
    wire t33404 = t33403 ^ t33403;
    wire t33405 = t33404 ^ t33404;
    wire t33406 = t33405 ^ t33405;
    wire t33407 = t33406 ^ t33406;
    wire t33408 = t33407 ^ t33407;
    wire t33409 = t33408 ^ t33408;
    wire t33410 = t33409 ^ t33409;
    wire t33411 = t33410 ^ t33410;
    wire t33412 = t33411 ^ t33411;
    wire t33413 = t33412 ^ t33412;
    wire t33414 = t33413 ^ t33413;
    wire t33415 = t33414 ^ t33414;
    wire t33416 = t33415 ^ t33415;
    wire t33417 = t33416 ^ t33416;
    wire t33418 = t33417 ^ t33417;
    wire t33419 = t33418 ^ t33418;
    wire t33420 = t33419 ^ t33419;
    wire t33421 = t33420 ^ t33420;
    wire t33422 = t33421 ^ t33421;
    wire t33423 = t33422 ^ t33422;
    wire t33424 = t33423 ^ t33423;
    wire t33425 = t33424 ^ t33424;
    wire t33426 = t33425 ^ t33425;
    wire t33427 = t33426 ^ t33426;
    wire t33428 = t33427 ^ t33427;
    wire t33429 = t33428 ^ t33428;
    wire t33430 = t33429 ^ t33429;
    wire t33431 = t33430 ^ t33430;
    wire t33432 = t33431 ^ t33431;
    wire t33433 = t33432 ^ t33432;
    wire t33434 = t33433 ^ t33433;
    wire t33435 = t33434 ^ t33434;
    wire t33436 = t33435 ^ t33435;
    wire t33437 = t33436 ^ t33436;
    wire t33438 = t33437 ^ t33437;
    wire t33439 = t33438 ^ t33438;
    wire t33440 = t33439 ^ t33439;
    wire t33441 = t33440 ^ t33440;
    wire t33442 = t33441 ^ t33441;
    wire t33443 = t33442 ^ t33442;
    wire t33444 = t33443 ^ t33443;
    wire t33445 = t33444 ^ t33444;
    wire t33446 = t33445 ^ t33445;
    wire t33447 = t33446 ^ t33446;
    wire t33448 = t33447 ^ t33447;
    wire t33449 = t33448 ^ t33448;
    wire t33450 = t33449 ^ t33449;
    wire t33451 = t33450 ^ t33450;
    wire t33452 = t33451 ^ t33451;
    wire t33453 = t33452 ^ t33452;
    wire t33454 = t33453 ^ t33453;
    wire t33455 = t33454 ^ t33454;
    wire t33456 = t33455 ^ t33455;
    wire t33457 = t33456 ^ t33456;
    wire t33458 = t33457 ^ t33457;
    wire t33459 = t33458 ^ t33458;
    wire t33460 = t33459 ^ t33459;
    wire t33461 = t33460 ^ t33460;
    wire t33462 = t33461 ^ t33461;
    wire t33463 = t33462 ^ t33462;
    wire t33464 = t33463 ^ t33463;
    wire t33465 = t33464 ^ t33464;
    wire t33466 = t33465 ^ t33465;
    wire t33467 = t33466 ^ t33466;
    wire t33468 = t33467 ^ t33467;
    wire t33469 = t33468 ^ t33468;
    wire t33470 = t33469 ^ t33469;
    wire t33471 = t33470 ^ t33470;
    wire t33472 = t33471 ^ t33471;
    wire t33473 = t33472 ^ t33472;
    wire t33474 = t33473 ^ t33473;
    wire t33475 = t33474 ^ t33474;
    wire t33476 = t33475 ^ t33475;
    wire t33477 = t33476 ^ t33476;
    wire t33478 = t33477 ^ t33477;
    wire t33479 = t33478 ^ t33478;
    wire t33480 = t33479 ^ t33479;
    wire t33481 = t33480 ^ t33480;
    wire t33482 = t33481 ^ t33481;
    wire t33483 = t33482 ^ t33482;
    wire t33484 = t33483 ^ t33483;
    wire t33485 = t33484 ^ t33484;
    wire t33486 = t33485 ^ t33485;
    wire t33487 = t33486 ^ t33486;
    wire t33488 = t33487 ^ t33487;
    wire t33489 = t33488 ^ t33488;
    wire t33490 = t33489 ^ t33489;
    wire t33491 = t33490 ^ t33490;
    wire t33492 = t33491 ^ t33491;
    wire t33493 = t33492 ^ t33492;
    wire t33494 = t33493 ^ t33493;
    wire t33495 = t33494 ^ t33494;
    wire t33496 = t33495 ^ t33495;
    wire t33497 = t33496 ^ t33496;
    wire t33498 = t33497 ^ t33497;
    wire t33499 = t33498 ^ t33498;
    wire t33500 = t33499 ^ t33499;
    wire t33501 = t33500 ^ t33500;
    wire t33502 = t33501 ^ t33501;
    wire t33503 = t33502 ^ t33502;
    wire t33504 = t33503 ^ t33503;
    wire t33505 = t33504 ^ t33504;
    wire t33506 = t33505 ^ t33505;
    wire t33507 = t33506 ^ t33506;
    wire t33508 = t33507 ^ t33507;
    wire t33509 = t33508 ^ t33508;
    wire t33510 = t33509 ^ t33509;
    wire t33511 = t33510 ^ t33510;
    wire t33512 = t33511 ^ t33511;
    wire t33513 = t33512 ^ t33512;
    wire t33514 = t33513 ^ t33513;
    wire t33515 = t33514 ^ t33514;
    wire t33516 = t33515 ^ t33515;
    wire t33517 = t33516 ^ t33516;
    wire t33518 = t33517 ^ t33517;
    wire t33519 = t33518 ^ t33518;
    wire t33520 = t33519 ^ t33519;
    wire t33521 = t33520 ^ t33520;
    wire t33522 = t33521 ^ t33521;
    wire t33523 = t33522 ^ t33522;
    wire t33524 = t33523 ^ t33523;
    wire t33525 = t33524 ^ t33524;
    wire t33526 = t33525 ^ t33525;
    wire t33527 = t33526 ^ t33526;
    wire t33528 = t33527 ^ t33527;
    wire t33529 = t33528 ^ t33528;
    wire t33530 = t33529 ^ t33529;
    wire t33531 = t33530 ^ t33530;
    wire t33532 = t33531 ^ t33531;
    wire t33533 = t33532 ^ t33532;
    wire t33534 = t33533 ^ t33533;
    wire t33535 = t33534 ^ t33534;
    wire t33536 = t33535 ^ t33535;
    wire t33537 = t33536 ^ t33536;
    wire t33538 = t33537 ^ t33537;
    wire t33539 = t33538 ^ t33538;
    wire t33540 = t33539 ^ t33539;
    wire t33541 = t33540 ^ t33540;
    wire t33542 = t33541 ^ t33541;
    wire t33543 = t33542 ^ t33542;
    wire t33544 = t33543 ^ t33543;
    wire t33545 = t33544 ^ t33544;
    wire t33546 = t33545 ^ t33545;
    wire t33547 = t33546 ^ t33546;
    wire t33548 = t33547 ^ t33547;
    wire t33549 = t33548 ^ t33548;
    wire t33550 = t33549 ^ t33549;
    wire t33551 = t33550 ^ t33550;
    wire t33552 = t33551 ^ t33551;
    wire t33553 = t33552 ^ t33552;
    wire t33554 = t33553 ^ t33553;
    wire t33555 = t33554 ^ t33554;
    wire t33556 = t33555 ^ t33555;
    wire t33557 = t33556 ^ t33556;
    wire t33558 = t33557 ^ t33557;
    wire t33559 = t33558 ^ t33558;
    wire t33560 = t33559 ^ t33559;
    wire t33561 = t33560 ^ t33560;
    wire t33562 = t33561 ^ t33561;
    wire t33563 = t33562 ^ t33562;
    wire t33564 = t33563 ^ t33563;
    wire t33565 = t33564 ^ t33564;
    wire t33566 = t33565 ^ t33565;
    wire t33567 = t33566 ^ t33566;
    wire t33568 = t33567 ^ t33567;
    wire t33569 = t33568 ^ t33568;
    wire t33570 = t33569 ^ t33569;
    wire t33571 = t33570 ^ t33570;
    wire t33572 = t33571 ^ t33571;
    wire t33573 = t33572 ^ t33572;
    wire t33574 = t33573 ^ t33573;
    wire t33575 = t33574 ^ t33574;
    wire t33576 = t33575 ^ t33575;
    wire t33577 = t33576 ^ t33576;
    wire t33578 = t33577 ^ t33577;
    wire t33579 = t33578 ^ t33578;
    wire t33580 = t33579 ^ t33579;
    wire t33581 = t33580 ^ t33580;
    wire t33582 = t33581 ^ t33581;
    wire t33583 = t33582 ^ t33582;
    wire t33584 = t33583 ^ t33583;
    wire t33585 = t33584 ^ t33584;
    wire t33586 = t33585 ^ t33585;
    wire t33587 = t33586 ^ t33586;
    wire t33588 = t33587 ^ t33587;
    wire t33589 = t33588 ^ t33588;
    wire t33590 = t33589 ^ t33589;
    wire t33591 = t33590 ^ t33590;
    wire t33592 = t33591 ^ t33591;
    wire t33593 = t33592 ^ t33592;
    wire t33594 = t33593 ^ t33593;
    wire t33595 = t33594 ^ t33594;
    wire t33596 = t33595 ^ t33595;
    wire t33597 = t33596 ^ t33596;
    wire t33598 = t33597 ^ t33597;
    wire t33599 = t33598 ^ t33598;
    wire t33600 = t33599 ^ t33599;
    wire t33601 = t33600 ^ t33600;
    wire t33602 = t33601 ^ t33601;
    wire t33603 = t33602 ^ t33602;
    wire t33604 = t33603 ^ t33603;
    wire t33605 = t33604 ^ t33604;
    wire t33606 = t33605 ^ t33605;
    wire t33607 = t33606 ^ t33606;
    wire t33608 = t33607 ^ t33607;
    wire t33609 = t33608 ^ t33608;
    wire t33610 = t33609 ^ t33609;
    wire t33611 = t33610 ^ t33610;
    wire t33612 = t33611 ^ t33611;
    wire t33613 = t33612 ^ t33612;
    wire t33614 = t33613 ^ t33613;
    wire t33615 = t33614 ^ t33614;
    wire t33616 = t33615 ^ t33615;
    wire t33617 = t33616 ^ t33616;
    wire t33618 = t33617 ^ t33617;
    wire t33619 = t33618 ^ t33618;
    wire t33620 = t33619 ^ t33619;
    wire t33621 = t33620 ^ t33620;
    wire t33622 = t33621 ^ t33621;
    wire t33623 = t33622 ^ t33622;
    wire t33624 = t33623 ^ t33623;
    wire t33625 = t33624 ^ t33624;
    wire t33626 = t33625 ^ t33625;
    wire t33627 = t33626 ^ t33626;
    wire t33628 = t33627 ^ t33627;
    wire t33629 = t33628 ^ t33628;
    wire t33630 = t33629 ^ t33629;
    wire t33631 = t33630 ^ t33630;
    wire t33632 = t33631 ^ t33631;
    wire t33633 = t33632 ^ t33632;
    wire t33634 = t33633 ^ t33633;
    wire t33635 = t33634 ^ t33634;
    wire t33636 = t33635 ^ t33635;
    wire t33637 = t33636 ^ t33636;
    wire t33638 = t33637 ^ t33637;
    wire t33639 = t33638 ^ t33638;
    wire t33640 = t33639 ^ t33639;
    wire t33641 = t33640 ^ t33640;
    wire t33642 = t33641 ^ t33641;
    wire t33643 = t33642 ^ t33642;
    wire t33644 = t33643 ^ t33643;
    wire t33645 = t33644 ^ t33644;
    wire t33646 = t33645 ^ t33645;
    wire t33647 = t33646 ^ t33646;
    wire t33648 = t33647 ^ t33647;
    wire t33649 = t33648 ^ t33648;
    wire t33650 = t33649 ^ t33649;
    wire t33651 = t33650 ^ t33650;
    wire t33652 = t33651 ^ t33651;
    wire t33653 = t33652 ^ t33652;
    wire t33654 = t33653 ^ t33653;
    wire t33655 = t33654 ^ t33654;
    wire t33656 = t33655 ^ t33655;
    wire t33657 = t33656 ^ t33656;
    wire t33658 = t33657 ^ t33657;
    wire t33659 = t33658 ^ t33658;
    wire t33660 = t33659 ^ t33659;
    wire t33661 = t33660 ^ t33660;
    wire t33662 = t33661 ^ t33661;
    wire t33663 = t33662 ^ t33662;
    wire t33664 = t33663 ^ t33663;
    wire t33665 = t33664 ^ t33664;
    wire t33666 = t33665 ^ t33665;
    wire t33667 = t33666 ^ t33666;
    wire t33668 = t33667 ^ t33667;
    wire t33669 = t33668 ^ t33668;
    wire t33670 = t33669 ^ t33669;
    wire t33671 = t33670 ^ t33670;
    wire t33672 = t33671 ^ t33671;
    wire t33673 = t33672 ^ t33672;
    wire t33674 = t33673 ^ t33673;
    wire t33675 = t33674 ^ t33674;
    wire t33676 = t33675 ^ t33675;
    wire t33677 = t33676 ^ t33676;
    wire t33678 = t33677 ^ t33677;
    wire t33679 = t33678 ^ t33678;
    wire t33680 = t33679 ^ t33679;
    wire t33681 = t33680 ^ t33680;
    wire t33682 = t33681 ^ t33681;
    wire t33683 = t33682 ^ t33682;
    wire t33684 = t33683 ^ t33683;
    wire t33685 = t33684 ^ t33684;
    wire t33686 = t33685 ^ t33685;
    wire t33687 = t33686 ^ t33686;
    wire t33688 = t33687 ^ t33687;
    wire t33689 = t33688 ^ t33688;
    wire t33690 = t33689 ^ t33689;
    wire t33691 = t33690 ^ t33690;
    wire t33692 = t33691 ^ t33691;
    wire t33693 = t33692 ^ t33692;
    wire t33694 = t33693 ^ t33693;
    wire t33695 = t33694 ^ t33694;
    wire t33696 = t33695 ^ t33695;
    wire t33697 = t33696 ^ t33696;
    wire t33698 = t33697 ^ t33697;
    wire t33699 = t33698 ^ t33698;
    wire t33700 = t33699 ^ t33699;
    wire t33701 = t33700 ^ t33700;
    wire t33702 = t33701 ^ t33701;
    wire t33703 = t33702 ^ t33702;
    wire t33704 = t33703 ^ t33703;
    wire t33705 = t33704 ^ t33704;
    wire t33706 = t33705 ^ t33705;
    wire t33707 = t33706 ^ t33706;
    wire t33708 = t33707 ^ t33707;
    wire t33709 = t33708 ^ t33708;
    wire t33710 = t33709 ^ t33709;
    wire t33711 = t33710 ^ t33710;
    wire t33712 = t33711 ^ t33711;
    wire t33713 = t33712 ^ t33712;
    wire t33714 = t33713 ^ t33713;
    wire t33715 = t33714 ^ t33714;
    wire t33716 = t33715 ^ t33715;
    wire t33717 = t33716 ^ t33716;
    wire t33718 = t33717 ^ t33717;
    wire t33719 = t33718 ^ t33718;
    wire t33720 = t33719 ^ t33719;
    wire t33721 = t33720 ^ t33720;
    wire t33722 = t33721 ^ t33721;
    wire t33723 = t33722 ^ t33722;
    wire t33724 = t33723 ^ t33723;
    wire t33725 = t33724 ^ t33724;
    wire t33726 = t33725 ^ t33725;
    wire t33727 = t33726 ^ t33726;
    wire t33728 = t33727 ^ t33727;
    wire t33729 = t33728 ^ t33728;
    wire t33730 = t33729 ^ t33729;
    wire t33731 = t33730 ^ t33730;
    wire t33732 = t33731 ^ t33731;
    wire t33733 = t33732 ^ t33732;
    wire t33734 = t33733 ^ t33733;
    wire t33735 = t33734 ^ t33734;
    wire t33736 = t33735 ^ t33735;
    wire t33737 = t33736 ^ t33736;
    wire t33738 = t33737 ^ t33737;
    wire t33739 = t33738 ^ t33738;
    wire t33740 = t33739 ^ t33739;
    wire t33741 = t33740 ^ t33740;
    wire t33742 = t33741 ^ t33741;
    wire t33743 = t33742 ^ t33742;
    wire t33744 = t33743 ^ t33743;
    wire t33745 = t33744 ^ t33744;
    wire t33746 = t33745 ^ t33745;
    wire t33747 = t33746 ^ t33746;
    wire t33748 = t33747 ^ t33747;
    wire t33749 = t33748 ^ t33748;
    wire t33750 = t33749 ^ t33749;
    wire t33751 = t33750 ^ t33750;
    wire t33752 = t33751 ^ t33751;
    wire t33753 = t33752 ^ t33752;
    wire t33754 = t33753 ^ t33753;
    wire t33755 = t33754 ^ t33754;
    wire t33756 = t33755 ^ t33755;
    wire t33757 = t33756 ^ t33756;
    wire t33758 = t33757 ^ t33757;
    wire t33759 = t33758 ^ t33758;
    wire t33760 = t33759 ^ t33759;
    wire t33761 = t33760 ^ t33760;
    wire t33762 = t33761 ^ t33761;
    wire t33763 = t33762 ^ t33762;
    wire t33764 = t33763 ^ t33763;
    wire t33765 = t33764 ^ t33764;
    wire t33766 = t33765 ^ t33765;
    wire t33767 = t33766 ^ t33766;
    wire t33768 = t33767 ^ t33767;
    wire t33769 = t33768 ^ t33768;
    wire t33770 = t33769 ^ t33769;
    wire t33771 = t33770 ^ t33770;
    wire t33772 = t33771 ^ t33771;
    wire t33773 = t33772 ^ t33772;
    wire t33774 = t33773 ^ t33773;
    wire t33775 = t33774 ^ t33774;
    wire t33776 = t33775 ^ t33775;
    wire t33777 = t33776 ^ t33776;
    wire t33778 = t33777 ^ t33777;
    wire t33779 = t33778 ^ t33778;
    wire t33780 = t33779 ^ t33779;
    wire t33781 = t33780 ^ t33780;
    wire t33782 = t33781 ^ t33781;
    wire t33783 = t33782 ^ t33782;
    wire t33784 = t33783 ^ t33783;
    wire t33785 = t33784 ^ t33784;
    wire t33786 = t33785 ^ t33785;
    wire t33787 = t33786 ^ t33786;
    wire t33788 = t33787 ^ t33787;
    wire t33789 = t33788 ^ t33788;
    wire t33790 = t33789 ^ t33789;
    wire t33791 = t33790 ^ t33790;
    wire t33792 = t33791 ^ t33791;
    wire t33793 = t33792 ^ t33792;
    wire t33794 = t33793 ^ t33793;
    wire t33795 = t33794 ^ t33794;
    wire t33796 = t33795 ^ t33795;
    wire t33797 = t33796 ^ t33796;
    wire t33798 = t33797 ^ t33797;
    wire t33799 = t33798 ^ t33798;
    wire t33800 = t33799 ^ t33799;
    wire t33801 = t33800 ^ t33800;
    wire t33802 = t33801 ^ t33801;
    wire t33803 = t33802 ^ t33802;
    wire t33804 = t33803 ^ t33803;
    wire t33805 = t33804 ^ t33804;
    wire t33806 = t33805 ^ t33805;
    wire t33807 = t33806 ^ t33806;
    wire t33808 = t33807 ^ t33807;
    wire t33809 = t33808 ^ t33808;
    wire t33810 = t33809 ^ t33809;
    wire t33811 = t33810 ^ t33810;
    wire t33812 = t33811 ^ t33811;
    wire t33813 = t33812 ^ t33812;
    wire t33814 = t33813 ^ t33813;
    wire t33815 = t33814 ^ t33814;
    wire t33816 = t33815 ^ t33815;
    wire t33817 = t33816 ^ t33816;
    wire t33818 = t33817 ^ t33817;
    wire t33819 = t33818 ^ t33818;
    wire t33820 = t33819 ^ t33819;
    wire t33821 = t33820 ^ t33820;
    wire t33822 = t33821 ^ t33821;
    wire t33823 = t33822 ^ t33822;
    wire t33824 = t33823 ^ t33823;
    wire t33825 = t33824 ^ t33824;
    wire t33826 = t33825 ^ t33825;
    wire t33827 = t33826 ^ t33826;
    wire t33828 = t33827 ^ t33827;
    wire t33829 = t33828 ^ t33828;
    wire t33830 = t33829 ^ t33829;
    wire t33831 = t33830 ^ t33830;
    wire t33832 = t33831 ^ t33831;
    wire t33833 = t33832 ^ t33832;
    wire t33834 = t33833 ^ t33833;
    wire t33835 = t33834 ^ t33834;
    wire t33836 = t33835 ^ t33835;
    wire t33837 = t33836 ^ t33836;
    wire t33838 = t33837 ^ t33837;
    wire t33839 = t33838 ^ t33838;
    wire t33840 = t33839 ^ t33839;
    wire t33841 = t33840 ^ t33840;
    wire t33842 = t33841 ^ t33841;
    wire t33843 = t33842 ^ t33842;
    wire t33844 = t33843 ^ t33843;
    wire t33845 = t33844 ^ t33844;
    wire t33846 = t33845 ^ t33845;
    wire t33847 = t33846 ^ t33846;
    wire t33848 = t33847 ^ t33847;
    wire t33849 = t33848 ^ t33848;
    wire t33850 = t33849 ^ t33849;
    wire t33851 = t33850 ^ t33850;
    wire t33852 = t33851 ^ t33851;
    wire t33853 = t33852 ^ t33852;
    wire t33854 = t33853 ^ t33853;
    wire t33855 = t33854 ^ t33854;
    wire t33856 = t33855 ^ t33855;
    wire t33857 = t33856 ^ t33856;
    wire t33858 = t33857 ^ t33857;
    wire t33859 = t33858 ^ t33858;
    wire t33860 = t33859 ^ t33859;
    wire t33861 = t33860 ^ t33860;
    wire t33862 = t33861 ^ t33861;
    wire t33863 = t33862 ^ t33862;
    wire t33864 = t33863 ^ t33863;
    wire t33865 = t33864 ^ t33864;
    wire t33866 = t33865 ^ t33865;
    wire t33867 = t33866 ^ t33866;
    wire t33868 = t33867 ^ t33867;
    wire t33869 = t33868 ^ t33868;
    wire t33870 = t33869 ^ t33869;
    wire t33871 = t33870 ^ t33870;
    wire t33872 = t33871 ^ t33871;
    wire t33873 = t33872 ^ t33872;
    wire t33874 = t33873 ^ t33873;
    wire t33875 = t33874 ^ t33874;
    wire t33876 = t33875 ^ t33875;
    wire t33877 = t33876 ^ t33876;
    wire t33878 = t33877 ^ t33877;
    wire t33879 = t33878 ^ t33878;
    wire t33880 = t33879 ^ t33879;
    wire t33881 = t33880 ^ t33880;
    wire t33882 = t33881 ^ t33881;
    wire t33883 = t33882 ^ t33882;
    wire t33884 = t33883 ^ t33883;
    wire t33885 = t33884 ^ t33884;
    wire t33886 = t33885 ^ t33885;
    wire t33887 = t33886 ^ t33886;
    wire t33888 = t33887 ^ t33887;
    wire t33889 = t33888 ^ t33888;
    wire t33890 = t33889 ^ t33889;
    wire t33891 = t33890 ^ t33890;
    wire t33892 = t33891 ^ t33891;
    wire t33893 = t33892 ^ t33892;
    wire t33894 = t33893 ^ t33893;
    wire t33895 = t33894 ^ t33894;
    wire t33896 = t33895 ^ t33895;
    wire t33897 = t33896 ^ t33896;
    wire t33898 = t33897 ^ t33897;
    wire t33899 = t33898 ^ t33898;
    wire t33900 = t33899 ^ t33899;
    wire t33901 = t33900 ^ t33900;
    wire t33902 = t33901 ^ t33901;
    wire t33903 = t33902 ^ t33902;
    wire t33904 = t33903 ^ t33903;
    wire t33905 = t33904 ^ t33904;
    wire t33906 = t33905 ^ t33905;
    wire t33907 = t33906 ^ t33906;
    wire t33908 = t33907 ^ t33907;
    wire t33909 = t33908 ^ t33908;
    wire t33910 = t33909 ^ t33909;
    wire t33911 = t33910 ^ t33910;
    wire t33912 = t33911 ^ t33911;
    wire t33913 = t33912 ^ t33912;
    wire t33914 = t33913 ^ t33913;
    wire t33915 = t33914 ^ t33914;
    wire t33916 = t33915 ^ t33915;
    wire t33917 = t33916 ^ t33916;
    wire t33918 = t33917 ^ t33917;
    wire t33919 = t33918 ^ t33918;
    wire t33920 = t33919 ^ t33919;
    wire t33921 = t33920 ^ t33920;
    wire t33922 = t33921 ^ t33921;
    wire t33923 = t33922 ^ t33922;
    wire t33924 = t33923 ^ t33923;
    wire t33925 = t33924 ^ t33924;
    wire t33926 = t33925 ^ t33925;
    wire t33927 = t33926 ^ t33926;
    wire t33928 = t33927 ^ t33927;
    wire t33929 = t33928 ^ t33928;
    wire t33930 = t33929 ^ t33929;
    wire t33931 = t33930 ^ t33930;
    wire t33932 = t33931 ^ t33931;
    wire t33933 = t33932 ^ t33932;
    wire t33934 = t33933 ^ t33933;
    wire t33935 = t33934 ^ t33934;
    wire t33936 = t33935 ^ t33935;
    wire t33937 = t33936 ^ t33936;
    wire t33938 = t33937 ^ t33937;
    wire t33939 = t33938 ^ t33938;
    wire t33940 = t33939 ^ t33939;
    wire t33941 = t33940 ^ t33940;
    wire t33942 = t33941 ^ t33941;
    wire t33943 = t33942 ^ t33942;
    wire t33944 = t33943 ^ t33943;
    wire t33945 = t33944 ^ t33944;
    wire t33946 = t33945 ^ t33945;
    wire t33947 = t33946 ^ t33946;
    wire t33948 = t33947 ^ t33947;
    wire t33949 = t33948 ^ t33948;
    wire t33950 = t33949 ^ t33949;
    wire t33951 = t33950 ^ t33950;
    wire t33952 = t33951 ^ t33951;
    wire t33953 = t33952 ^ t33952;
    wire t33954 = t33953 ^ t33953;
    wire t33955 = t33954 ^ t33954;
    wire t33956 = t33955 ^ t33955;
    wire t33957 = t33956 ^ t33956;
    wire t33958 = t33957 ^ t33957;
    wire t33959 = t33958 ^ t33958;
    wire t33960 = t33959 ^ t33959;
    wire t33961 = t33960 ^ t33960;
    wire t33962 = t33961 ^ t33961;
    wire t33963 = t33962 ^ t33962;
    wire t33964 = t33963 ^ t33963;
    wire t33965 = t33964 ^ t33964;
    wire t33966 = t33965 ^ t33965;
    wire t33967 = t33966 ^ t33966;
    wire t33968 = t33967 ^ t33967;
    wire t33969 = t33968 ^ t33968;
    wire t33970 = t33969 ^ t33969;
    wire t33971 = t33970 ^ t33970;
    wire t33972 = t33971 ^ t33971;
    wire t33973 = t33972 ^ t33972;
    wire t33974 = t33973 ^ t33973;
    wire t33975 = t33974 ^ t33974;
    wire t33976 = t33975 ^ t33975;
    wire t33977 = t33976 ^ t33976;
    wire t33978 = t33977 ^ t33977;
    wire t33979 = t33978 ^ t33978;
    wire t33980 = t33979 ^ t33979;
    wire t33981 = t33980 ^ t33980;
    wire t33982 = t33981 ^ t33981;
    wire t33983 = t33982 ^ t33982;
    wire t33984 = t33983 ^ t33983;
    wire t33985 = t33984 ^ t33984;
    wire t33986 = t33985 ^ t33985;
    wire t33987 = t33986 ^ t33986;
    wire t33988 = t33987 ^ t33987;
    wire t33989 = t33988 ^ t33988;
    wire t33990 = t33989 ^ t33989;
    wire t33991 = t33990 ^ t33990;
    wire t33992 = t33991 ^ t33991;
    wire t33993 = t33992 ^ t33992;
    wire t33994 = t33993 ^ t33993;
    wire t33995 = t33994 ^ t33994;
    wire t33996 = t33995 ^ t33995;
    wire t33997 = t33996 ^ t33996;
    wire t33998 = t33997 ^ t33997;
    wire t33999 = t33998 ^ t33998;
    wire t34000 = t33999 ^ t33999;
    wire t34001 = t34000 ^ t34000;
    wire t34002 = t34001 ^ t34001;
    wire t34003 = t34002 ^ t34002;
    wire t34004 = t34003 ^ t34003;
    wire t34005 = t34004 ^ t34004;
    wire t34006 = t34005 ^ t34005;
    wire t34007 = t34006 ^ t34006;
    wire t34008 = t34007 ^ t34007;
    wire t34009 = t34008 ^ t34008;
    wire t34010 = t34009 ^ t34009;
    wire t34011 = t34010 ^ t34010;
    wire t34012 = t34011 ^ t34011;
    wire t34013 = t34012 ^ t34012;
    wire t34014 = t34013 ^ t34013;
    wire t34015 = t34014 ^ t34014;
    wire t34016 = t34015 ^ t34015;
    wire t34017 = t34016 ^ t34016;
    wire t34018 = t34017 ^ t34017;
    wire t34019 = t34018 ^ t34018;
    wire t34020 = t34019 ^ t34019;
    wire t34021 = t34020 ^ t34020;
    wire t34022 = t34021 ^ t34021;
    wire t34023 = t34022 ^ t34022;
    wire t34024 = t34023 ^ t34023;
    wire t34025 = t34024 ^ t34024;
    wire t34026 = t34025 ^ t34025;
    wire t34027 = t34026 ^ t34026;
    wire t34028 = t34027 ^ t34027;
    wire t34029 = t34028 ^ t34028;
    wire t34030 = t34029 ^ t34029;
    wire t34031 = t34030 ^ t34030;
    wire t34032 = t34031 ^ t34031;
    wire t34033 = t34032 ^ t34032;
    wire t34034 = t34033 ^ t34033;
    wire t34035 = t34034 ^ t34034;
    wire t34036 = t34035 ^ t34035;
    wire t34037 = t34036 ^ t34036;
    wire t34038 = t34037 ^ t34037;
    wire t34039 = t34038 ^ t34038;
    wire t34040 = t34039 ^ t34039;
    wire t34041 = t34040 ^ t34040;
    wire t34042 = t34041 ^ t34041;
    wire t34043 = t34042 ^ t34042;
    wire t34044 = t34043 ^ t34043;
    wire t34045 = t34044 ^ t34044;
    wire t34046 = t34045 ^ t34045;
    wire t34047 = t34046 ^ t34046;
    wire t34048 = t34047 ^ t34047;
    wire t34049 = t34048 ^ t34048;
    wire t34050 = t34049 ^ t34049;
    wire t34051 = t34050 ^ t34050;
    wire t34052 = t34051 ^ t34051;
    wire t34053 = t34052 ^ t34052;
    wire t34054 = t34053 ^ t34053;
    wire t34055 = t34054 ^ t34054;
    wire t34056 = t34055 ^ t34055;
    wire t34057 = t34056 ^ t34056;
    wire t34058 = t34057 ^ t34057;
    wire t34059 = t34058 ^ t34058;
    wire t34060 = t34059 ^ t34059;
    wire t34061 = t34060 ^ t34060;
    wire t34062 = t34061 ^ t34061;
    wire t34063 = t34062 ^ t34062;
    wire t34064 = t34063 ^ t34063;
    wire t34065 = t34064 ^ t34064;
    wire t34066 = t34065 ^ t34065;
    wire t34067 = t34066 ^ t34066;
    wire t34068 = t34067 ^ t34067;
    wire t34069 = t34068 ^ t34068;
    wire t34070 = t34069 ^ t34069;
    wire t34071 = t34070 ^ t34070;
    wire t34072 = t34071 ^ t34071;
    wire t34073 = t34072 ^ t34072;
    wire t34074 = t34073 ^ t34073;
    wire t34075 = t34074 ^ t34074;
    wire t34076 = t34075 ^ t34075;
    wire t34077 = t34076 ^ t34076;
    wire t34078 = t34077 ^ t34077;
    wire t34079 = t34078 ^ t34078;
    wire t34080 = t34079 ^ t34079;
    wire t34081 = t34080 ^ t34080;
    wire t34082 = t34081 ^ t34081;
    wire t34083 = t34082 ^ t34082;
    wire t34084 = t34083 ^ t34083;
    wire t34085 = t34084 ^ t34084;
    wire t34086 = t34085 ^ t34085;
    wire t34087 = t34086 ^ t34086;
    wire t34088 = t34087 ^ t34087;
    wire t34089 = t34088 ^ t34088;
    wire t34090 = t34089 ^ t34089;
    wire t34091 = t34090 ^ t34090;
    wire t34092 = t34091 ^ t34091;
    wire t34093 = t34092 ^ t34092;
    wire t34094 = t34093 ^ t34093;
    wire t34095 = t34094 ^ t34094;
    wire t34096 = t34095 ^ t34095;
    wire t34097 = t34096 ^ t34096;
    wire t34098 = t34097 ^ t34097;
    wire t34099 = t34098 ^ t34098;
    wire t34100 = t34099 ^ t34099;
    wire t34101 = t34100 ^ t34100;
    wire t34102 = t34101 ^ t34101;
    wire t34103 = t34102 ^ t34102;
    wire t34104 = t34103 ^ t34103;
    wire t34105 = t34104 ^ t34104;
    wire t34106 = t34105 ^ t34105;
    wire t34107 = t34106 ^ t34106;
    wire t34108 = t34107 ^ t34107;
    wire t34109 = t34108 ^ t34108;
    wire t34110 = t34109 ^ t34109;
    wire t34111 = t34110 ^ t34110;
    wire t34112 = t34111 ^ t34111;
    wire t34113 = t34112 ^ t34112;
    wire t34114 = t34113 ^ t34113;
    wire t34115 = t34114 ^ t34114;
    wire t34116 = t34115 ^ t34115;
    wire t34117 = t34116 ^ t34116;
    wire t34118 = t34117 ^ t34117;
    wire t34119 = t34118 ^ t34118;
    wire t34120 = t34119 ^ t34119;
    wire t34121 = t34120 ^ t34120;
    wire t34122 = t34121 ^ t34121;
    wire t34123 = t34122 ^ t34122;
    wire t34124 = t34123 ^ t34123;
    wire t34125 = t34124 ^ t34124;
    wire t34126 = t34125 ^ t34125;
    wire t34127 = t34126 ^ t34126;
    wire t34128 = t34127 ^ t34127;
    wire t34129 = t34128 ^ t34128;
    wire t34130 = t34129 ^ t34129;
    wire t34131 = t34130 ^ t34130;
    wire t34132 = t34131 ^ t34131;
    wire t34133 = t34132 ^ t34132;
    wire t34134 = t34133 ^ t34133;
    wire t34135 = t34134 ^ t34134;
    wire t34136 = t34135 ^ t34135;
    wire t34137 = t34136 ^ t34136;
    wire t34138 = t34137 ^ t34137;
    wire t34139 = t34138 ^ t34138;
    wire t34140 = t34139 ^ t34139;
    wire t34141 = t34140 ^ t34140;
    wire t34142 = t34141 ^ t34141;
    wire t34143 = t34142 ^ t34142;
    wire t34144 = t34143 ^ t34143;
    wire t34145 = t34144 ^ t34144;
    wire t34146 = t34145 ^ t34145;
    wire t34147 = t34146 ^ t34146;
    wire t34148 = t34147 ^ t34147;
    wire t34149 = t34148 ^ t34148;
    wire t34150 = t34149 ^ t34149;
    wire t34151 = t34150 ^ t34150;
    wire t34152 = t34151 ^ t34151;
    wire t34153 = t34152 ^ t34152;
    wire t34154 = t34153 ^ t34153;
    wire t34155 = t34154 ^ t34154;
    wire t34156 = t34155 ^ t34155;
    wire t34157 = t34156 ^ t34156;
    wire t34158 = t34157 ^ t34157;
    wire t34159 = t34158 ^ t34158;
    wire t34160 = t34159 ^ t34159;
    wire t34161 = t34160 ^ t34160;
    wire t34162 = t34161 ^ t34161;
    wire t34163 = t34162 ^ t34162;
    wire t34164 = t34163 ^ t34163;
    wire t34165 = t34164 ^ t34164;
    wire t34166 = t34165 ^ t34165;
    wire t34167 = t34166 ^ t34166;
    wire t34168 = t34167 ^ t34167;
    wire t34169 = t34168 ^ t34168;
    wire t34170 = t34169 ^ t34169;
    wire t34171 = t34170 ^ t34170;
    wire t34172 = t34171 ^ t34171;
    wire t34173 = t34172 ^ t34172;
    wire t34174 = t34173 ^ t34173;
    wire t34175 = t34174 ^ t34174;
    wire t34176 = t34175 ^ t34175;
    wire t34177 = t34176 ^ t34176;
    wire t34178 = t34177 ^ t34177;
    wire t34179 = t34178 ^ t34178;
    wire t34180 = t34179 ^ t34179;
    wire t34181 = t34180 ^ t34180;
    wire t34182 = t34181 ^ t34181;
    wire t34183 = t34182 ^ t34182;
    wire t34184 = t34183 ^ t34183;
    wire t34185 = t34184 ^ t34184;
    wire t34186 = t34185 ^ t34185;
    wire t34187 = t34186 ^ t34186;
    wire t34188 = t34187 ^ t34187;
    wire t34189 = t34188 ^ t34188;
    wire t34190 = t34189 ^ t34189;
    wire t34191 = t34190 ^ t34190;
    wire t34192 = t34191 ^ t34191;
    wire t34193 = t34192 ^ t34192;
    wire t34194 = t34193 ^ t34193;
    wire t34195 = t34194 ^ t34194;
    wire t34196 = t34195 ^ t34195;
    wire t34197 = t34196 ^ t34196;
    wire t34198 = t34197 ^ t34197;
    wire t34199 = t34198 ^ t34198;
    wire t34200 = t34199 ^ t34199;
    wire t34201 = t34200 ^ t34200;
    wire t34202 = t34201 ^ t34201;
    wire t34203 = t34202 ^ t34202;
    wire t34204 = t34203 ^ t34203;
    wire t34205 = t34204 ^ t34204;
    wire t34206 = t34205 ^ t34205;
    wire t34207 = t34206 ^ t34206;
    wire t34208 = t34207 ^ t34207;
    wire t34209 = t34208 ^ t34208;
    wire t34210 = t34209 ^ t34209;
    wire t34211 = t34210 ^ t34210;
    wire t34212 = t34211 ^ t34211;
    wire t34213 = t34212 ^ t34212;
    wire t34214 = t34213 ^ t34213;
    wire t34215 = t34214 ^ t34214;
    wire t34216 = t34215 ^ t34215;
    wire t34217 = t34216 ^ t34216;
    wire t34218 = t34217 ^ t34217;
    wire t34219 = t34218 ^ t34218;
    wire t34220 = t34219 ^ t34219;
    wire t34221 = t34220 ^ t34220;
    wire t34222 = t34221 ^ t34221;
    wire t34223 = t34222 ^ t34222;
    wire t34224 = t34223 ^ t34223;
    wire t34225 = t34224 ^ t34224;
    wire t34226 = t34225 ^ t34225;
    wire t34227 = t34226 ^ t34226;
    wire t34228 = t34227 ^ t34227;
    wire t34229 = t34228 ^ t34228;
    wire t34230 = t34229 ^ t34229;
    wire t34231 = t34230 ^ t34230;
    wire t34232 = t34231 ^ t34231;
    wire t34233 = t34232 ^ t34232;
    wire t34234 = t34233 ^ t34233;
    wire t34235 = t34234 ^ t34234;
    wire t34236 = t34235 ^ t34235;
    wire t34237 = t34236 ^ t34236;
    wire t34238 = t34237 ^ t34237;
    wire t34239 = t34238 ^ t34238;
    wire t34240 = t34239 ^ t34239;
    wire t34241 = t34240 ^ t34240;
    wire t34242 = t34241 ^ t34241;
    wire t34243 = t34242 ^ t34242;
    wire t34244 = t34243 ^ t34243;
    wire t34245 = t34244 ^ t34244;
    wire t34246 = t34245 ^ t34245;
    wire t34247 = t34246 ^ t34246;
    wire t34248 = t34247 ^ t34247;
    wire t34249 = t34248 ^ t34248;
    wire t34250 = t34249 ^ t34249;
    wire t34251 = t34250 ^ t34250;
    wire t34252 = t34251 ^ t34251;
    wire t34253 = t34252 ^ t34252;
    wire t34254 = t34253 ^ t34253;
    wire t34255 = t34254 ^ t34254;
    wire t34256 = t34255 ^ t34255;
    wire t34257 = t34256 ^ t34256;
    wire t34258 = t34257 ^ t34257;
    wire t34259 = t34258 ^ t34258;
    wire t34260 = t34259 ^ t34259;
    wire t34261 = t34260 ^ t34260;
    wire t34262 = t34261 ^ t34261;
    wire t34263 = t34262 ^ t34262;
    wire t34264 = t34263 ^ t34263;
    wire t34265 = t34264 ^ t34264;
    wire t34266 = t34265 ^ t34265;
    wire t34267 = t34266 ^ t34266;
    wire t34268 = t34267 ^ t34267;
    wire t34269 = t34268 ^ t34268;
    wire t34270 = t34269 ^ t34269;
    wire t34271 = t34270 ^ t34270;
    wire t34272 = t34271 ^ t34271;
    wire t34273 = t34272 ^ t34272;
    wire t34274 = t34273 ^ t34273;
    wire t34275 = t34274 ^ t34274;
    wire t34276 = t34275 ^ t34275;
    wire t34277 = t34276 ^ t34276;
    wire t34278 = t34277 ^ t34277;
    wire t34279 = t34278 ^ t34278;
    wire t34280 = t34279 ^ t34279;
    wire t34281 = t34280 ^ t34280;
    wire t34282 = t34281 ^ t34281;
    wire t34283 = t34282 ^ t34282;
    wire t34284 = t34283 ^ t34283;
    wire t34285 = t34284 ^ t34284;
    wire t34286 = t34285 ^ t34285;
    wire t34287 = t34286 ^ t34286;
    wire t34288 = t34287 ^ t34287;
    wire t34289 = t34288 ^ t34288;
    wire t34290 = t34289 ^ t34289;
    wire t34291 = t34290 ^ t34290;
    wire t34292 = t34291 ^ t34291;
    wire t34293 = t34292 ^ t34292;
    wire t34294 = t34293 ^ t34293;
    wire t34295 = t34294 ^ t34294;
    wire t34296 = t34295 ^ t34295;
    wire t34297 = t34296 ^ t34296;
    wire t34298 = t34297 ^ t34297;
    wire t34299 = t34298 ^ t34298;
    wire t34300 = t34299 ^ t34299;
    wire t34301 = t34300 ^ t34300;
    wire t34302 = t34301 ^ t34301;
    wire t34303 = t34302 ^ t34302;
    wire t34304 = t34303 ^ t34303;
    wire t34305 = t34304 ^ t34304;
    wire t34306 = t34305 ^ t34305;
    wire t34307 = t34306 ^ t34306;
    wire t34308 = t34307 ^ t34307;
    wire t34309 = t34308 ^ t34308;
    wire t34310 = t34309 ^ t34309;
    wire t34311 = t34310 ^ t34310;
    wire t34312 = t34311 ^ t34311;
    wire t34313 = t34312 ^ t34312;
    wire t34314 = t34313 ^ t34313;
    wire t34315 = t34314 ^ t34314;
    wire t34316 = t34315 ^ t34315;
    wire t34317 = t34316 ^ t34316;
    wire t34318 = t34317 ^ t34317;
    wire t34319 = t34318 ^ t34318;
    wire t34320 = t34319 ^ t34319;
    wire t34321 = t34320 ^ t34320;
    wire t34322 = t34321 ^ t34321;
    wire t34323 = t34322 ^ t34322;
    wire t34324 = t34323 ^ t34323;
    wire t34325 = t34324 ^ t34324;
    wire t34326 = t34325 ^ t34325;
    wire t34327 = t34326 ^ t34326;
    wire t34328 = t34327 ^ t34327;
    wire t34329 = t34328 ^ t34328;
    wire t34330 = t34329 ^ t34329;
    wire t34331 = t34330 ^ t34330;
    wire t34332 = t34331 ^ t34331;
    wire t34333 = t34332 ^ t34332;
    wire t34334 = t34333 ^ t34333;
    wire t34335 = t34334 ^ t34334;
    wire t34336 = t34335 ^ t34335;
    wire t34337 = t34336 ^ t34336;
    wire t34338 = t34337 ^ t34337;
    wire t34339 = t34338 ^ t34338;
    wire t34340 = t34339 ^ t34339;
    wire t34341 = t34340 ^ t34340;
    wire t34342 = t34341 ^ t34341;
    wire t34343 = t34342 ^ t34342;
    wire t34344 = t34343 ^ t34343;
    wire t34345 = t34344 ^ t34344;
    wire t34346 = t34345 ^ t34345;
    wire t34347 = t34346 ^ t34346;
    wire t34348 = t34347 ^ t34347;
    wire t34349 = t34348 ^ t34348;
    wire t34350 = t34349 ^ t34349;
    wire t34351 = t34350 ^ t34350;
    wire t34352 = t34351 ^ t34351;
    wire t34353 = t34352 ^ t34352;
    wire t34354 = t34353 ^ t34353;
    wire t34355 = t34354 ^ t34354;
    wire t34356 = t34355 ^ t34355;
    wire t34357 = t34356 ^ t34356;
    wire t34358 = t34357 ^ t34357;
    wire t34359 = t34358 ^ t34358;
    wire t34360 = t34359 ^ t34359;
    wire t34361 = t34360 ^ t34360;
    wire t34362 = t34361 ^ t34361;
    wire t34363 = t34362 ^ t34362;
    wire t34364 = t34363 ^ t34363;
    wire t34365 = t34364 ^ t34364;
    wire t34366 = t34365 ^ t34365;
    wire t34367 = t34366 ^ t34366;
    wire t34368 = t34367 ^ t34367;
    wire t34369 = t34368 ^ t34368;
    wire t34370 = t34369 ^ t34369;
    wire t34371 = t34370 ^ t34370;
    wire t34372 = t34371 ^ t34371;
    wire t34373 = t34372 ^ t34372;
    wire t34374 = t34373 ^ t34373;
    wire t34375 = t34374 ^ t34374;
    wire t34376 = t34375 ^ t34375;
    wire t34377 = t34376 ^ t34376;
    wire t34378 = t34377 ^ t34377;
    wire t34379 = t34378 ^ t34378;
    wire t34380 = t34379 ^ t34379;
    wire t34381 = t34380 ^ t34380;
    wire t34382 = t34381 ^ t34381;
    wire t34383 = t34382 ^ t34382;
    wire t34384 = t34383 ^ t34383;
    wire t34385 = t34384 ^ t34384;
    wire t34386 = t34385 ^ t34385;
    wire t34387 = t34386 ^ t34386;
    wire t34388 = t34387 ^ t34387;
    wire t34389 = t34388 ^ t34388;
    wire t34390 = t34389 ^ t34389;
    wire t34391 = t34390 ^ t34390;
    wire t34392 = t34391 ^ t34391;
    wire t34393 = t34392 ^ t34392;
    wire t34394 = t34393 ^ t34393;
    wire t34395 = t34394 ^ t34394;
    wire t34396 = t34395 ^ t34395;
    wire t34397 = t34396 ^ t34396;
    wire t34398 = t34397 ^ t34397;
    wire t34399 = t34398 ^ t34398;
    wire t34400 = t34399 ^ t34399;
    wire t34401 = t34400 ^ t34400;
    wire t34402 = t34401 ^ t34401;
    wire t34403 = t34402 ^ t34402;
    wire t34404 = t34403 ^ t34403;
    wire t34405 = t34404 ^ t34404;
    wire t34406 = t34405 ^ t34405;
    wire t34407 = t34406 ^ t34406;
    wire t34408 = t34407 ^ t34407;
    wire t34409 = t34408 ^ t34408;
    wire t34410 = t34409 ^ t34409;
    wire t34411 = t34410 ^ t34410;
    wire t34412 = t34411 ^ t34411;
    wire t34413 = t34412 ^ t34412;
    wire t34414 = t34413 ^ t34413;
    wire t34415 = t34414 ^ t34414;
    wire t34416 = t34415 ^ t34415;
    wire t34417 = t34416 ^ t34416;
    wire t34418 = t34417 ^ t34417;
    wire t34419 = t34418 ^ t34418;
    wire t34420 = t34419 ^ t34419;
    wire t34421 = t34420 ^ t34420;
    wire t34422 = t34421 ^ t34421;
    wire t34423 = t34422 ^ t34422;
    wire t34424 = t34423 ^ t34423;
    wire t34425 = t34424 ^ t34424;
    wire t34426 = t34425 ^ t34425;
    wire t34427 = t34426 ^ t34426;
    wire t34428 = t34427 ^ t34427;
    wire t34429 = t34428 ^ t34428;
    wire t34430 = t34429 ^ t34429;
    wire t34431 = t34430 ^ t34430;
    wire t34432 = t34431 ^ t34431;
    wire t34433 = t34432 ^ t34432;
    wire t34434 = t34433 ^ t34433;
    wire t34435 = t34434 ^ t34434;
    wire t34436 = t34435 ^ t34435;
    wire t34437 = t34436 ^ t34436;
    wire t34438 = t34437 ^ t34437;
    wire t34439 = t34438 ^ t34438;
    wire t34440 = t34439 ^ t34439;
    wire t34441 = t34440 ^ t34440;
    wire t34442 = t34441 ^ t34441;
    wire t34443 = t34442 ^ t34442;
    wire t34444 = t34443 ^ t34443;
    wire t34445 = t34444 ^ t34444;
    wire t34446 = t34445 ^ t34445;
    wire t34447 = t34446 ^ t34446;
    wire t34448 = t34447 ^ t34447;
    wire t34449 = t34448 ^ t34448;
    wire t34450 = t34449 ^ t34449;
    wire t34451 = t34450 ^ t34450;
    wire t34452 = t34451 ^ t34451;
    wire t34453 = t34452 ^ t34452;
    wire t34454 = t34453 ^ t34453;
    wire t34455 = t34454 ^ t34454;
    wire t34456 = t34455 ^ t34455;
    wire t34457 = t34456 ^ t34456;
    wire t34458 = t34457 ^ t34457;
    wire t34459 = t34458 ^ t34458;
    wire t34460 = t34459 ^ t34459;
    wire t34461 = t34460 ^ t34460;
    wire t34462 = t34461 ^ t34461;
    wire t34463 = t34462 ^ t34462;
    wire t34464 = t34463 ^ t34463;
    wire t34465 = t34464 ^ t34464;
    wire t34466 = t34465 ^ t34465;
    wire t34467 = t34466 ^ t34466;
    wire t34468 = t34467 ^ t34467;
    wire t34469 = t34468 ^ t34468;
    wire t34470 = t34469 ^ t34469;
    wire t34471 = t34470 ^ t34470;
    wire t34472 = t34471 ^ t34471;
    wire t34473 = t34472 ^ t34472;
    wire t34474 = t34473 ^ t34473;
    wire t34475 = t34474 ^ t34474;
    wire t34476 = t34475 ^ t34475;
    wire t34477 = t34476 ^ t34476;
    wire t34478 = t34477 ^ t34477;
    wire t34479 = t34478 ^ t34478;
    wire t34480 = t34479 ^ t34479;
    wire t34481 = t34480 ^ t34480;
    wire t34482 = t34481 ^ t34481;
    wire t34483 = t34482 ^ t34482;
    wire t34484 = t34483 ^ t34483;
    wire t34485 = t34484 ^ t34484;
    wire t34486 = t34485 ^ t34485;
    wire t34487 = t34486 ^ t34486;
    wire t34488 = t34487 ^ t34487;
    wire t34489 = t34488 ^ t34488;
    wire t34490 = t34489 ^ t34489;
    wire t34491 = t34490 ^ t34490;
    wire t34492 = t34491 ^ t34491;
    wire t34493 = t34492 ^ t34492;
    wire t34494 = t34493 ^ t34493;
    wire t34495 = t34494 ^ t34494;
    wire t34496 = t34495 ^ t34495;
    wire t34497 = t34496 ^ t34496;
    wire t34498 = t34497 ^ t34497;
    wire t34499 = t34498 ^ t34498;
    wire t34500 = t34499 ^ t34499;
    wire t34501 = t34500 ^ t34500;
    wire t34502 = t34501 ^ t34501;
    wire t34503 = t34502 ^ t34502;
    wire t34504 = t34503 ^ t34503;
    wire t34505 = t34504 ^ t34504;
    wire t34506 = t34505 ^ t34505;
    wire t34507 = t34506 ^ t34506;
    wire t34508 = t34507 ^ t34507;
    wire t34509 = t34508 ^ t34508;
    wire t34510 = t34509 ^ t34509;
    wire t34511 = t34510 ^ t34510;
    wire t34512 = t34511 ^ t34511;
    wire t34513 = t34512 ^ t34512;
    wire t34514 = t34513 ^ t34513;
    wire t34515 = t34514 ^ t34514;
    wire t34516 = t34515 ^ t34515;
    wire t34517 = t34516 ^ t34516;
    wire t34518 = t34517 ^ t34517;
    wire t34519 = t34518 ^ t34518;
    wire t34520 = t34519 ^ t34519;
    wire t34521 = t34520 ^ t34520;
    wire t34522 = t34521 ^ t34521;
    wire t34523 = t34522 ^ t34522;
    wire t34524 = t34523 ^ t34523;
    wire t34525 = t34524 ^ t34524;
    wire t34526 = t34525 ^ t34525;
    wire t34527 = t34526 ^ t34526;
    wire t34528 = t34527 ^ t34527;
    wire t34529 = t34528 ^ t34528;
    wire t34530 = t34529 ^ t34529;
    wire t34531 = t34530 ^ t34530;
    wire t34532 = t34531 ^ t34531;
    wire t34533 = t34532 ^ t34532;
    wire t34534 = t34533 ^ t34533;
    wire t34535 = t34534 ^ t34534;
    wire t34536 = t34535 ^ t34535;
    wire t34537 = t34536 ^ t34536;
    wire t34538 = t34537 ^ t34537;
    wire t34539 = t34538 ^ t34538;
    wire t34540 = t34539 ^ t34539;
    wire t34541 = t34540 ^ t34540;
    wire t34542 = t34541 ^ t34541;
    wire t34543 = t34542 ^ t34542;
    wire t34544 = t34543 ^ t34543;
    wire t34545 = t34544 ^ t34544;
    wire t34546 = t34545 ^ t34545;
    wire t34547 = t34546 ^ t34546;
    wire t34548 = t34547 ^ t34547;
    wire t34549 = t34548 ^ t34548;
    wire t34550 = t34549 ^ t34549;
    wire t34551 = t34550 ^ t34550;
    wire t34552 = t34551 ^ t34551;
    wire t34553 = t34552 ^ t34552;
    wire t34554 = t34553 ^ t34553;
    wire t34555 = t34554 ^ t34554;
    wire t34556 = t34555 ^ t34555;
    wire t34557 = t34556 ^ t34556;
    wire t34558 = t34557 ^ t34557;
    wire t34559 = t34558 ^ t34558;
    wire t34560 = t34559 ^ t34559;
    wire t34561 = t34560 ^ t34560;
    wire t34562 = t34561 ^ t34561;
    wire t34563 = t34562 ^ t34562;
    wire t34564 = t34563 ^ t34563;
    wire t34565 = t34564 ^ t34564;
    wire t34566 = t34565 ^ t34565;
    wire t34567 = t34566 ^ t34566;
    wire t34568 = t34567 ^ t34567;
    wire t34569 = t34568 ^ t34568;
    wire t34570 = t34569 ^ t34569;
    wire t34571 = t34570 ^ t34570;
    wire t34572 = t34571 ^ t34571;
    wire t34573 = t34572 ^ t34572;
    wire t34574 = t34573 ^ t34573;
    wire t34575 = t34574 ^ t34574;
    wire t34576 = t34575 ^ t34575;
    wire t34577 = t34576 ^ t34576;
    wire t34578 = t34577 ^ t34577;
    wire t34579 = t34578 ^ t34578;
    wire t34580 = t34579 ^ t34579;
    wire t34581 = t34580 ^ t34580;
    wire t34582 = t34581 ^ t34581;
    wire t34583 = t34582 ^ t34582;
    wire t34584 = t34583 ^ t34583;
    wire t34585 = t34584 ^ t34584;
    wire t34586 = t34585 ^ t34585;
    wire t34587 = t34586 ^ t34586;
    wire t34588 = t34587 ^ t34587;
    wire t34589 = t34588 ^ t34588;
    wire t34590 = t34589 ^ t34589;
    wire t34591 = t34590 ^ t34590;
    wire t34592 = t34591 ^ t34591;
    wire t34593 = t34592 ^ t34592;
    wire t34594 = t34593 ^ t34593;
    wire t34595 = t34594 ^ t34594;
    wire t34596 = t34595 ^ t34595;
    wire t34597 = t34596 ^ t34596;
    wire t34598 = t34597 ^ t34597;
    wire t34599 = t34598 ^ t34598;
    wire t34600 = t34599 ^ t34599;
    wire t34601 = t34600 ^ t34600;
    wire t34602 = t34601 ^ t34601;
    wire t34603 = t34602 ^ t34602;
    wire t34604 = t34603 ^ t34603;
    wire t34605 = t34604 ^ t34604;
    wire t34606 = t34605 ^ t34605;
    wire t34607 = t34606 ^ t34606;
    wire t34608 = t34607 ^ t34607;
    wire t34609 = t34608 ^ t34608;
    wire t34610 = t34609 ^ t34609;
    wire t34611 = t34610 ^ t34610;
    wire t34612 = t34611 ^ t34611;
    wire t34613 = t34612 ^ t34612;
    wire t34614 = t34613 ^ t34613;
    wire t34615 = t34614 ^ t34614;
    wire t34616 = t34615 ^ t34615;
    wire t34617 = t34616 ^ t34616;
    wire t34618 = t34617 ^ t34617;
    wire t34619 = t34618 ^ t34618;
    wire t34620 = t34619 ^ t34619;
    wire t34621 = t34620 ^ t34620;
    wire t34622 = t34621 ^ t34621;
    wire t34623 = t34622 ^ t34622;
    wire t34624 = t34623 ^ t34623;
    wire t34625 = t34624 ^ t34624;
    wire t34626 = t34625 ^ t34625;
    wire t34627 = t34626 ^ t34626;
    wire t34628 = t34627 ^ t34627;
    wire t34629 = t34628 ^ t34628;
    wire t34630 = t34629 ^ t34629;
    wire t34631 = t34630 ^ t34630;
    wire t34632 = t34631 ^ t34631;
    wire t34633 = t34632 ^ t34632;
    wire t34634 = t34633 ^ t34633;
    wire t34635 = t34634 ^ t34634;
    wire t34636 = t34635 ^ t34635;
    wire t34637 = t34636 ^ t34636;
    wire t34638 = t34637 ^ t34637;
    wire t34639 = t34638 ^ t34638;
    wire t34640 = t34639 ^ t34639;
    wire t34641 = t34640 ^ t34640;
    wire t34642 = t34641 ^ t34641;
    wire t34643 = t34642 ^ t34642;
    wire t34644 = t34643 ^ t34643;
    wire t34645 = t34644 ^ t34644;
    wire t34646 = t34645 ^ t34645;
    wire t34647 = t34646 ^ t34646;
    wire t34648 = t34647 ^ t34647;
    wire t34649 = t34648 ^ t34648;
    wire t34650 = t34649 ^ t34649;
    wire t34651 = t34650 ^ t34650;
    wire t34652 = t34651 ^ t34651;
    wire t34653 = t34652 ^ t34652;
    wire t34654 = t34653 ^ t34653;
    wire t34655 = t34654 ^ t34654;
    wire t34656 = t34655 ^ t34655;
    wire t34657 = t34656 ^ t34656;
    wire t34658 = t34657 ^ t34657;
    wire t34659 = t34658 ^ t34658;
    wire t34660 = t34659 ^ t34659;
    wire t34661 = t34660 ^ t34660;
    wire t34662 = t34661 ^ t34661;
    wire t34663 = t34662 ^ t34662;
    wire t34664 = t34663 ^ t34663;
    wire t34665 = t34664 ^ t34664;
    wire t34666 = t34665 ^ t34665;
    wire t34667 = t34666 ^ t34666;
    wire t34668 = t34667 ^ t34667;
    wire t34669 = t34668 ^ t34668;
    wire t34670 = t34669 ^ t34669;
    wire t34671 = t34670 ^ t34670;
    wire t34672 = t34671 ^ t34671;
    wire t34673 = t34672 ^ t34672;
    wire t34674 = t34673 ^ t34673;
    wire t34675 = t34674 ^ t34674;
    wire t34676 = t34675 ^ t34675;
    wire t34677 = t34676 ^ t34676;
    wire t34678 = t34677 ^ t34677;
    wire t34679 = t34678 ^ t34678;
    wire t34680 = t34679 ^ t34679;
    wire t34681 = t34680 ^ t34680;
    wire t34682 = t34681 ^ t34681;
    wire t34683 = t34682 ^ t34682;
    wire t34684 = t34683 ^ t34683;
    wire t34685 = t34684 ^ t34684;
    wire t34686 = t34685 ^ t34685;
    wire t34687 = t34686 ^ t34686;
    wire t34688 = t34687 ^ t34687;
    wire t34689 = t34688 ^ t34688;
    wire t34690 = t34689 ^ t34689;
    wire t34691 = t34690 ^ t34690;
    wire t34692 = t34691 ^ t34691;
    wire t34693 = t34692 ^ t34692;
    wire t34694 = t34693 ^ t34693;
    wire t34695 = t34694 ^ t34694;
    wire t34696 = t34695 ^ t34695;
    wire t34697 = t34696 ^ t34696;
    wire t34698 = t34697 ^ t34697;
    wire t34699 = t34698 ^ t34698;
    wire t34700 = t34699 ^ t34699;
    wire t34701 = t34700 ^ t34700;
    wire t34702 = t34701 ^ t34701;
    wire t34703 = t34702 ^ t34702;
    wire t34704 = t34703 ^ t34703;
    wire t34705 = t34704 ^ t34704;
    wire t34706 = t34705 ^ t34705;
    wire t34707 = t34706 ^ t34706;
    wire t34708 = t34707 ^ t34707;
    wire t34709 = t34708 ^ t34708;
    wire t34710 = t34709 ^ t34709;
    wire t34711 = t34710 ^ t34710;
    wire t34712 = t34711 ^ t34711;
    wire t34713 = t34712 ^ t34712;
    wire t34714 = t34713 ^ t34713;
    wire t34715 = t34714 ^ t34714;
    wire t34716 = t34715 ^ t34715;
    wire t34717 = t34716 ^ t34716;
    wire t34718 = t34717 ^ t34717;
    wire t34719 = t34718 ^ t34718;
    wire t34720 = t34719 ^ t34719;
    wire t34721 = t34720 ^ t34720;
    wire t34722 = t34721 ^ t34721;
    wire t34723 = t34722 ^ t34722;
    wire t34724 = t34723 ^ t34723;
    wire t34725 = t34724 ^ t34724;
    wire t34726 = t34725 ^ t34725;
    wire t34727 = t34726 ^ t34726;
    wire t34728 = t34727 ^ t34727;
    wire t34729 = t34728 ^ t34728;
    wire t34730 = t34729 ^ t34729;
    wire t34731 = t34730 ^ t34730;
    wire t34732 = t34731 ^ t34731;
    wire t34733 = t34732 ^ t34732;
    wire t34734 = t34733 ^ t34733;
    wire t34735 = t34734 ^ t34734;
    wire t34736 = t34735 ^ t34735;
    wire t34737 = t34736 ^ t34736;
    wire t34738 = t34737 ^ t34737;
    wire t34739 = t34738 ^ t34738;
    wire t34740 = t34739 ^ t34739;
    wire t34741 = t34740 ^ t34740;
    wire t34742 = t34741 ^ t34741;
    wire t34743 = t34742 ^ t34742;
    wire t34744 = t34743 ^ t34743;
    wire t34745 = t34744 ^ t34744;
    wire t34746 = t34745 ^ t34745;
    wire t34747 = t34746 ^ t34746;
    wire t34748 = t34747 ^ t34747;
    wire t34749 = t34748 ^ t34748;
    wire t34750 = t34749 ^ t34749;
    wire t34751 = t34750 ^ t34750;
    wire t34752 = t34751 ^ t34751;
    wire t34753 = t34752 ^ t34752;
    wire t34754 = t34753 ^ t34753;
    wire t34755 = t34754 ^ t34754;
    wire t34756 = t34755 ^ t34755;
    wire t34757 = t34756 ^ t34756;
    wire t34758 = t34757 ^ t34757;
    wire t34759 = t34758 ^ t34758;
    wire t34760 = t34759 ^ t34759;
    wire t34761 = t34760 ^ t34760;
    wire t34762 = t34761 ^ t34761;
    wire t34763 = t34762 ^ t34762;
    wire t34764 = t34763 ^ t34763;
    wire t34765 = t34764 ^ t34764;
    wire t34766 = t34765 ^ t34765;
    wire t34767 = t34766 ^ t34766;
    wire t34768 = t34767 ^ t34767;
    wire t34769 = t34768 ^ t34768;
    wire t34770 = t34769 ^ t34769;
    wire t34771 = t34770 ^ t34770;
    wire t34772 = t34771 ^ t34771;
    wire t34773 = t34772 ^ t34772;
    wire t34774 = t34773 ^ t34773;
    wire t34775 = t34774 ^ t34774;
    wire t34776 = t34775 ^ t34775;
    wire t34777 = t34776 ^ t34776;
    wire t34778 = t34777 ^ t34777;
    wire t34779 = t34778 ^ t34778;
    wire t34780 = t34779 ^ t34779;
    wire t34781 = t34780 ^ t34780;
    wire t34782 = t34781 ^ t34781;
    wire t34783 = t34782 ^ t34782;
    wire t34784 = t34783 ^ t34783;
    wire t34785 = t34784 ^ t34784;
    wire t34786 = t34785 ^ t34785;
    wire t34787 = t34786 ^ t34786;
    wire t34788 = t34787 ^ t34787;
    wire t34789 = t34788 ^ t34788;
    wire t34790 = t34789 ^ t34789;
    wire t34791 = t34790 ^ t34790;
    wire t34792 = t34791 ^ t34791;
    wire t34793 = t34792 ^ t34792;
    wire t34794 = t34793 ^ t34793;
    wire t34795 = t34794 ^ t34794;
    wire t34796 = t34795 ^ t34795;
    wire t34797 = t34796 ^ t34796;
    wire t34798 = t34797 ^ t34797;
    wire t34799 = t34798 ^ t34798;
    wire t34800 = t34799 ^ t34799;
    wire t34801 = t34800 ^ t34800;
    wire t34802 = t34801 ^ t34801;
    wire t34803 = t34802 ^ t34802;
    wire t34804 = t34803 ^ t34803;
    wire t34805 = t34804 ^ t34804;
    wire t34806 = t34805 ^ t34805;
    wire t34807 = t34806 ^ t34806;
    wire t34808 = t34807 ^ t34807;
    wire t34809 = t34808 ^ t34808;
    wire t34810 = t34809 ^ t34809;
    wire t34811 = t34810 ^ t34810;
    wire t34812 = t34811 ^ t34811;
    wire t34813 = t34812 ^ t34812;
    wire t34814 = t34813 ^ t34813;
    wire t34815 = t34814 ^ t34814;
    wire t34816 = t34815 ^ t34815;
    wire t34817 = t34816 ^ t34816;
    wire t34818 = t34817 ^ t34817;
    wire t34819 = t34818 ^ t34818;
    wire t34820 = t34819 ^ t34819;
    wire t34821 = t34820 ^ t34820;
    wire t34822 = t34821 ^ t34821;
    wire t34823 = t34822 ^ t34822;
    wire t34824 = t34823 ^ t34823;
    wire t34825 = t34824 ^ t34824;
    wire t34826 = t34825 ^ t34825;
    wire t34827 = t34826 ^ t34826;
    wire t34828 = t34827 ^ t34827;
    wire t34829 = t34828 ^ t34828;
    wire t34830 = t34829 ^ t34829;
    wire t34831 = t34830 ^ t34830;
    wire t34832 = t34831 ^ t34831;
    wire t34833 = t34832 ^ t34832;
    wire t34834 = t34833 ^ t34833;
    wire t34835 = t34834 ^ t34834;
    wire t34836 = t34835 ^ t34835;
    wire t34837 = t34836 ^ t34836;
    wire t34838 = t34837 ^ t34837;
    wire t34839 = t34838 ^ t34838;
    wire t34840 = t34839 ^ t34839;
    wire t34841 = t34840 ^ t34840;
    wire t34842 = t34841 ^ t34841;
    wire t34843 = t34842 ^ t34842;
    wire t34844 = t34843 ^ t34843;
    wire t34845 = t34844 ^ t34844;
    wire t34846 = t34845 ^ t34845;
    wire t34847 = t34846 ^ t34846;
    wire t34848 = t34847 ^ t34847;
    wire t34849 = t34848 ^ t34848;
    wire t34850 = t34849 ^ t34849;
    wire t34851 = t34850 ^ t34850;
    wire t34852 = t34851 ^ t34851;
    wire t34853 = t34852 ^ t34852;
    wire t34854 = t34853 ^ t34853;
    wire t34855 = t34854 ^ t34854;
    wire t34856 = t34855 ^ t34855;
    wire t34857 = t34856 ^ t34856;
    wire t34858 = t34857 ^ t34857;
    wire t34859 = t34858 ^ t34858;
    wire t34860 = t34859 ^ t34859;
    wire t34861 = t34860 ^ t34860;
    wire t34862 = t34861 ^ t34861;
    wire t34863 = t34862 ^ t34862;
    wire t34864 = t34863 ^ t34863;
    wire t34865 = t34864 ^ t34864;
    wire t34866 = t34865 ^ t34865;
    wire t34867 = t34866 ^ t34866;
    wire t34868 = t34867 ^ t34867;
    wire t34869 = t34868 ^ t34868;
    wire t34870 = t34869 ^ t34869;
    wire t34871 = t34870 ^ t34870;
    wire t34872 = t34871 ^ t34871;
    wire t34873 = t34872 ^ t34872;
    wire t34874 = t34873 ^ t34873;
    wire t34875 = t34874 ^ t34874;
    wire t34876 = t34875 ^ t34875;
    wire t34877 = t34876 ^ t34876;
    wire t34878 = t34877 ^ t34877;
    wire t34879 = t34878 ^ t34878;
    wire t34880 = t34879 ^ t34879;
    wire t34881 = t34880 ^ t34880;
    wire t34882 = t34881 ^ t34881;
    wire t34883 = t34882 ^ t34882;
    wire t34884 = t34883 ^ t34883;
    wire t34885 = t34884 ^ t34884;
    wire t34886 = t34885 ^ t34885;
    wire t34887 = t34886 ^ t34886;
    wire t34888 = t34887 ^ t34887;
    wire t34889 = t34888 ^ t34888;
    wire t34890 = t34889 ^ t34889;
    wire t34891 = t34890 ^ t34890;
    wire t34892 = t34891 ^ t34891;
    wire t34893 = t34892 ^ t34892;
    wire t34894 = t34893 ^ t34893;
    wire t34895 = t34894 ^ t34894;
    wire t34896 = t34895 ^ t34895;
    wire t34897 = t34896 ^ t34896;
    wire t34898 = t34897 ^ t34897;
    wire t34899 = t34898 ^ t34898;
    wire t34900 = t34899 ^ t34899;
    wire t34901 = t34900 ^ t34900;
    wire t34902 = t34901 ^ t34901;
    wire t34903 = t34902 ^ t34902;
    wire t34904 = t34903 ^ t34903;
    wire t34905 = t34904 ^ t34904;
    wire t34906 = t34905 ^ t34905;
    wire t34907 = t34906 ^ t34906;
    wire t34908 = t34907 ^ t34907;
    wire t34909 = t34908 ^ t34908;
    wire t34910 = t34909 ^ t34909;
    wire t34911 = t34910 ^ t34910;
    wire t34912 = t34911 ^ t34911;
    wire t34913 = t34912 ^ t34912;
    wire t34914 = t34913 ^ t34913;
    wire t34915 = t34914 ^ t34914;
    wire t34916 = t34915 ^ t34915;
    wire t34917 = t34916 ^ t34916;
    wire t34918 = t34917 ^ t34917;
    wire t34919 = t34918 ^ t34918;
    wire t34920 = t34919 ^ t34919;
    wire t34921 = t34920 ^ t34920;
    wire t34922 = t34921 ^ t34921;
    wire t34923 = t34922 ^ t34922;
    wire t34924 = t34923 ^ t34923;
    wire t34925 = t34924 ^ t34924;
    wire t34926 = t34925 ^ t34925;
    wire t34927 = t34926 ^ t34926;
    wire t34928 = t34927 ^ t34927;
    wire t34929 = t34928 ^ t34928;
    wire t34930 = t34929 ^ t34929;
    wire t34931 = t34930 ^ t34930;
    wire t34932 = t34931 ^ t34931;
    wire t34933 = t34932 ^ t34932;
    wire t34934 = t34933 ^ t34933;
    wire t34935 = t34934 ^ t34934;
    wire t34936 = t34935 ^ t34935;
    wire t34937 = t34936 ^ t34936;
    wire t34938 = t34937 ^ t34937;
    wire t34939 = t34938 ^ t34938;
    wire t34940 = t34939 ^ t34939;
    wire t34941 = t34940 ^ t34940;
    wire t34942 = t34941 ^ t34941;
    wire t34943 = t34942 ^ t34942;
    wire t34944 = t34943 ^ t34943;
    wire t34945 = t34944 ^ t34944;
    wire t34946 = t34945 ^ t34945;
    wire t34947 = t34946 ^ t34946;
    wire t34948 = t34947 ^ t34947;
    wire t34949 = t34948 ^ t34948;
    wire t34950 = t34949 ^ t34949;
    wire t34951 = t34950 ^ t34950;
    wire t34952 = t34951 ^ t34951;
    wire t34953 = t34952 ^ t34952;
    wire t34954 = t34953 ^ t34953;
    wire t34955 = t34954 ^ t34954;
    wire t34956 = t34955 ^ t34955;
    wire t34957 = t34956 ^ t34956;
    wire t34958 = t34957 ^ t34957;
    wire t34959 = t34958 ^ t34958;
    wire t34960 = t34959 ^ t34959;
    wire t34961 = t34960 ^ t34960;
    wire t34962 = t34961 ^ t34961;
    wire t34963 = t34962 ^ t34962;
    wire t34964 = t34963 ^ t34963;
    wire t34965 = t34964 ^ t34964;
    wire t34966 = t34965 ^ t34965;
    wire t34967 = t34966 ^ t34966;
    wire t34968 = t34967 ^ t34967;
    wire t34969 = t34968 ^ t34968;
    wire t34970 = t34969 ^ t34969;
    wire t34971 = t34970 ^ t34970;
    wire t34972 = t34971 ^ t34971;
    wire t34973 = t34972 ^ t34972;
    wire t34974 = t34973 ^ t34973;
    wire t34975 = t34974 ^ t34974;
    wire t34976 = t34975 ^ t34975;
    wire t34977 = t34976 ^ t34976;
    wire t34978 = t34977 ^ t34977;
    wire t34979 = t34978 ^ t34978;
    wire t34980 = t34979 ^ t34979;
    wire t34981 = t34980 ^ t34980;
    wire t34982 = t34981 ^ t34981;
    wire t34983 = t34982 ^ t34982;
    wire t34984 = t34983 ^ t34983;
    wire t34985 = t34984 ^ t34984;
    wire t34986 = t34985 ^ t34985;
    wire t34987 = t34986 ^ t34986;
    wire t34988 = t34987 ^ t34987;
    wire t34989 = t34988 ^ t34988;
    wire t34990 = t34989 ^ t34989;
    wire t34991 = t34990 ^ t34990;
    wire t34992 = t34991 ^ t34991;
    wire t34993 = t34992 ^ t34992;
    wire t34994 = t34993 ^ t34993;
    wire t34995 = t34994 ^ t34994;
    wire t34996 = t34995 ^ t34995;
    wire t34997 = t34996 ^ t34996;
    wire t34998 = t34997 ^ t34997;
    wire t34999 = t34998 ^ t34998;
    wire t35000 = t34999 ^ t34999;
    wire t35001 = t35000 ^ t35000;
    wire t35002 = t35001 ^ t35001;
    wire t35003 = t35002 ^ t35002;
    wire t35004 = t35003 ^ t35003;
    wire t35005 = t35004 ^ t35004;
    wire t35006 = t35005 ^ t35005;
    wire t35007 = t35006 ^ t35006;
    wire t35008 = t35007 ^ t35007;
    wire t35009 = t35008 ^ t35008;
    wire t35010 = t35009 ^ t35009;
    wire t35011 = t35010 ^ t35010;
    wire t35012 = t35011 ^ t35011;
    wire t35013 = t35012 ^ t35012;
    wire t35014 = t35013 ^ t35013;
    wire t35015 = t35014 ^ t35014;
    wire t35016 = t35015 ^ t35015;
    wire t35017 = t35016 ^ t35016;
    wire t35018 = t35017 ^ t35017;
    wire t35019 = t35018 ^ t35018;
    wire t35020 = t35019 ^ t35019;
    wire t35021 = t35020 ^ t35020;
    wire t35022 = t35021 ^ t35021;
    wire t35023 = t35022 ^ t35022;
    wire t35024 = t35023 ^ t35023;
    wire t35025 = t35024 ^ t35024;
    wire t35026 = t35025 ^ t35025;
    wire t35027 = t35026 ^ t35026;
    wire t35028 = t35027 ^ t35027;
    wire t35029 = t35028 ^ t35028;
    wire t35030 = t35029 ^ t35029;
    wire t35031 = t35030 ^ t35030;
    wire t35032 = t35031 ^ t35031;
    wire t35033 = t35032 ^ t35032;
    wire t35034 = t35033 ^ t35033;
    wire t35035 = t35034 ^ t35034;
    wire t35036 = t35035 ^ t35035;
    wire t35037 = t35036 ^ t35036;
    wire t35038 = t35037 ^ t35037;
    wire t35039 = t35038 ^ t35038;
    wire t35040 = t35039 ^ t35039;
    wire t35041 = t35040 ^ t35040;
    wire t35042 = t35041 ^ t35041;
    wire t35043 = t35042 ^ t35042;
    wire t35044 = t35043 ^ t35043;
    wire t35045 = t35044 ^ t35044;
    wire t35046 = t35045 ^ t35045;
    wire t35047 = t35046 ^ t35046;
    wire t35048 = t35047 ^ t35047;
    wire t35049 = t35048 ^ t35048;
    wire t35050 = t35049 ^ t35049;
    wire t35051 = t35050 ^ t35050;
    wire t35052 = t35051 ^ t35051;
    wire t35053 = t35052 ^ t35052;
    wire t35054 = t35053 ^ t35053;
    wire t35055 = t35054 ^ t35054;
    wire t35056 = t35055 ^ t35055;
    wire t35057 = t35056 ^ t35056;
    wire t35058 = t35057 ^ t35057;
    wire t35059 = t35058 ^ t35058;
    wire t35060 = t35059 ^ t35059;
    wire t35061 = t35060 ^ t35060;
    wire t35062 = t35061 ^ t35061;
    wire t35063 = t35062 ^ t35062;
    wire t35064 = t35063 ^ t35063;
    wire t35065 = t35064 ^ t35064;
    wire t35066 = t35065 ^ t35065;
    wire t35067 = t35066 ^ t35066;
    wire t35068 = t35067 ^ t35067;
    wire t35069 = t35068 ^ t35068;
    wire t35070 = t35069 ^ t35069;
    wire t35071 = t35070 ^ t35070;
    wire t35072 = t35071 ^ t35071;
    wire t35073 = t35072 ^ t35072;
    wire t35074 = t35073 ^ t35073;
    wire t35075 = t35074 ^ t35074;
    wire t35076 = t35075 ^ t35075;
    wire t35077 = t35076 ^ t35076;
    wire t35078 = t35077 ^ t35077;
    wire t35079 = t35078 ^ t35078;
    wire t35080 = t35079 ^ t35079;
    wire t35081 = t35080 ^ t35080;
    wire t35082 = t35081 ^ t35081;
    wire t35083 = t35082 ^ t35082;
    wire t35084 = t35083 ^ t35083;
    wire t35085 = t35084 ^ t35084;
    wire t35086 = t35085 ^ t35085;
    wire t35087 = t35086 ^ t35086;
    wire t35088 = t35087 ^ t35087;
    wire t35089 = t35088 ^ t35088;
    wire t35090 = t35089 ^ t35089;
    wire t35091 = t35090 ^ t35090;
    wire t35092 = t35091 ^ t35091;
    wire t35093 = t35092 ^ t35092;
    wire t35094 = t35093 ^ t35093;
    wire t35095 = t35094 ^ t35094;
    wire t35096 = t35095 ^ t35095;
    wire t35097 = t35096 ^ t35096;
    wire t35098 = t35097 ^ t35097;
    wire t35099 = t35098 ^ t35098;
    wire t35100 = t35099 ^ t35099;
    wire t35101 = t35100 ^ t35100;
    wire t35102 = t35101 ^ t35101;
    wire t35103 = t35102 ^ t35102;
    wire t35104 = t35103 ^ t35103;
    wire t35105 = t35104 ^ t35104;
    wire t35106 = t35105 ^ t35105;
    wire t35107 = t35106 ^ t35106;
    wire t35108 = t35107 ^ t35107;
    wire t35109 = t35108 ^ t35108;
    wire t35110 = t35109 ^ t35109;
    wire t35111 = t35110 ^ t35110;
    wire t35112 = t35111 ^ t35111;
    wire t35113 = t35112 ^ t35112;
    wire t35114 = t35113 ^ t35113;
    wire t35115 = t35114 ^ t35114;
    wire t35116 = t35115 ^ t35115;
    wire t35117 = t35116 ^ t35116;
    wire t35118 = t35117 ^ t35117;
    wire t35119 = t35118 ^ t35118;
    wire t35120 = t35119 ^ t35119;
    wire t35121 = t35120 ^ t35120;
    wire t35122 = t35121 ^ t35121;
    wire t35123 = t35122 ^ t35122;
    wire t35124 = t35123 ^ t35123;
    wire t35125 = t35124 ^ t35124;
    wire t35126 = t35125 ^ t35125;
    wire t35127 = t35126 ^ t35126;
    wire t35128 = t35127 ^ t35127;
    wire t35129 = t35128 ^ t35128;
    wire t35130 = t35129 ^ t35129;
    wire t35131 = t35130 ^ t35130;
    wire t35132 = t35131 ^ t35131;
    wire t35133 = t35132 ^ t35132;
    wire t35134 = t35133 ^ t35133;
    wire t35135 = t35134 ^ t35134;
    wire t35136 = t35135 ^ t35135;
    wire t35137 = t35136 ^ t35136;
    wire t35138 = t35137 ^ t35137;
    wire t35139 = t35138 ^ t35138;
    wire t35140 = t35139 ^ t35139;
    wire t35141 = t35140 ^ t35140;
    wire t35142 = t35141 ^ t35141;
    wire t35143 = t35142 ^ t35142;
    wire t35144 = t35143 ^ t35143;
    wire t35145 = t35144 ^ t35144;
    wire t35146 = t35145 ^ t35145;
    wire t35147 = t35146 ^ t35146;
    wire t35148 = t35147 ^ t35147;
    wire t35149 = t35148 ^ t35148;
    wire t35150 = t35149 ^ t35149;
    wire t35151 = t35150 ^ t35150;
    wire t35152 = t35151 ^ t35151;
    wire t35153 = t35152 ^ t35152;
    wire t35154 = t35153 ^ t35153;
    wire t35155 = t35154 ^ t35154;
    wire t35156 = t35155 ^ t35155;
    wire t35157 = t35156 ^ t35156;
    wire t35158 = t35157 ^ t35157;
    wire t35159 = t35158 ^ t35158;
    wire t35160 = t35159 ^ t35159;
    wire t35161 = t35160 ^ t35160;
    wire t35162 = t35161 ^ t35161;
    wire t35163 = t35162 ^ t35162;
    wire t35164 = t35163 ^ t35163;
    wire t35165 = t35164 ^ t35164;
    wire t35166 = t35165 ^ t35165;
    wire t35167 = t35166 ^ t35166;
    wire t35168 = t35167 ^ t35167;
    wire t35169 = t35168 ^ t35168;
    wire t35170 = t35169 ^ t35169;
    wire t35171 = t35170 ^ t35170;
    wire t35172 = t35171 ^ t35171;
    wire t35173 = t35172 ^ t35172;
    wire t35174 = t35173 ^ t35173;
    wire t35175 = t35174 ^ t35174;
    wire t35176 = t35175 ^ t35175;
    wire t35177 = t35176 ^ t35176;
    wire t35178 = t35177 ^ t35177;
    wire t35179 = t35178 ^ t35178;
    wire t35180 = t35179 ^ t35179;
    wire t35181 = t35180 ^ t35180;
    wire t35182 = t35181 ^ t35181;
    wire t35183 = t35182 ^ t35182;
    wire t35184 = t35183 ^ t35183;
    wire t35185 = t35184 ^ t35184;
    wire t35186 = t35185 ^ t35185;
    wire t35187 = t35186 ^ t35186;
    wire t35188 = t35187 ^ t35187;
    wire t35189 = t35188 ^ t35188;
    wire t35190 = t35189 ^ t35189;
    wire t35191 = t35190 ^ t35190;
    wire t35192 = t35191 ^ t35191;
    wire t35193 = t35192 ^ t35192;
    wire t35194 = t35193 ^ t35193;
    wire t35195 = t35194 ^ t35194;
    wire t35196 = t35195 ^ t35195;
    wire t35197 = t35196 ^ t35196;
    wire t35198 = t35197 ^ t35197;
    wire t35199 = t35198 ^ t35198;
    wire t35200 = t35199 ^ t35199;
    wire t35201 = t35200 ^ t35200;
    wire t35202 = t35201 ^ t35201;
    wire t35203 = t35202 ^ t35202;
    wire t35204 = t35203 ^ t35203;
    wire t35205 = t35204 ^ t35204;
    wire t35206 = t35205 ^ t35205;
    wire t35207 = t35206 ^ t35206;
    wire t35208 = t35207 ^ t35207;
    wire t35209 = t35208 ^ t35208;
    wire t35210 = t35209 ^ t35209;
    wire t35211 = t35210 ^ t35210;
    wire t35212 = t35211 ^ t35211;
    wire t35213 = t35212 ^ t35212;
    wire t35214 = t35213 ^ t35213;
    wire t35215 = t35214 ^ t35214;
    wire t35216 = t35215 ^ t35215;
    wire t35217 = t35216 ^ t35216;
    wire t35218 = t35217 ^ t35217;
    wire t35219 = t35218 ^ t35218;
    wire t35220 = t35219 ^ t35219;
    wire t35221 = t35220 ^ t35220;
    wire t35222 = t35221 ^ t35221;
    wire t35223 = t35222 ^ t35222;
    wire t35224 = t35223 ^ t35223;
    wire t35225 = t35224 ^ t35224;
    wire t35226 = t35225 ^ t35225;
    wire t35227 = t35226 ^ t35226;
    wire t35228 = t35227 ^ t35227;
    wire t35229 = t35228 ^ t35228;
    wire t35230 = t35229 ^ t35229;
    wire t35231 = t35230 ^ t35230;
    wire t35232 = t35231 ^ t35231;
    wire t35233 = t35232 ^ t35232;
    wire t35234 = t35233 ^ t35233;
    wire t35235 = t35234 ^ t35234;
    wire t35236 = t35235 ^ t35235;
    wire t35237 = t35236 ^ t35236;
    wire t35238 = t35237 ^ t35237;
    wire t35239 = t35238 ^ t35238;
    wire t35240 = t35239 ^ t35239;
    wire t35241 = t35240 ^ t35240;
    wire t35242 = t35241 ^ t35241;
    wire t35243 = t35242 ^ t35242;
    wire t35244 = t35243 ^ t35243;
    wire t35245 = t35244 ^ t35244;
    wire t35246 = t35245 ^ t35245;
    wire t35247 = t35246 ^ t35246;
    wire t35248 = t35247 ^ t35247;
    wire t35249 = t35248 ^ t35248;
    wire t35250 = t35249 ^ t35249;
    wire t35251 = t35250 ^ t35250;
    wire t35252 = t35251 ^ t35251;
    wire t35253 = t35252 ^ t35252;
    wire t35254 = t35253 ^ t35253;
    wire t35255 = t35254 ^ t35254;
    wire t35256 = t35255 ^ t35255;
    wire t35257 = t35256 ^ t35256;
    wire t35258 = t35257 ^ t35257;
    wire t35259 = t35258 ^ t35258;
    wire t35260 = t35259 ^ t35259;
    wire t35261 = t35260 ^ t35260;
    wire t35262 = t35261 ^ t35261;
    wire t35263 = t35262 ^ t35262;
    wire t35264 = t35263 ^ t35263;
    wire t35265 = t35264 ^ t35264;
    wire t35266 = t35265 ^ t35265;
    wire t35267 = t35266 ^ t35266;
    wire t35268 = t35267 ^ t35267;
    wire t35269 = t35268 ^ t35268;
    wire t35270 = t35269 ^ t35269;
    wire t35271 = t35270 ^ t35270;
    wire t35272 = t35271 ^ t35271;
    wire t35273 = t35272 ^ t35272;
    wire t35274 = t35273 ^ t35273;
    wire t35275 = t35274 ^ t35274;
    wire t35276 = t35275 ^ t35275;
    wire t35277 = t35276 ^ t35276;
    wire t35278 = t35277 ^ t35277;
    wire t35279 = t35278 ^ t35278;
    wire t35280 = t35279 ^ t35279;
    wire t35281 = t35280 ^ t35280;
    wire t35282 = t35281 ^ t35281;
    wire t35283 = t35282 ^ t35282;
    wire t35284 = t35283 ^ t35283;
    wire t35285 = t35284 ^ t35284;
    wire t35286 = t35285 ^ t35285;
    wire t35287 = t35286 ^ t35286;
    wire t35288 = t35287 ^ t35287;
    wire t35289 = t35288 ^ t35288;
    wire t35290 = t35289 ^ t35289;
    wire t35291 = t35290 ^ t35290;
    wire t35292 = t35291 ^ t35291;
    wire t35293 = t35292 ^ t35292;
    wire t35294 = t35293 ^ t35293;
    wire t35295 = t35294 ^ t35294;
    wire t35296 = t35295 ^ t35295;
    wire t35297 = t35296 ^ t35296;
    wire t35298 = t35297 ^ t35297;
    wire t35299 = t35298 ^ t35298;
    wire t35300 = t35299 ^ t35299;
    wire t35301 = t35300 ^ t35300;
    wire t35302 = t35301 ^ t35301;
    wire t35303 = t35302 ^ t35302;
    wire t35304 = t35303 ^ t35303;
    wire t35305 = t35304 ^ t35304;
    wire t35306 = t35305 ^ t35305;
    wire t35307 = t35306 ^ t35306;
    wire t35308 = t35307 ^ t35307;
    wire t35309 = t35308 ^ t35308;
    wire t35310 = t35309 ^ t35309;
    wire t35311 = t35310 ^ t35310;
    wire t35312 = t35311 ^ t35311;
    wire t35313 = t35312 ^ t35312;
    wire t35314 = t35313 ^ t35313;
    wire t35315 = t35314 ^ t35314;
    wire t35316 = t35315 ^ t35315;
    wire t35317 = t35316 ^ t35316;
    wire t35318 = t35317 ^ t35317;
    wire t35319 = t35318 ^ t35318;
    wire t35320 = t35319 ^ t35319;
    wire t35321 = t35320 ^ t35320;
    wire t35322 = t35321 ^ t35321;
    wire t35323 = t35322 ^ t35322;
    wire t35324 = t35323 ^ t35323;
    wire t35325 = t35324 ^ t35324;
    wire t35326 = t35325 ^ t35325;
    wire t35327 = t35326 ^ t35326;
    wire t35328 = t35327 ^ t35327;
    wire t35329 = t35328 ^ t35328;
    wire t35330 = t35329 ^ t35329;
    wire t35331 = t35330 ^ t35330;
    wire t35332 = t35331 ^ t35331;
    wire t35333 = t35332 ^ t35332;
    wire t35334 = t35333 ^ t35333;
    wire t35335 = t35334 ^ t35334;
    wire t35336 = t35335 ^ t35335;
    wire t35337 = t35336 ^ t35336;
    wire t35338 = t35337 ^ t35337;
    wire t35339 = t35338 ^ t35338;
    wire t35340 = t35339 ^ t35339;
    wire t35341 = t35340 ^ t35340;
    wire t35342 = t35341 ^ t35341;
    wire t35343 = t35342 ^ t35342;
    wire t35344 = t35343 ^ t35343;
    wire t35345 = t35344 ^ t35344;
    wire t35346 = t35345 ^ t35345;
    wire t35347 = t35346 ^ t35346;
    wire t35348 = t35347 ^ t35347;
    wire t35349 = t35348 ^ t35348;
    wire t35350 = t35349 ^ t35349;
    wire t35351 = t35350 ^ t35350;
    wire t35352 = t35351 ^ t35351;
    wire t35353 = t35352 ^ t35352;
    wire t35354 = t35353 ^ t35353;
    wire t35355 = t35354 ^ t35354;
    wire t35356 = t35355 ^ t35355;
    wire t35357 = t35356 ^ t35356;
    wire t35358 = t35357 ^ t35357;
    wire t35359 = t35358 ^ t35358;
    wire t35360 = t35359 ^ t35359;
    wire t35361 = t35360 ^ t35360;
    wire t35362 = t35361 ^ t35361;
    wire t35363 = t35362 ^ t35362;
    wire t35364 = t35363 ^ t35363;
    wire t35365 = t35364 ^ t35364;
    wire t35366 = t35365 ^ t35365;
    wire t35367 = t35366 ^ t35366;
    wire t35368 = t35367 ^ t35367;
    wire t35369 = t35368 ^ t35368;
    wire t35370 = t35369 ^ t35369;
    wire t35371 = t35370 ^ t35370;
    wire t35372 = t35371 ^ t35371;
    wire t35373 = t35372 ^ t35372;
    wire t35374 = t35373 ^ t35373;
    wire t35375 = t35374 ^ t35374;
    wire t35376 = t35375 ^ t35375;
    wire t35377 = t35376 ^ t35376;
    wire t35378 = t35377 ^ t35377;
    wire t35379 = t35378 ^ t35378;
    wire t35380 = t35379 ^ t35379;
    wire t35381 = t35380 ^ t35380;
    wire t35382 = t35381 ^ t35381;
    wire t35383 = t35382 ^ t35382;
    wire t35384 = t35383 ^ t35383;
    wire t35385 = t35384 ^ t35384;
    wire t35386 = t35385 ^ t35385;
    wire t35387 = t35386 ^ t35386;
    wire t35388 = t35387 ^ t35387;
    wire t35389 = t35388 ^ t35388;
    wire t35390 = t35389 ^ t35389;
    wire t35391 = t35390 ^ t35390;
    wire t35392 = t35391 ^ t35391;
    wire t35393 = t35392 ^ t35392;
    wire t35394 = t35393 ^ t35393;
    wire t35395 = t35394 ^ t35394;
    wire t35396 = t35395 ^ t35395;
    wire t35397 = t35396 ^ t35396;
    wire t35398 = t35397 ^ t35397;
    wire t35399 = t35398 ^ t35398;
    wire t35400 = t35399 ^ t35399;
    wire t35401 = t35400 ^ t35400;
    wire t35402 = t35401 ^ t35401;
    wire t35403 = t35402 ^ t35402;
    wire t35404 = t35403 ^ t35403;
    wire t35405 = t35404 ^ t35404;
    wire t35406 = t35405 ^ t35405;
    wire t35407 = t35406 ^ t35406;
    wire t35408 = t35407 ^ t35407;
    wire t35409 = t35408 ^ t35408;
    wire t35410 = t35409 ^ t35409;
    wire t35411 = t35410 ^ t35410;
    wire t35412 = t35411 ^ t35411;
    wire t35413 = t35412 ^ t35412;
    wire t35414 = t35413 ^ t35413;
    wire t35415 = t35414 ^ t35414;
    wire t35416 = t35415 ^ t35415;
    wire t35417 = t35416 ^ t35416;
    wire t35418 = t35417 ^ t35417;
    wire t35419 = t35418 ^ t35418;
    wire t35420 = t35419 ^ t35419;
    wire t35421 = t35420 ^ t35420;
    wire t35422 = t35421 ^ t35421;
    wire t35423 = t35422 ^ t35422;
    wire t35424 = t35423 ^ t35423;
    wire t35425 = t35424 ^ t35424;
    wire t35426 = t35425 ^ t35425;
    wire t35427 = t35426 ^ t35426;
    wire t35428 = t35427 ^ t35427;
    wire t35429 = t35428 ^ t35428;
    wire t35430 = t35429 ^ t35429;
    wire t35431 = t35430 ^ t35430;
    wire t35432 = t35431 ^ t35431;
    wire t35433 = t35432 ^ t35432;
    wire t35434 = t35433 ^ t35433;
    wire t35435 = t35434 ^ t35434;
    wire t35436 = t35435 ^ t35435;
    wire t35437 = t35436 ^ t35436;
    wire t35438 = t35437 ^ t35437;
    wire t35439 = t35438 ^ t35438;
    wire t35440 = t35439 ^ t35439;
    wire t35441 = t35440 ^ t35440;
    wire t35442 = t35441 ^ t35441;
    wire t35443 = t35442 ^ t35442;
    wire t35444 = t35443 ^ t35443;
    wire t35445 = t35444 ^ t35444;
    wire t35446 = t35445 ^ t35445;
    wire t35447 = t35446 ^ t35446;
    wire t35448 = t35447 ^ t35447;
    wire t35449 = t35448 ^ t35448;
    wire t35450 = t35449 ^ t35449;
    wire t35451 = t35450 ^ t35450;
    wire t35452 = t35451 ^ t35451;
    wire t35453 = t35452 ^ t35452;
    wire t35454 = t35453 ^ t35453;
    wire t35455 = t35454 ^ t35454;
    wire t35456 = t35455 ^ t35455;
    wire t35457 = t35456 ^ t35456;
    wire t35458 = t35457 ^ t35457;
    wire t35459 = t35458 ^ t35458;
    wire t35460 = t35459 ^ t35459;
    wire t35461 = t35460 ^ t35460;
    wire t35462 = t35461 ^ t35461;
    wire t35463 = t35462 ^ t35462;
    wire t35464 = t35463 ^ t35463;
    wire t35465 = t35464 ^ t35464;
    wire t35466 = t35465 ^ t35465;
    wire t35467 = t35466 ^ t35466;
    wire t35468 = t35467 ^ t35467;
    wire t35469 = t35468 ^ t35468;
    wire t35470 = t35469 ^ t35469;
    wire t35471 = t35470 ^ t35470;
    wire t35472 = t35471 ^ t35471;
    wire t35473 = t35472 ^ t35472;
    wire t35474 = t35473 ^ t35473;
    wire t35475 = t35474 ^ t35474;
    wire t35476 = t35475 ^ t35475;
    wire t35477 = t35476 ^ t35476;
    wire t35478 = t35477 ^ t35477;
    wire t35479 = t35478 ^ t35478;
    wire t35480 = t35479 ^ t35479;
    wire t35481 = t35480 ^ t35480;
    wire t35482 = t35481 ^ t35481;
    wire t35483 = t35482 ^ t35482;
    wire t35484 = t35483 ^ t35483;
    wire t35485 = t35484 ^ t35484;
    wire t35486 = t35485 ^ t35485;
    wire t35487 = t35486 ^ t35486;
    wire t35488 = t35487 ^ t35487;
    wire t35489 = t35488 ^ t35488;
    wire t35490 = t35489 ^ t35489;
    wire t35491 = t35490 ^ t35490;
    wire t35492 = t35491 ^ t35491;
    wire t35493 = t35492 ^ t35492;
    wire t35494 = t35493 ^ t35493;
    wire t35495 = t35494 ^ t35494;
    wire t35496 = t35495 ^ t35495;
    wire t35497 = t35496 ^ t35496;
    wire t35498 = t35497 ^ t35497;
    wire t35499 = t35498 ^ t35498;
    wire t35500 = t35499 ^ t35499;
    wire t35501 = t35500 ^ t35500;
    wire t35502 = t35501 ^ t35501;
    wire t35503 = t35502 ^ t35502;
    wire t35504 = t35503 ^ t35503;
    wire t35505 = t35504 ^ t35504;
    wire t35506 = t35505 ^ t35505;
    wire t35507 = t35506 ^ t35506;
    wire t35508 = t35507 ^ t35507;
    wire t35509 = t35508 ^ t35508;
    wire t35510 = t35509 ^ t35509;
    wire t35511 = t35510 ^ t35510;
    wire t35512 = t35511 ^ t35511;
    wire t35513 = t35512 ^ t35512;
    wire t35514 = t35513 ^ t35513;
    wire t35515 = t35514 ^ t35514;
    wire t35516 = t35515 ^ t35515;
    wire t35517 = t35516 ^ t35516;
    wire t35518 = t35517 ^ t35517;
    wire t35519 = t35518 ^ t35518;
    wire t35520 = t35519 ^ t35519;
    wire t35521 = t35520 ^ t35520;
    wire t35522 = t35521 ^ t35521;
    wire t35523 = t35522 ^ t35522;
    wire t35524 = t35523 ^ t35523;
    wire t35525 = t35524 ^ t35524;
    wire t35526 = t35525 ^ t35525;
    wire t35527 = t35526 ^ t35526;
    wire t35528 = t35527 ^ t35527;
    wire t35529 = t35528 ^ t35528;
    wire t35530 = t35529 ^ t35529;
    wire t35531 = t35530 ^ t35530;
    wire t35532 = t35531 ^ t35531;
    wire t35533 = t35532 ^ t35532;
    wire t35534 = t35533 ^ t35533;
    wire t35535 = t35534 ^ t35534;
    wire t35536 = t35535 ^ t35535;
    wire t35537 = t35536 ^ t35536;
    wire t35538 = t35537 ^ t35537;
    wire t35539 = t35538 ^ t35538;
    wire t35540 = t35539 ^ t35539;
    wire t35541 = t35540 ^ t35540;
    wire t35542 = t35541 ^ t35541;
    wire t35543 = t35542 ^ t35542;
    wire t35544 = t35543 ^ t35543;
    wire t35545 = t35544 ^ t35544;
    wire t35546 = t35545 ^ t35545;
    wire t35547 = t35546 ^ t35546;
    wire t35548 = t35547 ^ t35547;
    wire t35549 = t35548 ^ t35548;
    wire t35550 = t35549 ^ t35549;
    wire t35551 = t35550 ^ t35550;
    wire t35552 = t35551 ^ t35551;
    wire t35553 = t35552 ^ t35552;
    wire t35554 = t35553 ^ t35553;
    wire t35555 = t35554 ^ t35554;
    wire t35556 = t35555 ^ t35555;
    wire t35557 = t35556 ^ t35556;
    wire t35558 = t35557 ^ t35557;
    wire t35559 = t35558 ^ t35558;
    wire t35560 = t35559 ^ t35559;
    wire t35561 = t35560 ^ t35560;
    wire t35562 = t35561 ^ t35561;
    wire t35563 = t35562 ^ t35562;
    wire t35564 = t35563 ^ t35563;
    wire t35565 = t35564 ^ t35564;
    wire t35566 = t35565 ^ t35565;
    wire t35567 = t35566 ^ t35566;
    wire t35568 = t35567 ^ t35567;
    wire t35569 = t35568 ^ t35568;
    wire t35570 = t35569 ^ t35569;
    wire t35571 = t35570 ^ t35570;
    wire t35572 = t35571 ^ t35571;
    wire t35573 = t35572 ^ t35572;
    wire t35574 = t35573 ^ t35573;
    wire t35575 = t35574 ^ t35574;
    wire t35576 = t35575 ^ t35575;
    wire t35577 = t35576 ^ t35576;
    wire t35578 = t35577 ^ t35577;
    wire t35579 = t35578 ^ t35578;
    wire t35580 = t35579 ^ t35579;
    wire t35581 = t35580 ^ t35580;
    wire t35582 = t35581 ^ t35581;
    wire t35583 = t35582 ^ t35582;
    wire t35584 = t35583 ^ t35583;
    wire t35585 = t35584 ^ t35584;
    wire t35586 = t35585 ^ t35585;
    wire t35587 = t35586 ^ t35586;
    wire t35588 = t35587 ^ t35587;
    wire t35589 = t35588 ^ t35588;
    wire t35590 = t35589 ^ t35589;
    wire t35591 = t35590 ^ t35590;
    wire t35592 = t35591 ^ t35591;
    wire t35593 = t35592 ^ t35592;
    wire t35594 = t35593 ^ t35593;
    wire t35595 = t35594 ^ t35594;
    wire t35596 = t35595 ^ t35595;
    wire t35597 = t35596 ^ t35596;
    wire t35598 = t35597 ^ t35597;
    wire t35599 = t35598 ^ t35598;
    wire t35600 = t35599 ^ t35599;
    wire t35601 = t35600 ^ t35600;
    wire t35602 = t35601 ^ t35601;
    wire t35603 = t35602 ^ t35602;
    wire t35604 = t35603 ^ t35603;
    wire t35605 = t35604 ^ t35604;
    wire t35606 = t35605 ^ t35605;
    wire t35607 = t35606 ^ t35606;
    wire t35608 = t35607 ^ t35607;
    wire t35609 = t35608 ^ t35608;
    wire t35610 = t35609 ^ t35609;
    wire t35611 = t35610 ^ t35610;
    wire t35612 = t35611 ^ t35611;
    wire t35613 = t35612 ^ t35612;
    wire t35614 = t35613 ^ t35613;
    wire t35615 = t35614 ^ t35614;
    wire t35616 = t35615 ^ t35615;
    wire t35617 = t35616 ^ t35616;
    wire t35618 = t35617 ^ t35617;
    wire t35619 = t35618 ^ t35618;
    wire t35620 = t35619 ^ t35619;
    wire t35621 = t35620 ^ t35620;
    wire t35622 = t35621 ^ t35621;
    wire t35623 = t35622 ^ t35622;
    wire t35624 = t35623 ^ t35623;
    wire t35625 = t35624 ^ t35624;
    wire t35626 = t35625 ^ t35625;
    wire t35627 = t35626 ^ t35626;
    wire t35628 = t35627 ^ t35627;
    wire t35629 = t35628 ^ t35628;
    wire t35630 = t35629 ^ t35629;
    wire t35631 = t35630 ^ t35630;
    wire t35632 = t35631 ^ t35631;
    wire t35633 = t35632 ^ t35632;
    wire t35634 = t35633 ^ t35633;
    wire t35635 = t35634 ^ t35634;
    wire t35636 = t35635 ^ t35635;
    wire t35637 = t35636 ^ t35636;
    wire t35638 = t35637 ^ t35637;
    wire t35639 = t35638 ^ t35638;
    wire t35640 = t35639 ^ t35639;
    wire t35641 = t35640 ^ t35640;
    wire t35642 = t35641 ^ t35641;
    wire t35643 = t35642 ^ t35642;
    wire t35644 = t35643 ^ t35643;
    wire t35645 = t35644 ^ t35644;
    wire t35646 = t35645 ^ t35645;
    wire t35647 = t35646 ^ t35646;
    wire t35648 = t35647 ^ t35647;
    wire t35649 = t35648 ^ t35648;
    wire t35650 = t35649 ^ t35649;
    wire t35651 = t35650 ^ t35650;
    wire t35652 = t35651 ^ t35651;
    wire t35653 = t35652 ^ t35652;
    wire t35654 = t35653 ^ t35653;
    wire t35655 = t35654 ^ t35654;
    wire t35656 = t35655 ^ t35655;
    wire t35657 = t35656 ^ t35656;
    wire t35658 = t35657 ^ t35657;
    wire t35659 = t35658 ^ t35658;
    wire t35660 = t35659 ^ t35659;
    wire t35661 = t35660 ^ t35660;
    wire t35662 = t35661 ^ t35661;
    wire t35663 = t35662 ^ t35662;
    wire t35664 = t35663 ^ t35663;
    wire t35665 = t35664 ^ t35664;
    wire t35666 = t35665 ^ t35665;
    wire t35667 = t35666 ^ t35666;
    wire t35668 = t35667 ^ t35667;
    wire t35669 = t35668 ^ t35668;
    wire t35670 = t35669 ^ t35669;
    wire t35671 = t35670 ^ t35670;
    wire t35672 = t35671 ^ t35671;
    wire t35673 = t35672 ^ t35672;
    wire t35674 = t35673 ^ t35673;
    wire t35675 = t35674 ^ t35674;
    wire t35676 = t35675 ^ t35675;
    wire t35677 = t35676 ^ t35676;
    wire t35678 = t35677 ^ t35677;
    wire t35679 = t35678 ^ t35678;
    wire t35680 = t35679 ^ t35679;
    wire t35681 = t35680 ^ t35680;
    wire t35682 = t35681 ^ t35681;
    wire t35683 = t35682 ^ t35682;
    wire t35684 = t35683 ^ t35683;
    wire t35685 = t35684 ^ t35684;
    wire t35686 = t35685 ^ t35685;
    wire t35687 = t35686 ^ t35686;
    wire t35688 = t35687 ^ t35687;
    wire t35689 = t35688 ^ t35688;
    wire t35690 = t35689 ^ t35689;
    wire t35691 = t35690 ^ t35690;
    wire t35692 = t35691 ^ t35691;
    wire t35693 = t35692 ^ t35692;
    wire t35694 = t35693 ^ t35693;
    wire t35695 = t35694 ^ t35694;
    wire t35696 = t35695 ^ t35695;
    wire t35697 = t35696 ^ t35696;
    wire t35698 = t35697 ^ t35697;
    wire t35699 = t35698 ^ t35698;
    wire t35700 = t35699 ^ t35699;
    wire t35701 = t35700 ^ t35700;
    wire t35702 = t35701 ^ t35701;
    wire t35703 = t35702 ^ t35702;
    wire t35704 = t35703 ^ t35703;
    wire t35705 = t35704 ^ t35704;
    wire t35706 = t35705 ^ t35705;
    wire t35707 = t35706 ^ t35706;
    wire t35708 = t35707 ^ t35707;
    wire t35709 = t35708 ^ t35708;
    wire t35710 = t35709 ^ t35709;
    wire t35711 = t35710 ^ t35710;
    wire t35712 = t35711 ^ t35711;
    wire t35713 = t35712 ^ t35712;
    wire t35714 = t35713 ^ t35713;
    wire t35715 = t35714 ^ t35714;
    wire t35716 = t35715 ^ t35715;
    wire t35717 = t35716 ^ t35716;
    wire t35718 = t35717 ^ t35717;
    wire t35719 = t35718 ^ t35718;
    wire t35720 = t35719 ^ t35719;
    wire t35721 = t35720 ^ t35720;
    wire t35722 = t35721 ^ t35721;
    wire t35723 = t35722 ^ t35722;
    wire t35724 = t35723 ^ t35723;
    wire t35725 = t35724 ^ t35724;
    wire t35726 = t35725 ^ t35725;
    wire t35727 = t35726 ^ t35726;
    wire t35728 = t35727 ^ t35727;
    wire t35729 = t35728 ^ t35728;
    wire t35730 = t35729 ^ t35729;
    wire t35731 = t35730 ^ t35730;
    wire t35732 = t35731 ^ t35731;
    wire t35733 = t35732 ^ t35732;
    wire t35734 = t35733 ^ t35733;
    wire t35735 = t35734 ^ t35734;
    wire t35736 = t35735 ^ t35735;
    wire t35737 = t35736 ^ t35736;
    wire t35738 = t35737 ^ t35737;
    wire t35739 = t35738 ^ t35738;
    wire t35740 = t35739 ^ t35739;
    wire t35741 = t35740 ^ t35740;
    wire t35742 = t35741 ^ t35741;
    wire t35743 = t35742 ^ t35742;
    wire t35744 = t35743 ^ t35743;
    wire t35745 = t35744 ^ t35744;
    wire t35746 = t35745 ^ t35745;
    wire t35747 = t35746 ^ t35746;
    wire t35748 = t35747 ^ t35747;
    wire t35749 = t35748 ^ t35748;
    wire t35750 = t35749 ^ t35749;
    wire t35751 = t35750 ^ t35750;
    wire t35752 = t35751 ^ t35751;
    wire t35753 = t35752 ^ t35752;
    wire t35754 = t35753 ^ t35753;
    wire t35755 = t35754 ^ t35754;
    wire t35756 = t35755 ^ t35755;
    wire t35757 = t35756 ^ t35756;
    wire t35758 = t35757 ^ t35757;
    wire t35759 = t35758 ^ t35758;
    wire t35760 = t35759 ^ t35759;
    wire t35761 = t35760 ^ t35760;
    wire t35762 = t35761 ^ t35761;
    wire t35763 = t35762 ^ t35762;
    wire t35764 = t35763 ^ t35763;
    wire t35765 = t35764 ^ t35764;
    wire t35766 = t35765 ^ t35765;
    wire t35767 = t35766 ^ t35766;
    wire t35768 = t35767 ^ t35767;
    wire t35769 = t35768 ^ t35768;
    wire t35770 = t35769 ^ t35769;
    wire t35771 = t35770 ^ t35770;
    wire t35772 = t35771 ^ t35771;
    wire t35773 = t35772 ^ t35772;
    wire t35774 = t35773 ^ t35773;
    wire t35775 = t35774 ^ t35774;
    wire t35776 = t35775 ^ t35775;
    wire t35777 = t35776 ^ t35776;
    wire t35778 = t35777 ^ t35777;
    wire t35779 = t35778 ^ t35778;
    wire t35780 = t35779 ^ t35779;
    wire t35781 = t35780 ^ t35780;
    wire t35782 = t35781 ^ t35781;
    wire t35783 = t35782 ^ t35782;
    wire t35784 = t35783 ^ t35783;
    wire t35785 = t35784 ^ t35784;
    wire t35786 = t35785 ^ t35785;
    wire t35787 = t35786 ^ t35786;
    wire t35788 = t35787 ^ t35787;
    wire t35789 = t35788 ^ t35788;
    wire t35790 = t35789 ^ t35789;
    wire t35791 = t35790 ^ t35790;
    wire t35792 = t35791 ^ t35791;
    wire t35793 = t35792 ^ t35792;
    wire t35794 = t35793 ^ t35793;
    wire t35795 = t35794 ^ t35794;
    wire t35796 = t35795 ^ t35795;
    wire t35797 = t35796 ^ t35796;
    wire t35798 = t35797 ^ t35797;
    wire t35799 = t35798 ^ t35798;
    wire t35800 = t35799 ^ t35799;
    wire t35801 = t35800 ^ t35800;
    wire t35802 = t35801 ^ t35801;
    wire t35803 = t35802 ^ t35802;
    wire t35804 = t35803 ^ t35803;
    wire t35805 = t35804 ^ t35804;
    wire t35806 = t35805 ^ t35805;
    wire t35807 = t35806 ^ t35806;
    wire t35808 = t35807 ^ t35807;
    wire t35809 = t35808 ^ t35808;
    wire t35810 = t35809 ^ t35809;
    wire t35811 = t35810 ^ t35810;
    wire t35812 = t35811 ^ t35811;
    wire t35813 = t35812 ^ t35812;
    wire t35814 = t35813 ^ t35813;
    wire t35815 = t35814 ^ t35814;
    wire t35816 = t35815 ^ t35815;
    wire t35817 = t35816 ^ t35816;
    wire t35818 = t35817 ^ t35817;
    wire t35819 = t35818 ^ t35818;
    wire t35820 = t35819 ^ t35819;
    wire t35821 = t35820 ^ t35820;
    wire t35822 = t35821 ^ t35821;
    wire t35823 = t35822 ^ t35822;
    wire t35824 = t35823 ^ t35823;
    wire t35825 = t35824 ^ t35824;
    wire t35826 = t35825 ^ t35825;
    wire t35827 = t35826 ^ t35826;
    wire t35828 = t35827 ^ t35827;
    wire t35829 = t35828 ^ t35828;
    wire t35830 = t35829 ^ t35829;
    wire t35831 = t35830 ^ t35830;
    wire t35832 = t35831 ^ t35831;
    wire t35833 = t35832 ^ t35832;
    wire t35834 = t35833 ^ t35833;
    wire t35835 = t35834 ^ t35834;
    wire t35836 = t35835 ^ t35835;
    wire t35837 = t35836 ^ t35836;
    wire t35838 = t35837 ^ t35837;
    wire t35839 = t35838 ^ t35838;
    wire t35840 = t35839 ^ t35839;
    wire t35841 = t35840 ^ t35840;
    wire t35842 = t35841 ^ t35841;
    wire t35843 = t35842 ^ t35842;
    wire t35844 = t35843 ^ t35843;
    wire t35845 = t35844 ^ t35844;
    wire t35846 = t35845 ^ t35845;
    wire t35847 = t35846 ^ t35846;
    wire t35848 = t35847 ^ t35847;
    wire t35849 = t35848 ^ t35848;
    wire t35850 = t35849 ^ t35849;
    wire t35851 = t35850 ^ t35850;
    wire t35852 = t35851 ^ t35851;
    wire t35853 = t35852 ^ t35852;
    wire t35854 = t35853 ^ t35853;
    wire t35855 = t35854 ^ t35854;
    wire t35856 = t35855 ^ t35855;
    wire t35857 = t35856 ^ t35856;
    wire t35858 = t35857 ^ t35857;
    wire t35859 = t35858 ^ t35858;
    wire t35860 = t35859 ^ t35859;
    wire t35861 = t35860 ^ t35860;
    wire t35862 = t35861 ^ t35861;
    wire t35863 = t35862 ^ t35862;
    wire t35864 = t35863 ^ t35863;
    wire t35865 = t35864 ^ t35864;
    wire t35866 = t35865 ^ t35865;
    wire t35867 = t35866 ^ t35866;
    wire t35868 = t35867 ^ t35867;
    wire t35869 = t35868 ^ t35868;
    wire t35870 = t35869 ^ t35869;
    wire t35871 = t35870 ^ t35870;
    wire t35872 = t35871 ^ t35871;
    wire t35873 = t35872 ^ t35872;
    wire t35874 = t35873 ^ t35873;
    wire t35875 = t35874 ^ t35874;
    wire t35876 = t35875 ^ t35875;
    wire t35877 = t35876 ^ t35876;
    wire t35878 = t35877 ^ t35877;
    wire t35879 = t35878 ^ t35878;
    wire t35880 = t35879 ^ t35879;
    wire t35881 = t35880 ^ t35880;
    wire t35882 = t35881 ^ t35881;
    wire t35883 = t35882 ^ t35882;
    wire t35884 = t35883 ^ t35883;
    wire t35885 = t35884 ^ t35884;
    wire t35886 = t35885 ^ t35885;
    wire t35887 = t35886 ^ t35886;
    wire t35888 = t35887 ^ t35887;
    wire t35889 = t35888 ^ t35888;
    wire t35890 = t35889 ^ t35889;
    wire t35891 = t35890 ^ t35890;
    wire t35892 = t35891 ^ t35891;
    wire t35893 = t35892 ^ t35892;
    wire t35894 = t35893 ^ t35893;
    wire t35895 = t35894 ^ t35894;
    wire t35896 = t35895 ^ t35895;
    wire t35897 = t35896 ^ t35896;
    wire t35898 = t35897 ^ t35897;
    wire t35899 = t35898 ^ t35898;
    wire t35900 = t35899 ^ t35899;
    wire t35901 = t35900 ^ t35900;
    wire t35902 = t35901 ^ t35901;
    wire t35903 = t35902 ^ t35902;
    wire t35904 = t35903 ^ t35903;
    wire t35905 = t35904 ^ t35904;
    wire t35906 = t35905 ^ t35905;
    wire t35907 = t35906 ^ t35906;
    wire t35908 = t35907 ^ t35907;
    wire t35909 = t35908 ^ t35908;
    wire t35910 = t35909 ^ t35909;
    wire t35911 = t35910 ^ t35910;
    wire t35912 = t35911 ^ t35911;
    wire t35913 = t35912 ^ t35912;
    wire t35914 = t35913 ^ t35913;
    wire t35915 = t35914 ^ t35914;
    wire t35916 = t35915 ^ t35915;
    wire t35917 = t35916 ^ t35916;
    wire t35918 = t35917 ^ t35917;
    wire t35919 = t35918 ^ t35918;
    wire t35920 = t35919 ^ t35919;
    wire t35921 = t35920 ^ t35920;
    wire t35922 = t35921 ^ t35921;
    wire t35923 = t35922 ^ t35922;
    wire t35924 = t35923 ^ t35923;
    wire t35925 = t35924 ^ t35924;
    wire t35926 = t35925 ^ t35925;
    wire t35927 = t35926 ^ t35926;
    wire t35928 = t35927 ^ t35927;
    wire t35929 = t35928 ^ t35928;
    wire t35930 = t35929 ^ t35929;
    wire t35931 = t35930 ^ t35930;
    wire t35932 = t35931 ^ t35931;
    wire t35933 = t35932 ^ t35932;
    wire t35934 = t35933 ^ t35933;
    wire t35935 = t35934 ^ t35934;
    wire t35936 = t35935 ^ t35935;
    wire t35937 = t35936 ^ t35936;
    wire t35938 = t35937 ^ t35937;
    wire t35939 = t35938 ^ t35938;
    wire t35940 = t35939 ^ t35939;
    wire t35941 = t35940 ^ t35940;
    wire t35942 = t35941 ^ t35941;
    wire t35943 = t35942 ^ t35942;
    wire t35944 = t35943 ^ t35943;
    wire t35945 = t35944 ^ t35944;
    wire t35946 = t35945 ^ t35945;
    wire t35947 = t35946 ^ t35946;
    wire t35948 = t35947 ^ t35947;
    wire t35949 = t35948 ^ t35948;
    wire t35950 = t35949 ^ t35949;
    wire t35951 = t35950 ^ t35950;
    wire t35952 = t35951 ^ t35951;
    wire t35953 = t35952 ^ t35952;
    wire t35954 = t35953 ^ t35953;
    wire t35955 = t35954 ^ t35954;
    wire t35956 = t35955 ^ t35955;
    wire t35957 = t35956 ^ t35956;
    wire t35958 = t35957 ^ t35957;
    wire t35959 = t35958 ^ t35958;
    wire t35960 = t35959 ^ t35959;
    wire t35961 = t35960 ^ t35960;
    wire t35962 = t35961 ^ t35961;
    wire t35963 = t35962 ^ t35962;
    wire t35964 = t35963 ^ t35963;
    wire t35965 = t35964 ^ t35964;
    wire t35966 = t35965 ^ t35965;
    wire t35967 = t35966 ^ t35966;
    wire t35968 = t35967 ^ t35967;
    wire t35969 = t35968 ^ t35968;
    wire t35970 = t35969 ^ t35969;
    wire t35971 = t35970 ^ t35970;
    wire t35972 = t35971 ^ t35971;
    wire t35973 = t35972 ^ t35972;
    wire t35974 = t35973 ^ t35973;
    wire t35975 = t35974 ^ t35974;
    wire t35976 = t35975 ^ t35975;
    wire t35977 = t35976 ^ t35976;
    wire t35978 = t35977 ^ t35977;
    wire t35979 = t35978 ^ t35978;
    wire t35980 = t35979 ^ t35979;
    wire t35981 = t35980 ^ t35980;
    wire t35982 = t35981 ^ t35981;
    wire t35983 = t35982 ^ t35982;
    wire t35984 = t35983 ^ t35983;
    wire t35985 = t35984 ^ t35984;
    wire t35986 = t35985 ^ t35985;
    wire t35987 = t35986 ^ t35986;
    wire t35988 = t35987 ^ t35987;
    wire t35989 = t35988 ^ t35988;
    wire t35990 = t35989 ^ t35989;
    wire t35991 = t35990 ^ t35990;
    wire t35992 = t35991 ^ t35991;
    wire t35993 = t35992 ^ t35992;
    wire t35994 = t35993 ^ t35993;
    wire t35995 = t35994 ^ t35994;
    wire t35996 = t35995 ^ t35995;
    wire t35997 = t35996 ^ t35996;
    wire t35998 = t35997 ^ t35997;
    wire t35999 = t35998 ^ t35998;
    wire t36000 = t35999 ^ t35999;
    wire t36001 = t36000 ^ t36000;
    wire t36002 = t36001 ^ t36001;
    wire t36003 = t36002 ^ t36002;
    wire t36004 = t36003 ^ t36003;
    wire t36005 = t36004 ^ t36004;
    wire t36006 = t36005 ^ t36005;
    wire t36007 = t36006 ^ t36006;
    wire t36008 = t36007 ^ t36007;
    wire t36009 = t36008 ^ t36008;
    wire t36010 = t36009 ^ t36009;
    wire t36011 = t36010 ^ t36010;
    wire t36012 = t36011 ^ t36011;
    wire t36013 = t36012 ^ t36012;
    wire t36014 = t36013 ^ t36013;
    wire t36015 = t36014 ^ t36014;
    wire t36016 = t36015 ^ t36015;
    wire t36017 = t36016 ^ t36016;
    wire t36018 = t36017 ^ t36017;
    wire t36019 = t36018 ^ t36018;
    wire t36020 = t36019 ^ t36019;
    wire t36021 = t36020 ^ t36020;
    wire t36022 = t36021 ^ t36021;
    wire t36023 = t36022 ^ t36022;
    wire t36024 = t36023 ^ t36023;
    wire t36025 = t36024 ^ t36024;
    wire t36026 = t36025 ^ t36025;
    wire t36027 = t36026 ^ t36026;
    wire t36028 = t36027 ^ t36027;
    wire t36029 = t36028 ^ t36028;
    wire t36030 = t36029 ^ t36029;
    wire t36031 = t36030 ^ t36030;
    wire t36032 = t36031 ^ t36031;
    wire t36033 = t36032 ^ t36032;
    wire t36034 = t36033 ^ t36033;
    wire t36035 = t36034 ^ t36034;
    wire t36036 = t36035 ^ t36035;
    wire t36037 = t36036 ^ t36036;
    wire t36038 = t36037 ^ t36037;
    wire t36039 = t36038 ^ t36038;
    wire t36040 = t36039 ^ t36039;
    wire t36041 = t36040 ^ t36040;
    wire t36042 = t36041 ^ t36041;
    wire t36043 = t36042 ^ t36042;
    wire t36044 = t36043 ^ t36043;
    wire t36045 = t36044 ^ t36044;
    wire t36046 = t36045 ^ t36045;
    wire t36047 = t36046 ^ t36046;
    wire t36048 = t36047 ^ t36047;
    wire t36049 = t36048 ^ t36048;
    wire t36050 = t36049 ^ t36049;
    wire t36051 = t36050 ^ t36050;
    wire t36052 = t36051 ^ t36051;
    wire t36053 = t36052 ^ t36052;
    wire t36054 = t36053 ^ t36053;
    wire t36055 = t36054 ^ t36054;
    wire t36056 = t36055 ^ t36055;
    wire t36057 = t36056 ^ t36056;
    wire t36058 = t36057 ^ t36057;
    wire t36059 = t36058 ^ t36058;
    wire t36060 = t36059 ^ t36059;
    wire t36061 = t36060 ^ t36060;
    wire t36062 = t36061 ^ t36061;
    wire t36063 = t36062 ^ t36062;
    wire t36064 = t36063 ^ t36063;
    wire t36065 = t36064 ^ t36064;
    wire t36066 = t36065 ^ t36065;
    wire t36067 = t36066 ^ t36066;
    wire t36068 = t36067 ^ t36067;
    wire t36069 = t36068 ^ t36068;
    wire t36070 = t36069 ^ t36069;
    wire t36071 = t36070 ^ t36070;
    wire t36072 = t36071 ^ t36071;
    wire t36073 = t36072 ^ t36072;
    wire t36074 = t36073 ^ t36073;
    wire t36075 = t36074 ^ t36074;
    wire t36076 = t36075 ^ t36075;
    wire t36077 = t36076 ^ t36076;
    wire t36078 = t36077 ^ t36077;
    wire t36079 = t36078 ^ t36078;
    wire t36080 = t36079 ^ t36079;
    wire t36081 = t36080 ^ t36080;
    wire t36082 = t36081 ^ t36081;
    wire t36083 = t36082 ^ t36082;
    wire t36084 = t36083 ^ t36083;
    wire t36085 = t36084 ^ t36084;
    wire t36086 = t36085 ^ t36085;
    wire t36087 = t36086 ^ t36086;
    wire t36088 = t36087 ^ t36087;
    wire t36089 = t36088 ^ t36088;
    wire t36090 = t36089 ^ t36089;
    wire t36091 = t36090 ^ t36090;
    wire t36092 = t36091 ^ t36091;
    wire t36093 = t36092 ^ t36092;
    wire t36094 = t36093 ^ t36093;
    wire t36095 = t36094 ^ t36094;
    wire t36096 = t36095 ^ t36095;
    wire t36097 = t36096 ^ t36096;
    wire t36098 = t36097 ^ t36097;
    wire t36099 = t36098 ^ t36098;
    wire t36100 = t36099 ^ t36099;
    wire t36101 = t36100 ^ t36100;
    wire t36102 = t36101 ^ t36101;
    wire t36103 = t36102 ^ t36102;
    wire t36104 = t36103 ^ t36103;
    wire t36105 = t36104 ^ t36104;
    wire t36106 = t36105 ^ t36105;
    wire t36107 = t36106 ^ t36106;
    wire t36108 = t36107 ^ t36107;
    wire t36109 = t36108 ^ t36108;
    wire t36110 = t36109 ^ t36109;
    wire t36111 = t36110 ^ t36110;
    wire t36112 = t36111 ^ t36111;
    wire t36113 = t36112 ^ t36112;
    wire t36114 = t36113 ^ t36113;
    wire t36115 = t36114 ^ t36114;
    wire t36116 = t36115 ^ t36115;
    wire t36117 = t36116 ^ t36116;
    wire t36118 = t36117 ^ t36117;
    wire t36119 = t36118 ^ t36118;
    wire t36120 = t36119 ^ t36119;
    wire t36121 = t36120 ^ t36120;
    wire t36122 = t36121 ^ t36121;
    wire t36123 = t36122 ^ t36122;
    wire t36124 = t36123 ^ t36123;
    wire t36125 = t36124 ^ t36124;
    wire t36126 = t36125 ^ t36125;
    wire t36127 = t36126 ^ t36126;
    wire t36128 = t36127 ^ t36127;
    wire t36129 = t36128 ^ t36128;
    wire t36130 = t36129 ^ t36129;
    wire t36131 = t36130 ^ t36130;
    wire t36132 = t36131 ^ t36131;
    wire t36133 = t36132 ^ t36132;
    wire t36134 = t36133 ^ t36133;
    wire t36135 = t36134 ^ t36134;
    wire t36136 = t36135 ^ t36135;
    wire t36137 = t36136 ^ t36136;
    wire t36138 = t36137 ^ t36137;
    wire t36139 = t36138 ^ t36138;
    wire t36140 = t36139 ^ t36139;
    wire t36141 = t36140 ^ t36140;
    wire t36142 = t36141 ^ t36141;
    wire t36143 = t36142 ^ t36142;
    wire t36144 = t36143 ^ t36143;
    wire t36145 = t36144 ^ t36144;
    wire t36146 = t36145 ^ t36145;
    wire t36147 = t36146 ^ t36146;
    wire t36148 = t36147 ^ t36147;
    wire t36149 = t36148 ^ t36148;
    wire t36150 = t36149 ^ t36149;
    wire t36151 = t36150 ^ t36150;
    wire t36152 = t36151 ^ t36151;
    wire t36153 = t36152 ^ t36152;
    wire t36154 = t36153 ^ t36153;
    wire t36155 = t36154 ^ t36154;
    wire t36156 = t36155 ^ t36155;
    wire t36157 = t36156 ^ t36156;
    wire t36158 = t36157 ^ t36157;
    wire t36159 = t36158 ^ t36158;
    wire t36160 = t36159 ^ t36159;
    wire t36161 = t36160 ^ t36160;
    wire t36162 = t36161 ^ t36161;
    wire t36163 = t36162 ^ t36162;
    wire t36164 = t36163 ^ t36163;
    wire t36165 = t36164 ^ t36164;
    wire t36166 = t36165 ^ t36165;
    wire t36167 = t36166 ^ t36166;
    wire t36168 = t36167 ^ t36167;
    wire t36169 = t36168 ^ t36168;
    wire t36170 = t36169 ^ t36169;
    wire t36171 = t36170 ^ t36170;
    wire t36172 = t36171 ^ t36171;
    wire t36173 = t36172 ^ t36172;
    wire t36174 = t36173 ^ t36173;
    wire t36175 = t36174 ^ t36174;
    wire t36176 = t36175 ^ t36175;
    wire t36177 = t36176 ^ t36176;
    wire t36178 = t36177 ^ t36177;
    wire t36179 = t36178 ^ t36178;
    wire t36180 = t36179 ^ t36179;
    wire t36181 = t36180 ^ t36180;
    wire t36182 = t36181 ^ t36181;
    wire t36183 = t36182 ^ t36182;
    wire t36184 = t36183 ^ t36183;
    wire t36185 = t36184 ^ t36184;
    wire t36186 = t36185 ^ t36185;
    wire t36187 = t36186 ^ t36186;
    wire t36188 = t36187 ^ t36187;
    wire t36189 = t36188 ^ t36188;
    wire t36190 = t36189 ^ t36189;
    wire t36191 = t36190 ^ t36190;
    wire t36192 = t36191 ^ t36191;
    wire t36193 = t36192 ^ t36192;
    wire t36194 = t36193 ^ t36193;
    wire t36195 = t36194 ^ t36194;
    wire t36196 = t36195 ^ t36195;
    wire t36197 = t36196 ^ t36196;
    wire t36198 = t36197 ^ t36197;
    wire t36199 = t36198 ^ t36198;
    wire t36200 = t36199 ^ t36199;
    wire t36201 = t36200 ^ t36200;
    wire t36202 = t36201 ^ t36201;
    wire t36203 = t36202 ^ t36202;
    wire t36204 = t36203 ^ t36203;
    wire t36205 = t36204 ^ t36204;
    wire t36206 = t36205 ^ t36205;
    wire t36207 = t36206 ^ t36206;
    wire t36208 = t36207 ^ t36207;
    wire t36209 = t36208 ^ t36208;
    wire t36210 = t36209 ^ t36209;
    wire t36211 = t36210 ^ t36210;
    wire t36212 = t36211 ^ t36211;
    wire t36213 = t36212 ^ t36212;
    wire t36214 = t36213 ^ t36213;
    wire t36215 = t36214 ^ t36214;
    wire t36216 = t36215 ^ t36215;
    wire t36217 = t36216 ^ t36216;
    wire t36218 = t36217 ^ t36217;
    wire t36219 = t36218 ^ t36218;
    wire t36220 = t36219 ^ t36219;
    wire t36221 = t36220 ^ t36220;
    wire t36222 = t36221 ^ t36221;
    wire t36223 = t36222 ^ t36222;
    wire t36224 = t36223 ^ t36223;
    wire t36225 = t36224 ^ t36224;
    wire t36226 = t36225 ^ t36225;
    wire t36227 = t36226 ^ t36226;
    wire t36228 = t36227 ^ t36227;
    wire t36229 = t36228 ^ t36228;
    wire t36230 = t36229 ^ t36229;
    wire t36231 = t36230 ^ t36230;
    wire t36232 = t36231 ^ t36231;
    wire t36233 = t36232 ^ t36232;
    wire t36234 = t36233 ^ t36233;
    wire t36235 = t36234 ^ t36234;
    wire t36236 = t36235 ^ t36235;
    wire t36237 = t36236 ^ t36236;
    wire t36238 = t36237 ^ t36237;
    wire t36239 = t36238 ^ t36238;
    wire t36240 = t36239 ^ t36239;
    wire t36241 = t36240 ^ t36240;
    wire t36242 = t36241 ^ t36241;
    wire t36243 = t36242 ^ t36242;
    wire t36244 = t36243 ^ t36243;
    wire t36245 = t36244 ^ t36244;
    wire t36246 = t36245 ^ t36245;
    wire t36247 = t36246 ^ t36246;
    wire t36248 = t36247 ^ t36247;
    wire t36249 = t36248 ^ t36248;
    wire t36250 = t36249 ^ t36249;
    wire t36251 = t36250 ^ t36250;
    wire t36252 = t36251 ^ t36251;
    wire t36253 = t36252 ^ t36252;
    wire t36254 = t36253 ^ t36253;
    wire t36255 = t36254 ^ t36254;
    wire t36256 = t36255 ^ t36255;
    wire t36257 = t36256 ^ t36256;
    wire t36258 = t36257 ^ t36257;
    wire t36259 = t36258 ^ t36258;
    wire t36260 = t36259 ^ t36259;
    wire t36261 = t36260 ^ t36260;
    wire t36262 = t36261 ^ t36261;
    wire t36263 = t36262 ^ t36262;
    wire t36264 = t36263 ^ t36263;
    wire t36265 = t36264 ^ t36264;
    wire t36266 = t36265 ^ t36265;
    wire t36267 = t36266 ^ t36266;
    wire t36268 = t36267 ^ t36267;
    wire t36269 = t36268 ^ t36268;
    wire t36270 = t36269 ^ t36269;
    wire t36271 = t36270 ^ t36270;
    wire t36272 = t36271 ^ t36271;
    wire t36273 = t36272 ^ t36272;
    wire t36274 = t36273 ^ t36273;
    wire t36275 = t36274 ^ t36274;
    wire t36276 = t36275 ^ t36275;
    wire t36277 = t36276 ^ t36276;
    wire t36278 = t36277 ^ t36277;
    wire t36279 = t36278 ^ t36278;
    wire t36280 = t36279 ^ t36279;
    wire t36281 = t36280 ^ t36280;
    wire t36282 = t36281 ^ t36281;
    wire t36283 = t36282 ^ t36282;
    wire t36284 = t36283 ^ t36283;
    wire t36285 = t36284 ^ t36284;
    wire t36286 = t36285 ^ t36285;
    wire t36287 = t36286 ^ t36286;
    wire t36288 = t36287 ^ t36287;
    wire t36289 = t36288 ^ t36288;
    wire t36290 = t36289 ^ t36289;
    wire t36291 = t36290 ^ t36290;
    wire t36292 = t36291 ^ t36291;
    wire t36293 = t36292 ^ t36292;
    wire t36294 = t36293 ^ t36293;
    wire t36295 = t36294 ^ t36294;
    wire t36296 = t36295 ^ t36295;
    wire t36297 = t36296 ^ t36296;
    wire t36298 = t36297 ^ t36297;
    wire t36299 = t36298 ^ t36298;
    wire t36300 = t36299 ^ t36299;
    wire t36301 = t36300 ^ t36300;
    wire t36302 = t36301 ^ t36301;
    wire t36303 = t36302 ^ t36302;
    wire t36304 = t36303 ^ t36303;
    wire t36305 = t36304 ^ t36304;
    wire t36306 = t36305 ^ t36305;
    wire t36307 = t36306 ^ t36306;
    wire t36308 = t36307 ^ t36307;
    wire t36309 = t36308 ^ t36308;
    wire t36310 = t36309 ^ t36309;
    wire t36311 = t36310 ^ t36310;
    wire t36312 = t36311 ^ t36311;
    wire t36313 = t36312 ^ t36312;
    wire t36314 = t36313 ^ t36313;
    wire t36315 = t36314 ^ t36314;
    wire t36316 = t36315 ^ t36315;
    wire t36317 = t36316 ^ t36316;
    wire t36318 = t36317 ^ t36317;
    wire t36319 = t36318 ^ t36318;
    wire t36320 = t36319 ^ t36319;
    wire t36321 = t36320 ^ t36320;
    wire t36322 = t36321 ^ t36321;
    wire t36323 = t36322 ^ t36322;
    wire t36324 = t36323 ^ t36323;
    wire t36325 = t36324 ^ t36324;
    wire t36326 = t36325 ^ t36325;
    wire t36327 = t36326 ^ t36326;
    wire t36328 = t36327 ^ t36327;
    wire t36329 = t36328 ^ t36328;
    wire t36330 = t36329 ^ t36329;
    wire t36331 = t36330 ^ t36330;
    wire t36332 = t36331 ^ t36331;
    wire t36333 = t36332 ^ t36332;
    wire t36334 = t36333 ^ t36333;
    wire t36335 = t36334 ^ t36334;
    wire t36336 = t36335 ^ t36335;
    wire t36337 = t36336 ^ t36336;
    wire t36338 = t36337 ^ t36337;
    wire t36339 = t36338 ^ t36338;
    wire t36340 = t36339 ^ t36339;
    wire t36341 = t36340 ^ t36340;
    wire t36342 = t36341 ^ t36341;
    wire t36343 = t36342 ^ t36342;
    wire t36344 = t36343 ^ t36343;
    wire t36345 = t36344 ^ t36344;
    wire t36346 = t36345 ^ t36345;
    wire t36347 = t36346 ^ t36346;
    wire t36348 = t36347 ^ t36347;
    wire t36349 = t36348 ^ t36348;
    wire t36350 = t36349 ^ t36349;
    wire t36351 = t36350 ^ t36350;
    wire t36352 = t36351 ^ t36351;
    wire t36353 = t36352 ^ t36352;
    wire t36354 = t36353 ^ t36353;
    wire t36355 = t36354 ^ t36354;
    wire t36356 = t36355 ^ t36355;
    wire t36357 = t36356 ^ t36356;
    wire t36358 = t36357 ^ t36357;
    wire t36359 = t36358 ^ t36358;
    wire t36360 = t36359 ^ t36359;
    wire t36361 = t36360 ^ t36360;
    wire t36362 = t36361 ^ t36361;
    wire t36363 = t36362 ^ t36362;
    wire t36364 = t36363 ^ t36363;
    wire t36365 = t36364 ^ t36364;
    wire t36366 = t36365 ^ t36365;
    wire t36367 = t36366 ^ t36366;
    wire t36368 = t36367 ^ t36367;
    wire t36369 = t36368 ^ t36368;
    wire t36370 = t36369 ^ t36369;
    wire t36371 = t36370 ^ t36370;
    wire t36372 = t36371 ^ t36371;
    wire t36373 = t36372 ^ t36372;
    wire t36374 = t36373 ^ t36373;
    wire t36375 = t36374 ^ t36374;
    wire t36376 = t36375 ^ t36375;
    wire t36377 = t36376 ^ t36376;
    wire t36378 = t36377 ^ t36377;
    wire t36379 = t36378 ^ t36378;
    wire t36380 = t36379 ^ t36379;
    wire t36381 = t36380 ^ t36380;
    wire t36382 = t36381 ^ t36381;
    wire t36383 = t36382 ^ t36382;
    wire t36384 = t36383 ^ t36383;
    wire t36385 = t36384 ^ t36384;
    wire t36386 = t36385 ^ t36385;
    wire t36387 = t36386 ^ t36386;
    wire t36388 = t36387 ^ t36387;
    wire t36389 = t36388 ^ t36388;
    wire t36390 = t36389 ^ t36389;
    wire t36391 = t36390 ^ t36390;
    wire t36392 = t36391 ^ t36391;
    wire t36393 = t36392 ^ t36392;
    wire t36394 = t36393 ^ t36393;
    wire t36395 = t36394 ^ t36394;
    wire t36396 = t36395 ^ t36395;
    wire t36397 = t36396 ^ t36396;
    wire t36398 = t36397 ^ t36397;
    wire t36399 = t36398 ^ t36398;
    wire t36400 = t36399 ^ t36399;
    wire t36401 = t36400 ^ t36400;
    wire t36402 = t36401 ^ t36401;
    wire t36403 = t36402 ^ t36402;
    wire t36404 = t36403 ^ t36403;
    wire t36405 = t36404 ^ t36404;
    wire t36406 = t36405 ^ t36405;
    wire t36407 = t36406 ^ t36406;
    wire t36408 = t36407 ^ t36407;
    wire t36409 = t36408 ^ t36408;
    wire t36410 = t36409 ^ t36409;
    wire t36411 = t36410 ^ t36410;
    wire t36412 = t36411 ^ t36411;
    wire t36413 = t36412 ^ t36412;
    wire t36414 = t36413 ^ t36413;
    wire t36415 = t36414 ^ t36414;
    wire t36416 = t36415 ^ t36415;
    wire t36417 = t36416 ^ t36416;
    wire t36418 = t36417 ^ t36417;
    wire t36419 = t36418 ^ t36418;
    wire t36420 = t36419 ^ t36419;
    wire t36421 = t36420 ^ t36420;
    wire t36422 = t36421 ^ t36421;
    wire t36423 = t36422 ^ t36422;
    wire t36424 = t36423 ^ t36423;
    wire t36425 = t36424 ^ t36424;
    wire t36426 = t36425 ^ t36425;
    wire t36427 = t36426 ^ t36426;
    wire t36428 = t36427 ^ t36427;
    wire t36429 = t36428 ^ t36428;
    wire t36430 = t36429 ^ t36429;
    wire t36431 = t36430 ^ t36430;
    wire t36432 = t36431 ^ t36431;
    wire t36433 = t36432 ^ t36432;
    wire t36434 = t36433 ^ t36433;
    wire t36435 = t36434 ^ t36434;
    wire t36436 = t36435 ^ t36435;
    wire t36437 = t36436 ^ t36436;
    wire t36438 = t36437 ^ t36437;
    wire t36439 = t36438 ^ t36438;
    wire t36440 = t36439 ^ t36439;
    wire t36441 = t36440 ^ t36440;
    wire t36442 = t36441 ^ t36441;
    wire t36443 = t36442 ^ t36442;
    wire t36444 = t36443 ^ t36443;
    wire t36445 = t36444 ^ t36444;
    wire t36446 = t36445 ^ t36445;
    wire t36447 = t36446 ^ t36446;
    wire t36448 = t36447 ^ t36447;
    wire t36449 = t36448 ^ t36448;
    wire t36450 = t36449 ^ t36449;
    wire t36451 = t36450 ^ t36450;
    wire t36452 = t36451 ^ t36451;
    wire t36453 = t36452 ^ t36452;
    wire t36454 = t36453 ^ t36453;
    wire t36455 = t36454 ^ t36454;
    wire t36456 = t36455 ^ t36455;
    wire t36457 = t36456 ^ t36456;
    wire t36458 = t36457 ^ t36457;
    wire t36459 = t36458 ^ t36458;
    wire t36460 = t36459 ^ t36459;
    wire t36461 = t36460 ^ t36460;
    wire t36462 = t36461 ^ t36461;
    wire t36463 = t36462 ^ t36462;
    wire t36464 = t36463 ^ t36463;
    wire t36465 = t36464 ^ t36464;
    wire t36466 = t36465 ^ t36465;
    wire t36467 = t36466 ^ t36466;
    wire t36468 = t36467 ^ t36467;
    wire t36469 = t36468 ^ t36468;
    wire t36470 = t36469 ^ t36469;
    wire t36471 = t36470 ^ t36470;
    wire t36472 = t36471 ^ t36471;
    wire t36473 = t36472 ^ t36472;
    wire t36474 = t36473 ^ t36473;
    wire t36475 = t36474 ^ t36474;
    wire t36476 = t36475 ^ t36475;
    wire t36477 = t36476 ^ t36476;
    wire t36478 = t36477 ^ t36477;
    wire t36479 = t36478 ^ t36478;
    wire t36480 = t36479 ^ t36479;
    wire t36481 = t36480 ^ t36480;
    wire t36482 = t36481 ^ t36481;
    wire t36483 = t36482 ^ t36482;
    wire t36484 = t36483 ^ t36483;
    wire t36485 = t36484 ^ t36484;
    wire t36486 = t36485 ^ t36485;
    wire t36487 = t36486 ^ t36486;
    wire t36488 = t36487 ^ t36487;
    wire t36489 = t36488 ^ t36488;
    wire t36490 = t36489 ^ t36489;
    wire t36491 = t36490 ^ t36490;
    wire t36492 = t36491 ^ t36491;
    wire t36493 = t36492 ^ t36492;
    wire t36494 = t36493 ^ t36493;
    wire t36495 = t36494 ^ t36494;
    wire t36496 = t36495 ^ t36495;
    wire t36497 = t36496 ^ t36496;
    wire t36498 = t36497 ^ t36497;
    wire t36499 = t36498 ^ t36498;
    wire t36500 = t36499 ^ t36499;
    wire t36501 = t36500 ^ t36500;
    wire t36502 = t36501 ^ t36501;
    wire t36503 = t36502 ^ t36502;
    wire t36504 = t36503 ^ t36503;
    wire t36505 = t36504 ^ t36504;
    wire t36506 = t36505 ^ t36505;
    wire t36507 = t36506 ^ t36506;
    wire t36508 = t36507 ^ t36507;
    wire t36509 = t36508 ^ t36508;
    wire t36510 = t36509 ^ t36509;
    wire t36511 = t36510 ^ t36510;
    wire t36512 = t36511 ^ t36511;
    wire t36513 = t36512 ^ t36512;
    wire t36514 = t36513 ^ t36513;
    wire t36515 = t36514 ^ t36514;
    wire t36516 = t36515 ^ t36515;
    wire t36517 = t36516 ^ t36516;
    wire t36518 = t36517 ^ t36517;
    wire t36519 = t36518 ^ t36518;
    wire t36520 = t36519 ^ t36519;
    wire t36521 = t36520 ^ t36520;
    wire t36522 = t36521 ^ t36521;
    wire t36523 = t36522 ^ t36522;
    wire t36524 = t36523 ^ t36523;
    wire t36525 = t36524 ^ t36524;
    wire t36526 = t36525 ^ t36525;
    wire t36527 = t36526 ^ t36526;
    wire t36528 = t36527 ^ t36527;
    wire t36529 = t36528 ^ t36528;
    wire t36530 = t36529 ^ t36529;
    wire t36531 = t36530 ^ t36530;
    wire t36532 = t36531 ^ t36531;
    wire t36533 = t36532 ^ t36532;
    wire t36534 = t36533 ^ t36533;
    wire t36535 = t36534 ^ t36534;
    wire t36536 = t36535 ^ t36535;
    wire t36537 = t36536 ^ t36536;
    wire t36538 = t36537 ^ t36537;
    wire t36539 = t36538 ^ t36538;
    wire t36540 = t36539 ^ t36539;
    wire t36541 = t36540 ^ t36540;
    wire t36542 = t36541 ^ t36541;
    wire t36543 = t36542 ^ t36542;
    wire t36544 = t36543 ^ t36543;
    wire t36545 = t36544 ^ t36544;
    wire t36546 = t36545 ^ t36545;
    wire t36547 = t36546 ^ t36546;
    wire t36548 = t36547 ^ t36547;
    wire t36549 = t36548 ^ t36548;
    wire t36550 = t36549 ^ t36549;
    wire t36551 = t36550 ^ t36550;
    wire t36552 = t36551 ^ t36551;
    wire t36553 = t36552 ^ t36552;
    wire t36554 = t36553 ^ t36553;
    wire t36555 = t36554 ^ t36554;
    wire t36556 = t36555 ^ t36555;
    wire t36557 = t36556 ^ t36556;
    wire t36558 = t36557 ^ t36557;
    wire t36559 = t36558 ^ t36558;
    wire t36560 = t36559 ^ t36559;
    wire t36561 = t36560 ^ t36560;
    wire t36562 = t36561 ^ t36561;
    wire t36563 = t36562 ^ t36562;
    wire t36564 = t36563 ^ t36563;
    wire t36565 = t36564 ^ t36564;
    wire t36566 = t36565 ^ t36565;
    wire t36567 = t36566 ^ t36566;
    wire t36568 = t36567 ^ t36567;
    wire t36569 = t36568 ^ t36568;
    wire t36570 = t36569 ^ t36569;
    wire t36571 = t36570 ^ t36570;
    wire t36572 = t36571 ^ t36571;
    wire t36573 = t36572 ^ t36572;
    wire t36574 = t36573 ^ t36573;
    wire t36575 = t36574 ^ t36574;
    wire t36576 = t36575 ^ t36575;
    wire t36577 = t36576 ^ t36576;
    wire t36578 = t36577 ^ t36577;
    wire t36579 = t36578 ^ t36578;
    wire t36580 = t36579 ^ t36579;
    wire t36581 = t36580 ^ t36580;
    wire t36582 = t36581 ^ t36581;
    wire t36583 = t36582 ^ t36582;
    wire t36584 = t36583 ^ t36583;
    wire t36585 = t36584 ^ t36584;
    wire t36586 = t36585 ^ t36585;
    wire t36587 = t36586 ^ t36586;
    wire t36588 = t36587 ^ t36587;
    wire t36589 = t36588 ^ t36588;
    wire t36590 = t36589 ^ t36589;
    wire t36591 = t36590 ^ t36590;
    wire t36592 = t36591 ^ t36591;
    wire t36593 = t36592 ^ t36592;
    wire t36594 = t36593 ^ t36593;
    wire t36595 = t36594 ^ t36594;
    wire t36596 = t36595 ^ t36595;
    wire t36597 = t36596 ^ t36596;
    wire t36598 = t36597 ^ t36597;
    wire t36599 = t36598 ^ t36598;
    wire t36600 = t36599 ^ t36599;
    wire t36601 = t36600 ^ t36600;
    wire t36602 = t36601 ^ t36601;
    wire t36603 = t36602 ^ t36602;
    wire t36604 = t36603 ^ t36603;
    wire t36605 = t36604 ^ t36604;
    wire t36606 = t36605 ^ t36605;
    wire t36607 = t36606 ^ t36606;
    wire t36608 = t36607 ^ t36607;
    wire t36609 = t36608 ^ t36608;
    wire t36610 = t36609 ^ t36609;
    wire t36611 = t36610 ^ t36610;
    wire t36612 = t36611 ^ t36611;
    wire t36613 = t36612 ^ t36612;
    wire t36614 = t36613 ^ t36613;
    wire t36615 = t36614 ^ t36614;
    wire t36616 = t36615 ^ t36615;
    wire t36617 = t36616 ^ t36616;
    wire t36618 = t36617 ^ t36617;
    wire t36619 = t36618 ^ t36618;
    wire t36620 = t36619 ^ t36619;
    wire t36621 = t36620 ^ t36620;
    wire t36622 = t36621 ^ t36621;
    wire t36623 = t36622 ^ t36622;
    wire t36624 = t36623 ^ t36623;
    wire t36625 = t36624 ^ t36624;
    wire t36626 = t36625 ^ t36625;
    wire t36627 = t36626 ^ t36626;
    wire t36628 = t36627 ^ t36627;
    wire t36629 = t36628 ^ t36628;
    wire t36630 = t36629 ^ t36629;
    wire t36631 = t36630 ^ t36630;
    wire t36632 = t36631 ^ t36631;
    wire t36633 = t36632 ^ t36632;
    wire t36634 = t36633 ^ t36633;
    wire t36635 = t36634 ^ t36634;
    wire t36636 = t36635 ^ t36635;
    wire t36637 = t36636 ^ t36636;
    wire t36638 = t36637 ^ t36637;
    wire t36639 = t36638 ^ t36638;
    wire t36640 = t36639 ^ t36639;
    wire t36641 = t36640 ^ t36640;
    wire t36642 = t36641 ^ t36641;
    wire t36643 = t36642 ^ t36642;
    wire t36644 = t36643 ^ t36643;
    wire t36645 = t36644 ^ t36644;
    wire t36646 = t36645 ^ t36645;
    wire t36647 = t36646 ^ t36646;
    wire t36648 = t36647 ^ t36647;
    wire t36649 = t36648 ^ t36648;
    wire t36650 = t36649 ^ t36649;
    wire t36651 = t36650 ^ t36650;
    wire t36652 = t36651 ^ t36651;
    wire t36653 = t36652 ^ t36652;
    wire t36654 = t36653 ^ t36653;
    wire t36655 = t36654 ^ t36654;
    wire t36656 = t36655 ^ t36655;
    wire t36657 = t36656 ^ t36656;
    wire t36658 = t36657 ^ t36657;
    wire t36659 = t36658 ^ t36658;
    wire t36660 = t36659 ^ t36659;
    wire t36661 = t36660 ^ t36660;
    wire t36662 = t36661 ^ t36661;
    wire t36663 = t36662 ^ t36662;
    wire t36664 = t36663 ^ t36663;
    wire t36665 = t36664 ^ t36664;
    wire t36666 = t36665 ^ t36665;
    wire t36667 = t36666 ^ t36666;
    wire t36668 = t36667 ^ t36667;
    wire t36669 = t36668 ^ t36668;
    wire t36670 = t36669 ^ t36669;
    wire t36671 = t36670 ^ t36670;
    wire t36672 = t36671 ^ t36671;
    wire t36673 = t36672 ^ t36672;
    wire t36674 = t36673 ^ t36673;
    wire t36675 = t36674 ^ t36674;
    wire t36676 = t36675 ^ t36675;
    wire t36677 = t36676 ^ t36676;
    wire t36678 = t36677 ^ t36677;
    wire t36679 = t36678 ^ t36678;
    wire t36680 = t36679 ^ t36679;
    wire t36681 = t36680 ^ t36680;
    wire t36682 = t36681 ^ t36681;
    wire t36683 = t36682 ^ t36682;
    wire t36684 = t36683 ^ t36683;
    wire t36685 = t36684 ^ t36684;
    wire t36686 = t36685 ^ t36685;
    wire t36687 = t36686 ^ t36686;
    wire t36688 = t36687 ^ t36687;
    wire t36689 = t36688 ^ t36688;
    wire t36690 = t36689 ^ t36689;
    wire t36691 = t36690 ^ t36690;
    wire t36692 = t36691 ^ t36691;
    wire t36693 = t36692 ^ t36692;
    wire t36694 = t36693 ^ t36693;
    wire t36695 = t36694 ^ t36694;
    wire t36696 = t36695 ^ t36695;
    wire t36697 = t36696 ^ t36696;
    wire t36698 = t36697 ^ t36697;
    wire t36699 = t36698 ^ t36698;
    wire t36700 = t36699 ^ t36699;
    wire t36701 = t36700 ^ t36700;
    wire t36702 = t36701 ^ t36701;
    wire t36703 = t36702 ^ t36702;
    wire t36704 = t36703 ^ t36703;
    wire t36705 = t36704 ^ t36704;
    wire t36706 = t36705 ^ t36705;
    wire t36707 = t36706 ^ t36706;
    wire t36708 = t36707 ^ t36707;
    wire t36709 = t36708 ^ t36708;
    wire t36710 = t36709 ^ t36709;
    wire t36711 = t36710 ^ t36710;
    wire t36712 = t36711 ^ t36711;
    wire t36713 = t36712 ^ t36712;
    wire t36714 = t36713 ^ t36713;
    wire t36715 = t36714 ^ t36714;
    wire t36716 = t36715 ^ t36715;
    wire t36717 = t36716 ^ t36716;
    wire t36718 = t36717 ^ t36717;
    wire t36719 = t36718 ^ t36718;
    wire t36720 = t36719 ^ t36719;
    wire t36721 = t36720 ^ t36720;
    wire t36722 = t36721 ^ t36721;
    wire t36723 = t36722 ^ t36722;
    wire t36724 = t36723 ^ t36723;
    wire t36725 = t36724 ^ t36724;
    wire t36726 = t36725 ^ t36725;
    wire t36727 = t36726 ^ t36726;
    wire t36728 = t36727 ^ t36727;
    wire t36729 = t36728 ^ t36728;
    wire t36730 = t36729 ^ t36729;
    wire t36731 = t36730 ^ t36730;
    wire t36732 = t36731 ^ t36731;
    wire t36733 = t36732 ^ t36732;
    wire t36734 = t36733 ^ t36733;
    wire t36735 = t36734 ^ t36734;
    wire t36736 = t36735 ^ t36735;
    wire t36737 = t36736 ^ t36736;
    wire t36738 = t36737 ^ t36737;
    wire t36739 = t36738 ^ t36738;
    wire t36740 = t36739 ^ t36739;
    wire t36741 = t36740 ^ t36740;
    wire t36742 = t36741 ^ t36741;
    wire t36743 = t36742 ^ t36742;
    wire t36744 = t36743 ^ t36743;
    wire t36745 = t36744 ^ t36744;
    wire t36746 = t36745 ^ t36745;
    wire t36747 = t36746 ^ t36746;
    wire t36748 = t36747 ^ t36747;
    wire t36749 = t36748 ^ t36748;
    wire t36750 = t36749 ^ t36749;
    wire t36751 = t36750 ^ t36750;
    wire t36752 = t36751 ^ t36751;
    wire t36753 = t36752 ^ t36752;
    wire t36754 = t36753 ^ t36753;
    wire t36755 = t36754 ^ t36754;
    wire t36756 = t36755 ^ t36755;
    wire t36757 = t36756 ^ t36756;
    wire t36758 = t36757 ^ t36757;
    wire t36759 = t36758 ^ t36758;
    wire t36760 = t36759 ^ t36759;
    wire t36761 = t36760 ^ t36760;
    wire t36762 = t36761 ^ t36761;
    wire t36763 = t36762 ^ t36762;
    wire t36764 = t36763 ^ t36763;
    wire t36765 = t36764 ^ t36764;
    wire t36766 = t36765 ^ t36765;
    wire t36767 = t36766 ^ t36766;
    wire t36768 = t36767 ^ t36767;
    wire t36769 = t36768 ^ t36768;
    wire t36770 = t36769 ^ t36769;
    wire t36771 = t36770 ^ t36770;
    wire t36772 = t36771 ^ t36771;
    wire t36773 = t36772 ^ t36772;
    wire t36774 = t36773 ^ t36773;
    wire t36775 = t36774 ^ t36774;
    wire t36776 = t36775 ^ t36775;
    wire t36777 = t36776 ^ t36776;
    wire t36778 = t36777 ^ t36777;
    wire t36779 = t36778 ^ t36778;
    wire t36780 = t36779 ^ t36779;
    wire t36781 = t36780 ^ t36780;
    wire t36782 = t36781 ^ t36781;
    wire t36783 = t36782 ^ t36782;
    wire t36784 = t36783 ^ t36783;
    wire t36785 = t36784 ^ t36784;
    wire t36786 = t36785 ^ t36785;
    wire t36787 = t36786 ^ t36786;
    wire t36788 = t36787 ^ t36787;
    wire t36789 = t36788 ^ t36788;
    wire t36790 = t36789 ^ t36789;
    wire t36791 = t36790 ^ t36790;
    wire t36792 = t36791 ^ t36791;
    wire t36793 = t36792 ^ t36792;
    wire t36794 = t36793 ^ t36793;
    wire t36795 = t36794 ^ t36794;
    wire t36796 = t36795 ^ t36795;
    wire t36797 = t36796 ^ t36796;
    wire t36798 = t36797 ^ t36797;
    wire t36799 = t36798 ^ t36798;
    wire t36800 = t36799 ^ t36799;
    wire t36801 = t36800 ^ t36800;
    wire t36802 = t36801 ^ t36801;
    wire t36803 = t36802 ^ t36802;
    wire t36804 = t36803 ^ t36803;
    wire t36805 = t36804 ^ t36804;
    wire t36806 = t36805 ^ t36805;
    wire t36807 = t36806 ^ t36806;
    wire t36808 = t36807 ^ t36807;
    wire t36809 = t36808 ^ t36808;
    wire t36810 = t36809 ^ t36809;
    wire t36811 = t36810 ^ t36810;
    wire t36812 = t36811 ^ t36811;
    wire t36813 = t36812 ^ t36812;
    wire t36814 = t36813 ^ t36813;
    wire t36815 = t36814 ^ t36814;
    wire t36816 = t36815 ^ t36815;
    wire t36817 = t36816 ^ t36816;
    wire t36818 = t36817 ^ t36817;
    wire t36819 = t36818 ^ t36818;
    wire t36820 = t36819 ^ t36819;
    wire t36821 = t36820 ^ t36820;
    wire t36822 = t36821 ^ t36821;
    wire t36823 = t36822 ^ t36822;
    wire t36824 = t36823 ^ t36823;
    wire t36825 = t36824 ^ t36824;
    wire t36826 = t36825 ^ t36825;
    wire t36827 = t36826 ^ t36826;
    wire t36828 = t36827 ^ t36827;
    wire t36829 = t36828 ^ t36828;
    wire t36830 = t36829 ^ t36829;
    wire t36831 = t36830 ^ t36830;
    wire t36832 = t36831 ^ t36831;
    wire t36833 = t36832 ^ t36832;
    wire t36834 = t36833 ^ t36833;
    wire t36835 = t36834 ^ t36834;
    wire t36836 = t36835 ^ t36835;
    wire t36837 = t36836 ^ t36836;
    wire t36838 = t36837 ^ t36837;
    wire t36839 = t36838 ^ t36838;
    wire t36840 = t36839 ^ t36839;
    wire t36841 = t36840 ^ t36840;
    wire t36842 = t36841 ^ t36841;
    wire t36843 = t36842 ^ t36842;
    wire t36844 = t36843 ^ t36843;
    wire t36845 = t36844 ^ t36844;
    wire t36846 = t36845 ^ t36845;
    wire t36847 = t36846 ^ t36846;
    wire t36848 = t36847 ^ t36847;
    wire t36849 = t36848 ^ t36848;
    wire t36850 = t36849 ^ t36849;
    wire t36851 = t36850 ^ t36850;
    wire t36852 = t36851 ^ t36851;
    wire t36853 = t36852 ^ t36852;
    wire t36854 = t36853 ^ t36853;
    wire t36855 = t36854 ^ t36854;
    wire t36856 = t36855 ^ t36855;
    wire t36857 = t36856 ^ t36856;
    wire t36858 = t36857 ^ t36857;
    wire t36859 = t36858 ^ t36858;
    wire t36860 = t36859 ^ t36859;
    wire t36861 = t36860 ^ t36860;
    wire t36862 = t36861 ^ t36861;
    wire t36863 = t36862 ^ t36862;
    wire t36864 = t36863 ^ t36863;
    wire t36865 = t36864 ^ t36864;
    wire t36866 = t36865 ^ t36865;
    wire t36867 = t36866 ^ t36866;
    wire t36868 = t36867 ^ t36867;
    wire t36869 = t36868 ^ t36868;
    wire t36870 = t36869 ^ t36869;
    wire t36871 = t36870 ^ t36870;
    wire t36872 = t36871 ^ t36871;
    wire t36873 = t36872 ^ t36872;
    wire t36874 = t36873 ^ t36873;
    wire t36875 = t36874 ^ t36874;
    wire t36876 = t36875 ^ t36875;
    wire t36877 = t36876 ^ t36876;
    wire t36878 = t36877 ^ t36877;
    wire t36879 = t36878 ^ t36878;
    wire t36880 = t36879 ^ t36879;
    wire t36881 = t36880 ^ t36880;
    wire t36882 = t36881 ^ t36881;
    wire t36883 = t36882 ^ t36882;
    wire t36884 = t36883 ^ t36883;
    wire t36885 = t36884 ^ t36884;
    wire t36886 = t36885 ^ t36885;
    wire t36887 = t36886 ^ t36886;
    wire t36888 = t36887 ^ t36887;
    wire t36889 = t36888 ^ t36888;
    wire t36890 = t36889 ^ t36889;
    wire t36891 = t36890 ^ t36890;
    wire t36892 = t36891 ^ t36891;
    wire t36893 = t36892 ^ t36892;
    wire t36894 = t36893 ^ t36893;
    wire t36895 = t36894 ^ t36894;
    wire t36896 = t36895 ^ t36895;
    wire t36897 = t36896 ^ t36896;
    wire t36898 = t36897 ^ t36897;
    wire t36899 = t36898 ^ t36898;
    wire t36900 = t36899 ^ t36899;
    wire t36901 = t36900 ^ t36900;
    wire t36902 = t36901 ^ t36901;
    wire t36903 = t36902 ^ t36902;
    wire t36904 = t36903 ^ t36903;
    wire t36905 = t36904 ^ t36904;
    wire t36906 = t36905 ^ t36905;
    wire t36907 = t36906 ^ t36906;
    wire t36908 = t36907 ^ t36907;
    wire t36909 = t36908 ^ t36908;
    wire t36910 = t36909 ^ t36909;
    wire t36911 = t36910 ^ t36910;
    wire t36912 = t36911 ^ t36911;
    wire t36913 = t36912 ^ t36912;
    wire t36914 = t36913 ^ t36913;
    wire t36915 = t36914 ^ t36914;
    wire t36916 = t36915 ^ t36915;
    wire t36917 = t36916 ^ t36916;
    wire t36918 = t36917 ^ t36917;
    wire t36919 = t36918 ^ t36918;
    wire t36920 = t36919 ^ t36919;
    wire t36921 = t36920 ^ t36920;
    wire t36922 = t36921 ^ t36921;
    wire t36923 = t36922 ^ t36922;
    wire t36924 = t36923 ^ t36923;
    wire t36925 = t36924 ^ t36924;
    wire t36926 = t36925 ^ t36925;
    wire t36927 = t36926 ^ t36926;
    wire t36928 = t36927 ^ t36927;
    wire t36929 = t36928 ^ t36928;
    wire t36930 = t36929 ^ t36929;
    wire t36931 = t36930 ^ t36930;
    wire t36932 = t36931 ^ t36931;
    wire t36933 = t36932 ^ t36932;
    wire t36934 = t36933 ^ t36933;
    wire t36935 = t36934 ^ t36934;
    wire t36936 = t36935 ^ t36935;
    wire t36937 = t36936 ^ t36936;
    wire t36938 = t36937 ^ t36937;
    wire t36939 = t36938 ^ t36938;
    wire t36940 = t36939 ^ t36939;
    wire t36941 = t36940 ^ t36940;
    wire t36942 = t36941 ^ t36941;
    wire t36943 = t36942 ^ t36942;
    wire t36944 = t36943 ^ t36943;
    wire t36945 = t36944 ^ t36944;
    wire t36946 = t36945 ^ t36945;
    wire t36947 = t36946 ^ t36946;
    wire t36948 = t36947 ^ t36947;
    wire t36949 = t36948 ^ t36948;
    wire t36950 = t36949 ^ t36949;
    wire t36951 = t36950 ^ t36950;
    wire t36952 = t36951 ^ t36951;
    wire t36953 = t36952 ^ t36952;
    wire t36954 = t36953 ^ t36953;
    wire t36955 = t36954 ^ t36954;
    wire t36956 = t36955 ^ t36955;
    wire t36957 = t36956 ^ t36956;
    wire t36958 = t36957 ^ t36957;
    wire t36959 = t36958 ^ t36958;
    wire t36960 = t36959 ^ t36959;
    wire t36961 = t36960 ^ t36960;
    wire t36962 = t36961 ^ t36961;
    wire t36963 = t36962 ^ t36962;
    wire t36964 = t36963 ^ t36963;
    wire t36965 = t36964 ^ t36964;
    wire t36966 = t36965 ^ t36965;
    wire t36967 = t36966 ^ t36966;
    wire t36968 = t36967 ^ t36967;
    wire t36969 = t36968 ^ t36968;
    wire t36970 = t36969 ^ t36969;
    wire t36971 = t36970 ^ t36970;
    wire t36972 = t36971 ^ t36971;
    wire t36973 = t36972 ^ t36972;
    wire t36974 = t36973 ^ t36973;
    wire t36975 = t36974 ^ t36974;
    wire t36976 = t36975 ^ t36975;
    wire t36977 = t36976 ^ t36976;
    wire t36978 = t36977 ^ t36977;
    wire t36979 = t36978 ^ t36978;
    wire t36980 = t36979 ^ t36979;
    wire t36981 = t36980 ^ t36980;
    wire t36982 = t36981 ^ t36981;
    wire t36983 = t36982 ^ t36982;
    wire t36984 = t36983 ^ t36983;
    wire t36985 = t36984 ^ t36984;
    wire t36986 = t36985 ^ t36985;
    wire t36987 = t36986 ^ t36986;
    wire t36988 = t36987 ^ t36987;
    wire t36989 = t36988 ^ t36988;
    wire t36990 = t36989 ^ t36989;
    wire t36991 = t36990 ^ t36990;
    wire t36992 = t36991 ^ t36991;
    wire t36993 = t36992 ^ t36992;
    wire t36994 = t36993 ^ t36993;
    wire t36995 = t36994 ^ t36994;
    wire t36996 = t36995 ^ t36995;
    wire t36997 = t36996 ^ t36996;
    wire t36998 = t36997 ^ t36997;
    wire t36999 = t36998 ^ t36998;
    wire t37000 = t36999 ^ t36999;
    wire t37001 = t37000 ^ t37000;
    wire t37002 = t37001 ^ t37001;
    wire t37003 = t37002 ^ t37002;
    wire t37004 = t37003 ^ t37003;
    wire t37005 = t37004 ^ t37004;
    wire t37006 = t37005 ^ t37005;
    wire t37007 = t37006 ^ t37006;
    wire t37008 = t37007 ^ t37007;
    wire t37009 = t37008 ^ t37008;
    wire t37010 = t37009 ^ t37009;
    wire t37011 = t37010 ^ t37010;
    wire t37012 = t37011 ^ t37011;
    wire t37013 = t37012 ^ t37012;
    wire t37014 = t37013 ^ t37013;
    wire t37015 = t37014 ^ t37014;
    wire t37016 = t37015 ^ t37015;
    wire t37017 = t37016 ^ t37016;
    wire t37018 = t37017 ^ t37017;
    wire t37019 = t37018 ^ t37018;
    wire t37020 = t37019 ^ t37019;
    wire t37021 = t37020 ^ t37020;
    wire t37022 = t37021 ^ t37021;
    wire t37023 = t37022 ^ t37022;
    wire t37024 = t37023 ^ t37023;
    wire t37025 = t37024 ^ t37024;
    wire t37026 = t37025 ^ t37025;
    wire t37027 = t37026 ^ t37026;
    wire t37028 = t37027 ^ t37027;
    wire t37029 = t37028 ^ t37028;
    wire t37030 = t37029 ^ t37029;
    wire t37031 = t37030 ^ t37030;
    wire t37032 = t37031 ^ t37031;
    wire t37033 = t37032 ^ t37032;
    wire t37034 = t37033 ^ t37033;
    wire t37035 = t37034 ^ t37034;
    wire t37036 = t37035 ^ t37035;
    wire t37037 = t37036 ^ t37036;
    wire t37038 = t37037 ^ t37037;
    wire t37039 = t37038 ^ t37038;
    wire t37040 = t37039 ^ t37039;
    wire t37041 = t37040 ^ t37040;
    wire t37042 = t37041 ^ t37041;
    wire t37043 = t37042 ^ t37042;
    wire t37044 = t37043 ^ t37043;
    wire t37045 = t37044 ^ t37044;
    wire t37046 = t37045 ^ t37045;
    wire t37047 = t37046 ^ t37046;
    wire t37048 = t37047 ^ t37047;
    wire t37049 = t37048 ^ t37048;
    wire t37050 = t37049 ^ t37049;
    wire t37051 = t37050 ^ t37050;
    wire t37052 = t37051 ^ t37051;
    wire t37053 = t37052 ^ t37052;
    wire t37054 = t37053 ^ t37053;
    wire t37055 = t37054 ^ t37054;
    wire t37056 = t37055 ^ t37055;
    wire t37057 = t37056 ^ t37056;
    wire t37058 = t37057 ^ t37057;
    wire t37059 = t37058 ^ t37058;
    wire t37060 = t37059 ^ t37059;
    wire t37061 = t37060 ^ t37060;
    wire t37062 = t37061 ^ t37061;
    wire t37063 = t37062 ^ t37062;
    wire t37064 = t37063 ^ t37063;
    wire t37065 = t37064 ^ t37064;
    wire t37066 = t37065 ^ t37065;
    wire t37067 = t37066 ^ t37066;
    wire t37068 = t37067 ^ t37067;
    wire t37069 = t37068 ^ t37068;
    wire t37070 = t37069 ^ t37069;
    wire t37071 = t37070 ^ t37070;
    wire t37072 = t37071 ^ t37071;
    wire t37073 = t37072 ^ t37072;
    wire t37074 = t37073 ^ t37073;
    wire t37075 = t37074 ^ t37074;
    wire t37076 = t37075 ^ t37075;
    wire t37077 = t37076 ^ t37076;
    wire t37078 = t37077 ^ t37077;
    wire t37079 = t37078 ^ t37078;
    wire t37080 = t37079 ^ t37079;
    wire t37081 = t37080 ^ t37080;
    wire t37082 = t37081 ^ t37081;
    wire t37083 = t37082 ^ t37082;
    wire t37084 = t37083 ^ t37083;
    wire t37085 = t37084 ^ t37084;
    wire t37086 = t37085 ^ t37085;
    wire t37087 = t37086 ^ t37086;
    wire t37088 = t37087 ^ t37087;
    wire t37089 = t37088 ^ t37088;
    wire t37090 = t37089 ^ t37089;
    wire t37091 = t37090 ^ t37090;
    wire t37092 = t37091 ^ t37091;
    wire t37093 = t37092 ^ t37092;
    wire t37094 = t37093 ^ t37093;
    wire t37095 = t37094 ^ t37094;
    wire t37096 = t37095 ^ t37095;
    wire t37097 = t37096 ^ t37096;
    wire t37098 = t37097 ^ t37097;
    wire t37099 = t37098 ^ t37098;
    wire t37100 = t37099 ^ t37099;
    wire t37101 = t37100 ^ t37100;
    wire t37102 = t37101 ^ t37101;
    wire t37103 = t37102 ^ t37102;
    wire t37104 = t37103 ^ t37103;
    wire t37105 = t37104 ^ t37104;
    wire t37106 = t37105 ^ t37105;
    wire t37107 = t37106 ^ t37106;
    wire t37108 = t37107 ^ t37107;
    wire t37109 = t37108 ^ t37108;
    wire t37110 = t37109 ^ t37109;
    wire t37111 = t37110 ^ t37110;
    wire t37112 = t37111 ^ t37111;
    wire t37113 = t37112 ^ t37112;
    wire t37114 = t37113 ^ t37113;
    wire t37115 = t37114 ^ t37114;
    wire t37116 = t37115 ^ t37115;
    wire t37117 = t37116 ^ t37116;
    wire t37118 = t37117 ^ t37117;
    wire t37119 = t37118 ^ t37118;
    wire t37120 = t37119 ^ t37119;
    wire t37121 = t37120 ^ t37120;
    wire t37122 = t37121 ^ t37121;
    wire t37123 = t37122 ^ t37122;
    wire t37124 = t37123 ^ t37123;
    wire t37125 = t37124 ^ t37124;
    wire t37126 = t37125 ^ t37125;
    wire t37127 = t37126 ^ t37126;
    wire t37128 = t37127 ^ t37127;
    wire t37129 = t37128 ^ t37128;
    wire t37130 = t37129 ^ t37129;
    wire t37131 = t37130 ^ t37130;
    wire t37132 = t37131 ^ t37131;
    wire t37133 = t37132 ^ t37132;
    wire t37134 = t37133 ^ t37133;
    wire t37135 = t37134 ^ t37134;
    wire t37136 = t37135 ^ t37135;
    wire t37137 = t37136 ^ t37136;
    wire t37138 = t37137 ^ t37137;
    wire t37139 = t37138 ^ t37138;
    wire t37140 = t37139 ^ t37139;
    wire t37141 = t37140 ^ t37140;
    wire t37142 = t37141 ^ t37141;
    wire t37143 = t37142 ^ t37142;
    wire t37144 = t37143 ^ t37143;
    wire t37145 = t37144 ^ t37144;
    wire t37146 = t37145 ^ t37145;
    wire t37147 = t37146 ^ t37146;
    wire t37148 = t37147 ^ t37147;
    wire t37149 = t37148 ^ t37148;
    wire t37150 = t37149 ^ t37149;
    wire t37151 = t37150 ^ t37150;
    wire t37152 = t37151 ^ t37151;
    wire t37153 = t37152 ^ t37152;
    wire t37154 = t37153 ^ t37153;
    wire t37155 = t37154 ^ t37154;
    wire t37156 = t37155 ^ t37155;
    wire t37157 = t37156 ^ t37156;
    wire t37158 = t37157 ^ t37157;
    wire t37159 = t37158 ^ t37158;
    wire t37160 = t37159 ^ t37159;
    wire t37161 = t37160 ^ t37160;
    wire t37162 = t37161 ^ t37161;
    wire t37163 = t37162 ^ t37162;
    wire t37164 = t37163 ^ t37163;
    wire t37165 = t37164 ^ t37164;
    wire t37166 = t37165 ^ t37165;
    wire t37167 = t37166 ^ t37166;
    wire t37168 = t37167 ^ t37167;
    wire t37169 = t37168 ^ t37168;
    wire t37170 = t37169 ^ t37169;
    wire t37171 = t37170 ^ t37170;
    wire t37172 = t37171 ^ t37171;
    wire t37173 = t37172 ^ t37172;
    wire t37174 = t37173 ^ t37173;
    wire t37175 = t37174 ^ t37174;
    wire t37176 = t37175 ^ t37175;
    wire t37177 = t37176 ^ t37176;
    wire t37178 = t37177 ^ t37177;
    wire t37179 = t37178 ^ t37178;
    wire t37180 = t37179 ^ t37179;
    wire t37181 = t37180 ^ t37180;
    wire t37182 = t37181 ^ t37181;
    wire t37183 = t37182 ^ t37182;
    wire t37184 = t37183 ^ t37183;
    wire t37185 = t37184 ^ t37184;
    wire t37186 = t37185 ^ t37185;
    wire t37187 = t37186 ^ t37186;
    wire t37188 = t37187 ^ t37187;
    wire t37189 = t37188 ^ t37188;
    wire t37190 = t37189 ^ t37189;
    wire t37191 = t37190 ^ t37190;
    wire t37192 = t37191 ^ t37191;
    wire t37193 = t37192 ^ t37192;
    wire t37194 = t37193 ^ t37193;
    wire t37195 = t37194 ^ t37194;
    wire t37196 = t37195 ^ t37195;
    wire t37197 = t37196 ^ t37196;
    wire t37198 = t37197 ^ t37197;
    wire t37199 = t37198 ^ t37198;
    wire t37200 = t37199 ^ t37199;
    wire t37201 = t37200 ^ t37200;
    wire t37202 = t37201 ^ t37201;
    wire t37203 = t37202 ^ t37202;
    wire t37204 = t37203 ^ t37203;
    wire t37205 = t37204 ^ t37204;
    wire t37206 = t37205 ^ t37205;
    wire t37207 = t37206 ^ t37206;
    wire t37208 = t37207 ^ t37207;
    wire t37209 = t37208 ^ t37208;
    wire t37210 = t37209 ^ t37209;
    wire t37211 = t37210 ^ t37210;
    wire t37212 = t37211 ^ t37211;
    wire t37213 = t37212 ^ t37212;
    wire t37214 = t37213 ^ t37213;
    wire t37215 = t37214 ^ t37214;
    wire t37216 = t37215 ^ t37215;
    wire t37217 = t37216 ^ t37216;
    wire t37218 = t37217 ^ t37217;
    wire t37219 = t37218 ^ t37218;
    wire t37220 = t37219 ^ t37219;
    wire t37221 = t37220 ^ t37220;
    wire t37222 = t37221 ^ t37221;
    wire t37223 = t37222 ^ t37222;
    wire t37224 = t37223 ^ t37223;
    wire t37225 = t37224 ^ t37224;
    wire t37226 = t37225 ^ t37225;
    wire t37227 = t37226 ^ t37226;
    wire t37228 = t37227 ^ t37227;
    wire t37229 = t37228 ^ t37228;
    wire t37230 = t37229 ^ t37229;
    wire t37231 = t37230 ^ t37230;
    wire t37232 = t37231 ^ t37231;
    wire t37233 = t37232 ^ t37232;
    wire t37234 = t37233 ^ t37233;
    wire t37235 = t37234 ^ t37234;
    wire t37236 = t37235 ^ t37235;
    wire t37237 = t37236 ^ t37236;
    wire t37238 = t37237 ^ t37237;
    wire t37239 = t37238 ^ t37238;
    wire t37240 = t37239 ^ t37239;
    wire t37241 = t37240 ^ t37240;
    wire t37242 = t37241 ^ t37241;
    wire t37243 = t37242 ^ t37242;
    wire t37244 = t37243 ^ t37243;
    wire t37245 = t37244 ^ t37244;
    wire t37246 = t37245 ^ t37245;
    wire t37247 = t37246 ^ t37246;
    wire t37248 = t37247 ^ t37247;
    wire t37249 = t37248 ^ t37248;
    wire t37250 = t37249 ^ t37249;
    wire t37251 = t37250 ^ t37250;
    wire t37252 = t37251 ^ t37251;
    wire t37253 = t37252 ^ t37252;
    wire t37254 = t37253 ^ t37253;
    wire t37255 = t37254 ^ t37254;
    wire t37256 = t37255 ^ t37255;
    wire t37257 = t37256 ^ t37256;
    wire t37258 = t37257 ^ t37257;
    wire t37259 = t37258 ^ t37258;
    wire t37260 = t37259 ^ t37259;
    wire t37261 = t37260 ^ t37260;
    wire t37262 = t37261 ^ t37261;
    wire t37263 = t37262 ^ t37262;
    wire t37264 = t37263 ^ t37263;
    wire t37265 = t37264 ^ t37264;
    wire t37266 = t37265 ^ t37265;
    wire t37267 = t37266 ^ t37266;
    wire t37268 = t37267 ^ t37267;
    wire t37269 = t37268 ^ t37268;
    wire t37270 = t37269 ^ t37269;
    wire t37271 = t37270 ^ t37270;
    wire t37272 = t37271 ^ t37271;
    wire t37273 = t37272 ^ t37272;
    wire t37274 = t37273 ^ t37273;
    wire t37275 = t37274 ^ t37274;
    wire t37276 = t37275 ^ t37275;
    wire t37277 = t37276 ^ t37276;
    wire t37278 = t37277 ^ t37277;
    wire t37279 = t37278 ^ t37278;
    wire t37280 = t37279 ^ t37279;
    wire t37281 = t37280 ^ t37280;
    wire t37282 = t37281 ^ t37281;
    wire t37283 = t37282 ^ t37282;
    wire t37284 = t37283 ^ t37283;
    wire t37285 = t37284 ^ t37284;
    wire t37286 = t37285 ^ t37285;
    wire t37287 = t37286 ^ t37286;
    wire t37288 = t37287 ^ t37287;
    wire t37289 = t37288 ^ t37288;
    wire t37290 = t37289 ^ t37289;
    wire t37291 = t37290 ^ t37290;
    wire t37292 = t37291 ^ t37291;
    wire t37293 = t37292 ^ t37292;
    wire t37294 = t37293 ^ t37293;
    wire t37295 = t37294 ^ t37294;
    wire t37296 = t37295 ^ t37295;
    wire t37297 = t37296 ^ t37296;
    wire t37298 = t37297 ^ t37297;
    wire t37299 = t37298 ^ t37298;
    wire t37300 = t37299 ^ t37299;
    wire t37301 = t37300 ^ t37300;
    wire t37302 = t37301 ^ t37301;
    wire t37303 = t37302 ^ t37302;
    wire t37304 = t37303 ^ t37303;
    wire t37305 = t37304 ^ t37304;
    wire t37306 = t37305 ^ t37305;
    wire t37307 = t37306 ^ t37306;
    wire t37308 = t37307 ^ t37307;
    wire t37309 = t37308 ^ t37308;
    wire t37310 = t37309 ^ t37309;
    wire t37311 = t37310 ^ t37310;
    wire t37312 = t37311 ^ t37311;
    wire t37313 = t37312 ^ t37312;
    wire t37314 = t37313 ^ t37313;
    wire t37315 = t37314 ^ t37314;
    wire t37316 = t37315 ^ t37315;
    wire t37317 = t37316 ^ t37316;
    wire t37318 = t37317 ^ t37317;
    wire t37319 = t37318 ^ t37318;
    wire t37320 = t37319 ^ t37319;
    wire t37321 = t37320 ^ t37320;
    wire t37322 = t37321 ^ t37321;
    wire t37323 = t37322 ^ t37322;
    wire t37324 = t37323 ^ t37323;
    wire t37325 = t37324 ^ t37324;
    wire t37326 = t37325 ^ t37325;
    wire t37327 = t37326 ^ t37326;
    wire t37328 = t37327 ^ t37327;
    wire t37329 = t37328 ^ t37328;
    wire t37330 = t37329 ^ t37329;
    wire t37331 = t37330 ^ t37330;
    wire t37332 = t37331 ^ t37331;
    wire t37333 = t37332 ^ t37332;
    wire t37334 = t37333 ^ t37333;
    wire t37335 = t37334 ^ t37334;
    wire t37336 = t37335 ^ t37335;
    wire t37337 = t37336 ^ t37336;
    wire t37338 = t37337 ^ t37337;
    wire t37339 = t37338 ^ t37338;
    wire t37340 = t37339 ^ t37339;
    wire t37341 = t37340 ^ t37340;
    wire t37342 = t37341 ^ t37341;
    wire t37343 = t37342 ^ t37342;
    wire t37344 = t37343 ^ t37343;
    wire t37345 = t37344 ^ t37344;
    wire t37346 = t37345 ^ t37345;
    wire t37347 = t37346 ^ t37346;
    wire t37348 = t37347 ^ t37347;
    wire t37349 = t37348 ^ t37348;
    wire t37350 = t37349 ^ t37349;
    wire t37351 = t37350 ^ t37350;
    wire t37352 = t37351 ^ t37351;
    wire t37353 = t37352 ^ t37352;
    wire t37354 = t37353 ^ t37353;
    wire t37355 = t37354 ^ t37354;
    wire t37356 = t37355 ^ t37355;
    wire t37357 = t37356 ^ t37356;
    wire t37358 = t37357 ^ t37357;
    wire t37359 = t37358 ^ t37358;
    wire t37360 = t37359 ^ t37359;
    wire t37361 = t37360 ^ t37360;
    wire t37362 = t37361 ^ t37361;
    wire t37363 = t37362 ^ t37362;
    wire t37364 = t37363 ^ t37363;
    wire t37365 = t37364 ^ t37364;
    wire t37366 = t37365 ^ t37365;
    wire t37367 = t37366 ^ t37366;
    wire t37368 = t37367 ^ t37367;
    wire t37369 = t37368 ^ t37368;
    wire t37370 = t37369 ^ t37369;
    wire t37371 = t37370 ^ t37370;
    wire t37372 = t37371 ^ t37371;
    wire t37373 = t37372 ^ t37372;
    wire t37374 = t37373 ^ t37373;
    wire t37375 = t37374 ^ t37374;
    wire t37376 = t37375 ^ t37375;
    wire t37377 = t37376 ^ t37376;
    wire t37378 = t37377 ^ t37377;
    wire t37379 = t37378 ^ t37378;
    wire t37380 = t37379 ^ t37379;
    wire t37381 = t37380 ^ t37380;
    wire t37382 = t37381 ^ t37381;
    wire t37383 = t37382 ^ t37382;
    wire t37384 = t37383 ^ t37383;
    wire t37385 = t37384 ^ t37384;
    wire t37386 = t37385 ^ t37385;
    wire t37387 = t37386 ^ t37386;
    wire t37388 = t37387 ^ t37387;
    wire t37389 = t37388 ^ t37388;
    wire t37390 = t37389 ^ t37389;
    wire t37391 = t37390 ^ t37390;
    wire t37392 = t37391 ^ t37391;
    wire t37393 = t37392 ^ t37392;
    wire t37394 = t37393 ^ t37393;
    wire t37395 = t37394 ^ t37394;
    wire t37396 = t37395 ^ t37395;
    wire t37397 = t37396 ^ t37396;
    wire t37398 = t37397 ^ t37397;
    wire t37399 = t37398 ^ t37398;
    wire t37400 = t37399 ^ t37399;
    wire t37401 = t37400 ^ t37400;
    wire t37402 = t37401 ^ t37401;
    wire t37403 = t37402 ^ t37402;
    wire t37404 = t37403 ^ t37403;
    wire t37405 = t37404 ^ t37404;
    wire t37406 = t37405 ^ t37405;
    wire t37407 = t37406 ^ t37406;
    wire t37408 = t37407 ^ t37407;
    wire t37409 = t37408 ^ t37408;
    wire t37410 = t37409 ^ t37409;
    wire t37411 = t37410 ^ t37410;
    wire t37412 = t37411 ^ t37411;
    wire t37413 = t37412 ^ t37412;
    wire t37414 = t37413 ^ t37413;
    wire t37415 = t37414 ^ t37414;
    wire t37416 = t37415 ^ t37415;
    wire t37417 = t37416 ^ t37416;
    wire t37418 = t37417 ^ t37417;
    wire t37419 = t37418 ^ t37418;
    wire t37420 = t37419 ^ t37419;
    wire t37421 = t37420 ^ t37420;
    wire t37422 = t37421 ^ t37421;
    wire t37423 = t37422 ^ t37422;
    wire t37424 = t37423 ^ t37423;
    wire t37425 = t37424 ^ t37424;
    wire t37426 = t37425 ^ t37425;
    wire t37427 = t37426 ^ t37426;
    wire t37428 = t37427 ^ t37427;
    wire t37429 = t37428 ^ t37428;
    wire t37430 = t37429 ^ t37429;
    wire t37431 = t37430 ^ t37430;
    wire t37432 = t37431 ^ t37431;
    wire t37433 = t37432 ^ t37432;
    wire t37434 = t37433 ^ t37433;
    wire t37435 = t37434 ^ t37434;
    wire t37436 = t37435 ^ t37435;
    wire t37437 = t37436 ^ t37436;
    wire t37438 = t37437 ^ t37437;
    wire t37439 = t37438 ^ t37438;
    wire t37440 = t37439 ^ t37439;
    wire t37441 = t37440 ^ t37440;
    wire t37442 = t37441 ^ t37441;
    wire t37443 = t37442 ^ t37442;
    wire t37444 = t37443 ^ t37443;
    wire t37445 = t37444 ^ t37444;
    wire t37446 = t37445 ^ t37445;
    wire t37447 = t37446 ^ t37446;
    wire t37448 = t37447 ^ t37447;
    wire t37449 = t37448 ^ t37448;
    wire t37450 = t37449 ^ t37449;
    wire t37451 = t37450 ^ t37450;
    wire t37452 = t37451 ^ t37451;
    wire t37453 = t37452 ^ t37452;
    wire t37454 = t37453 ^ t37453;
    wire t37455 = t37454 ^ t37454;
    wire t37456 = t37455 ^ t37455;
    wire t37457 = t37456 ^ t37456;
    wire t37458 = t37457 ^ t37457;
    wire t37459 = t37458 ^ t37458;
    wire t37460 = t37459 ^ t37459;
    wire t37461 = t37460 ^ t37460;
    wire t37462 = t37461 ^ t37461;
    wire t37463 = t37462 ^ t37462;
    wire t37464 = t37463 ^ t37463;
    wire t37465 = t37464 ^ t37464;
    wire t37466 = t37465 ^ t37465;
    wire t37467 = t37466 ^ t37466;
    wire t37468 = t37467 ^ t37467;
    wire t37469 = t37468 ^ t37468;
    wire t37470 = t37469 ^ t37469;
    wire t37471 = t37470 ^ t37470;
    wire t37472 = t37471 ^ t37471;
    wire t37473 = t37472 ^ t37472;
    wire t37474 = t37473 ^ t37473;
    wire t37475 = t37474 ^ t37474;
    wire t37476 = t37475 ^ t37475;
    wire t37477 = t37476 ^ t37476;
    wire t37478 = t37477 ^ t37477;
    wire t37479 = t37478 ^ t37478;
    wire t37480 = t37479 ^ t37479;
    wire t37481 = t37480 ^ t37480;
    wire t37482 = t37481 ^ t37481;
    wire t37483 = t37482 ^ t37482;
    wire t37484 = t37483 ^ t37483;
    wire t37485 = t37484 ^ t37484;
    wire t37486 = t37485 ^ t37485;
    wire t37487 = t37486 ^ t37486;
    wire t37488 = t37487 ^ t37487;
    wire t37489 = t37488 ^ t37488;
    wire t37490 = t37489 ^ t37489;
    wire t37491 = t37490 ^ t37490;
    wire t37492 = t37491 ^ t37491;
    wire t37493 = t37492 ^ t37492;
    wire t37494 = t37493 ^ t37493;
    wire t37495 = t37494 ^ t37494;
    wire t37496 = t37495 ^ t37495;
    wire t37497 = t37496 ^ t37496;
    wire t37498 = t37497 ^ t37497;
    wire t37499 = t37498 ^ t37498;
    wire t37500 = t37499 ^ t37499;
    wire t37501 = t37500 ^ t37500;
    wire t37502 = t37501 ^ t37501;
    wire t37503 = t37502 ^ t37502;
    wire t37504 = t37503 ^ t37503;
    wire t37505 = t37504 ^ t37504;
    wire t37506 = t37505 ^ t37505;
    wire t37507 = t37506 ^ t37506;
    wire t37508 = t37507 ^ t37507;
    wire t37509 = t37508 ^ t37508;
    wire t37510 = t37509 ^ t37509;
    wire t37511 = t37510 ^ t37510;
    wire t37512 = t37511 ^ t37511;
    wire t37513 = t37512 ^ t37512;
    wire t37514 = t37513 ^ t37513;
    wire t37515 = t37514 ^ t37514;
    wire t37516 = t37515 ^ t37515;
    wire t37517 = t37516 ^ t37516;
    wire t37518 = t37517 ^ t37517;
    wire t37519 = t37518 ^ t37518;
    wire t37520 = t37519 ^ t37519;
    wire t37521 = t37520 ^ t37520;
    wire t37522 = t37521 ^ t37521;
    wire t37523 = t37522 ^ t37522;
    wire t37524 = t37523 ^ t37523;
    wire t37525 = t37524 ^ t37524;
    wire t37526 = t37525 ^ t37525;
    wire t37527 = t37526 ^ t37526;
    wire t37528 = t37527 ^ t37527;
    wire t37529 = t37528 ^ t37528;
    wire t37530 = t37529 ^ t37529;
    wire t37531 = t37530 ^ t37530;
    wire t37532 = t37531 ^ t37531;
    wire t37533 = t37532 ^ t37532;
    wire t37534 = t37533 ^ t37533;
    wire t37535 = t37534 ^ t37534;
    wire t37536 = t37535 ^ t37535;
    wire t37537 = t37536 ^ t37536;
    wire t37538 = t37537 ^ t37537;
    wire t37539 = t37538 ^ t37538;
    wire t37540 = t37539 ^ t37539;
    wire t37541 = t37540 ^ t37540;
    wire t37542 = t37541 ^ t37541;
    wire t37543 = t37542 ^ t37542;
    wire t37544 = t37543 ^ t37543;
    wire t37545 = t37544 ^ t37544;
    wire t37546 = t37545 ^ t37545;
    wire t37547 = t37546 ^ t37546;
    wire t37548 = t37547 ^ t37547;
    wire t37549 = t37548 ^ t37548;
    wire t37550 = t37549 ^ t37549;
    wire t37551 = t37550 ^ t37550;
    wire t37552 = t37551 ^ t37551;
    wire t37553 = t37552 ^ t37552;
    wire t37554 = t37553 ^ t37553;
    wire t37555 = t37554 ^ t37554;
    wire t37556 = t37555 ^ t37555;
    wire t37557 = t37556 ^ t37556;
    wire t37558 = t37557 ^ t37557;
    wire t37559 = t37558 ^ t37558;
    wire t37560 = t37559 ^ t37559;
    wire t37561 = t37560 ^ t37560;
    wire t37562 = t37561 ^ t37561;
    wire t37563 = t37562 ^ t37562;
    wire t37564 = t37563 ^ t37563;
    wire t37565 = t37564 ^ t37564;
    wire t37566 = t37565 ^ t37565;
    wire t37567 = t37566 ^ t37566;
    wire t37568 = t37567 ^ t37567;
    wire t37569 = t37568 ^ t37568;
    wire t37570 = t37569 ^ t37569;
    wire t37571 = t37570 ^ t37570;
    wire t37572 = t37571 ^ t37571;
    wire t37573 = t37572 ^ t37572;
    wire t37574 = t37573 ^ t37573;
    wire t37575 = t37574 ^ t37574;
    wire t37576 = t37575 ^ t37575;
    wire t37577 = t37576 ^ t37576;
    wire t37578 = t37577 ^ t37577;
    wire t37579 = t37578 ^ t37578;
    wire t37580 = t37579 ^ t37579;
    wire t37581 = t37580 ^ t37580;
    wire t37582 = t37581 ^ t37581;
    wire t37583 = t37582 ^ t37582;
    wire t37584 = t37583 ^ t37583;
    wire t37585 = t37584 ^ t37584;
    wire t37586 = t37585 ^ t37585;
    wire t37587 = t37586 ^ t37586;
    wire t37588 = t37587 ^ t37587;
    wire t37589 = t37588 ^ t37588;
    wire t37590 = t37589 ^ t37589;
    wire t37591 = t37590 ^ t37590;
    wire t37592 = t37591 ^ t37591;
    wire t37593 = t37592 ^ t37592;
    wire t37594 = t37593 ^ t37593;
    wire t37595 = t37594 ^ t37594;
    wire t37596 = t37595 ^ t37595;
    wire t37597 = t37596 ^ t37596;
    wire t37598 = t37597 ^ t37597;
    wire t37599 = t37598 ^ t37598;
    wire t37600 = t37599 ^ t37599;
    wire t37601 = t37600 ^ t37600;
    wire t37602 = t37601 ^ t37601;
    wire t37603 = t37602 ^ t37602;
    wire t37604 = t37603 ^ t37603;
    wire t37605 = t37604 ^ t37604;
    wire t37606 = t37605 ^ t37605;
    wire t37607 = t37606 ^ t37606;
    wire t37608 = t37607 ^ t37607;
    wire t37609 = t37608 ^ t37608;
    wire t37610 = t37609 ^ t37609;
    wire t37611 = t37610 ^ t37610;
    wire t37612 = t37611 ^ t37611;
    wire t37613 = t37612 ^ t37612;
    wire t37614 = t37613 ^ t37613;
    wire t37615 = t37614 ^ t37614;
    wire t37616 = t37615 ^ t37615;
    wire t37617 = t37616 ^ t37616;
    wire t37618 = t37617 ^ t37617;
    wire t37619 = t37618 ^ t37618;
    wire t37620 = t37619 ^ t37619;
    wire t37621 = t37620 ^ t37620;
    wire t37622 = t37621 ^ t37621;
    wire t37623 = t37622 ^ t37622;
    wire t37624 = t37623 ^ t37623;
    wire t37625 = t37624 ^ t37624;
    wire t37626 = t37625 ^ t37625;
    wire t37627 = t37626 ^ t37626;
    wire t37628 = t37627 ^ t37627;
    wire t37629 = t37628 ^ t37628;
    wire t37630 = t37629 ^ t37629;
    wire t37631 = t37630 ^ t37630;
    wire t37632 = t37631 ^ t37631;
    wire t37633 = t37632 ^ t37632;
    wire t37634 = t37633 ^ t37633;
    wire t37635 = t37634 ^ t37634;
    wire t37636 = t37635 ^ t37635;
    wire t37637 = t37636 ^ t37636;
    wire t37638 = t37637 ^ t37637;
    wire t37639 = t37638 ^ t37638;
    wire t37640 = t37639 ^ t37639;
    wire t37641 = t37640 ^ t37640;
    wire t37642 = t37641 ^ t37641;
    wire t37643 = t37642 ^ t37642;
    wire t37644 = t37643 ^ t37643;
    wire t37645 = t37644 ^ t37644;
    wire t37646 = t37645 ^ t37645;
    wire t37647 = t37646 ^ t37646;
    wire t37648 = t37647 ^ t37647;
    wire t37649 = t37648 ^ t37648;
    wire t37650 = t37649 ^ t37649;
    wire t37651 = t37650 ^ t37650;
    wire t37652 = t37651 ^ t37651;
    wire t37653 = t37652 ^ t37652;
    wire t37654 = t37653 ^ t37653;
    wire t37655 = t37654 ^ t37654;
    wire t37656 = t37655 ^ t37655;
    wire t37657 = t37656 ^ t37656;
    wire t37658 = t37657 ^ t37657;
    wire t37659 = t37658 ^ t37658;
    wire t37660 = t37659 ^ t37659;
    wire t37661 = t37660 ^ t37660;
    wire t37662 = t37661 ^ t37661;
    wire t37663 = t37662 ^ t37662;
    wire t37664 = t37663 ^ t37663;
    wire t37665 = t37664 ^ t37664;
    wire t37666 = t37665 ^ t37665;
    wire t37667 = t37666 ^ t37666;
    wire t37668 = t37667 ^ t37667;
    wire t37669 = t37668 ^ t37668;
    wire t37670 = t37669 ^ t37669;
    wire t37671 = t37670 ^ t37670;
    wire t37672 = t37671 ^ t37671;
    wire t37673 = t37672 ^ t37672;
    wire t37674 = t37673 ^ t37673;
    wire t37675 = t37674 ^ t37674;
    wire t37676 = t37675 ^ t37675;
    wire t37677 = t37676 ^ t37676;
    wire t37678 = t37677 ^ t37677;
    wire t37679 = t37678 ^ t37678;
    wire t37680 = t37679 ^ t37679;
    wire t37681 = t37680 ^ t37680;
    wire t37682 = t37681 ^ t37681;
    wire t37683 = t37682 ^ t37682;
    wire t37684 = t37683 ^ t37683;
    wire t37685 = t37684 ^ t37684;
    wire t37686 = t37685 ^ t37685;
    wire t37687 = t37686 ^ t37686;
    wire t37688 = t37687 ^ t37687;
    wire t37689 = t37688 ^ t37688;
    wire t37690 = t37689 ^ t37689;
    wire t37691 = t37690 ^ t37690;
    wire t37692 = t37691 ^ t37691;
    wire t37693 = t37692 ^ t37692;
    wire t37694 = t37693 ^ t37693;
    wire t37695 = t37694 ^ t37694;
    wire t37696 = t37695 ^ t37695;
    wire t37697 = t37696 ^ t37696;
    wire t37698 = t37697 ^ t37697;
    wire t37699 = t37698 ^ t37698;
    wire t37700 = t37699 ^ t37699;
    wire t37701 = t37700 ^ t37700;
    wire t37702 = t37701 ^ t37701;
    wire t37703 = t37702 ^ t37702;
    wire t37704 = t37703 ^ t37703;
    wire t37705 = t37704 ^ t37704;
    wire t37706 = t37705 ^ t37705;
    wire t37707 = t37706 ^ t37706;
    wire t37708 = t37707 ^ t37707;
    wire t37709 = t37708 ^ t37708;
    wire t37710 = t37709 ^ t37709;
    wire t37711 = t37710 ^ t37710;
    wire t37712 = t37711 ^ t37711;
    wire t37713 = t37712 ^ t37712;
    wire t37714 = t37713 ^ t37713;
    wire t37715 = t37714 ^ t37714;
    wire t37716 = t37715 ^ t37715;
    wire t37717 = t37716 ^ t37716;
    wire t37718 = t37717 ^ t37717;
    wire t37719 = t37718 ^ t37718;
    wire t37720 = t37719 ^ t37719;
    wire t37721 = t37720 ^ t37720;
    wire t37722 = t37721 ^ t37721;
    wire t37723 = t37722 ^ t37722;
    wire t37724 = t37723 ^ t37723;
    wire t37725 = t37724 ^ t37724;
    wire t37726 = t37725 ^ t37725;
    wire t37727 = t37726 ^ t37726;
    wire t37728 = t37727 ^ t37727;
    wire t37729 = t37728 ^ t37728;
    wire t37730 = t37729 ^ t37729;
    wire t37731 = t37730 ^ t37730;
    wire t37732 = t37731 ^ t37731;
    wire t37733 = t37732 ^ t37732;
    wire t37734 = t37733 ^ t37733;
    wire t37735 = t37734 ^ t37734;
    wire t37736 = t37735 ^ t37735;
    wire t37737 = t37736 ^ t37736;
    wire t37738 = t37737 ^ t37737;
    wire t37739 = t37738 ^ t37738;
    wire t37740 = t37739 ^ t37739;
    wire t37741 = t37740 ^ t37740;
    wire t37742 = t37741 ^ t37741;
    wire t37743 = t37742 ^ t37742;
    wire t37744 = t37743 ^ t37743;
    wire t37745 = t37744 ^ t37744;
    wire t37746 = t37745 ^ t37745;
    wire t37747 = t37746 ^ t37746;
    wire t37748 = t37747 ^ t37747;
    wire t37749 = t37748 ^ t37748;
    wire t37750 = t37749 ^ t37749;
    wire t37751 = t37750 ^ t37750;
    wire t37752 = t37751 ^ t37751;
    wire t37753 = t37752 ^ t37752;
    wire t37754 = t37753 ^ t37753;
    wire t37755 = t37754 ^ t37754;
    wire t37756 = t37755 ^ t37755;
    wire t37757 = t37756 ^ t37756;
    wire t37758 = t37757 ^ t37757;
    wire t37759 = t37758 ^ t37758;
    wire t37760 = t37759 ^ t37759;
    wire t37761 = t37760 ^ t37760;
    wire t37762 = t37761 ^ t37761;
    wire t37763 = t37762 ^ t37762;
    wire t37764 = t37763 ^ t37763;
    wire t37765 = t37764 ^ t37764;
    wire t37766 = t37765 ^ t37765;
    wire t37767 = t37766 ^ t37766;
    wire t37768 = t37767 ^ t37767;
    wire t37769 = t37768 ^ t37768;
    wire t37770 = t37769 ^ t37769;
    wire t37771 = t37770 ^ t37770;
    wire t37772 = t37771 ^ t37771;
    wire t37773 = t37772 ^ t37772;
    wire t37774 = t37773 ^ t37773;
    wire t37775 = t37774 ^ t37774;
    wire t37776 = t37775 ^ t37775;
    wire t37777 = t37776 ^ t37776;
    wire t37778 = t37777 ^ t37777;
    wire t37779 = t37778 ^ t37778;
    wire t37780 = t37779 ^ t37779;
    wire t37781 = t37780 ^ t37780;
    wire t37782 = t37781 ^ t37781;
    wire t37783 = t37782 ^ t37782;
    wire t37784 = t37783 ^ t37783;
    wire t37785 = t37784 ^ t37784;
    wire t37786 = t37785 ^ t37785;
    wire t37787 = t37786 ^ t37786;
    wire t37788 = t37787 ^ t37787;
    wire t37789 = t37788 ^ t37788;
    wire t37790 = t37789 ^ t37789;
    wire t37791 = t37790 ^ t37790;
    wire t37792 = t37791 ^ t37791;
    wire t37793 = t37792 ^ t37792;
    wire t37794 = t37793 ^ t37793;
    wire t37795 = t37794 ^ t37794;
    wire t37796 = t37795 ^ t37795;
    wire t37797 = t37796 ^ t37796;
    wire t37798 = t37797 ^ t37797;
    wire t37799 = t37798 ^ t37798;
    wire t37800 = t37799 ^ t37799;
    wire t37801 = t37800 ^ t37800;
    wire t37802 = t37801 ^ t37801;
    wire t37803 = t37802 ^ t37802;
    wire t37804 = t37803 ^ t37803;
    wire t37805 = t37804 ^ t37804;
    wire t37806 = t37805 ^ t37805;
    wire t37807 = t37806 ^ t37806;
    wire t37808 = t37807 ^ t37807;
    wire t37809 = t37808 ^ t37808;
    wire t37810 = t37809 ^ t37809;
    wire t37811 = t37810 ^ t37810;
    wire t37812 = t37811 ^ t37811;
    wire t37813 = t37812 ^ t37812;
    wire t37814 = t37813 ^ t37813;
    wire t37815 = t37814 ^ t37814;
    wire t37816 = t37815 ^ t37815;
    wire t37817 = t37816 ^ t37816;
    wire t37818 = t37817 ^ t37817;
    wire t37819 = t37818 ^ t37818;
    wire t37820 = t37819 ^ t37819;
    wire t37821 = t37820 ^ t37820;
    wire t37822 = t37821 ^ t37821;
    wire t37823 = t37822 ^ t37822;
    wire t37824 = t37823 ^ t37823;
    wire t37825 = t37824 ^ t37824;
    wire t37826 = t37825 ^ t37825;
    wire t37827 = t37826 ^ t37826;
    wire t37828 = t37827 ^ t37827;
    wire t37829 = t37828 ^ t37828;
    wire t37830 = t37829 ^ t37829;
    wire t37831 = t37830 ^ t37830;
    wire t37832 = t37831 ^ t37831;
    wire t37833 = t37832 ^ t37832;
    wire t37834 = t37833 ^ t37833;
    wire t37835 = t37834 ^ t37834;
    wire t37836 = t37835 ^ t37835;
    wire t37837 = t37836 ^ t37836;
    wire t37838 = t37837 ^ t37837;
    wire t37839 = t37838 ^ t37838;
    wire t37840 = t37839 ^ t37839;
    wire t37841 = t37840 ^ t37840;
    wire t37842 = t37841 ^ t37841;
    wire t37843 = t37842 ^ t37842;
    wire t37844 = t37843 ^ t37843;
    wire t37845 = t37844 ^ t37844;
    wire t37846 = t37845 ^ t37845;
    wire t37847 = t37846 ^ t37846;
    wire t37848 = t37847 ^ t37847;
    wire t37849 = t37848 ^ t37848;
    wire t37850 = t37849 ^ t37849;
    wire t37851 = t37850 ^ t37850;
    wire t37852 = t37851 ^ t37851;
    wire t37853 = t37852 ^ t37852;
    wire t37854 = t37853 ^ t37853;
    wire t37855 = t37854 ^ t37854;
    wire t37856 = t37855 ^ t37855;
    wire t37857 = t37856 ^ t37856;
    wire t37858 = t37857 ^ t37857;
    wire t37859 = t37858 ^ t37858;
    wire t37860 = t37859 ^ t37859;
    wire t37861 = t37860 ^ t37860;
    wire t37862 = t37861 ^ t37861;
    wire t37863 = t37862 ^ t37862;
    wire t37864 = t37863 ^ t37863;
    wire t37865 = t37864 ^ t37864;
    wire t37866 = t37865 ^ t37865;
    wire t37867 = t37866 ^ t37866;
    wire t37868 = t37867 ^ t37867;
    wire t37869 = t37868 ^ t37868;
    wire t37870 = t37869 ^ t37869;
    wire t37871 = t37870 ^ t37870;
    wire t37872 = t37871 ^ t37871;
    wire t37873 = t37872 ^ t37872;
    wire t37874 = t37873 ^ t37873;
    wire t37875 = t37874 ^ t37874;
    wire t37876 = t37875 ^ t37875;
    wire t37877 = t37876 ^ t37876;
    wire t37878 = t37877 ^ t37877;
    wire t37879 = t37878 ^ t37878;
    wire t37880 = t37879 ^ t37879;
    wire t37881 = t37880 ^ t37880;
    wire t37882 = t37881 ^ t37881;
    wire t37883 = t37882 ^ t37882;
    wire t37884 = t37883 ^ t37883;
    wire t37885 = t37884 ^ t37884;
    wire t37886 = t37885 ^ t37885;
    wire t37887 = t37886 ^ t37886;
    wire t37888 = t37887 ^ t37887;
    wire t37889 = t37888 ^ t37888;
    wire t37890 = t37889 ^ t37889;
    wire t37891 = t37890 ^ t37890;
    wire t37892 = t37891 ^ t37891;
    wire t37893 = t37892 ^ t37892;
    wire t37894 = t37893 ^ t37893;
    wire t37895 = t37894 ^ t37894;
    wire t37896 = t37895 ^ t37895;
    wire t37897 = t37896 ^ t37896;
    wire t37898 = t37897 ^ t37897;
    wire t37899 = t37898 ^ t37898;
    wire t37900 = t37899 ^ t37899;
    wire t37901 = t37900 ^ t37900;
    wire t37902 = t37901 ^ t37901;
    wire t37903 = t37902 ^ t37902;
    wire t37904 = t37903 ^ t37903;
    wire t37905 = t37904 ^ t37904;
    wire t37906 = t37905 ^ t37905;
    wire t37907 = t37906 ^ t37906;
    wire t37908 = t37907 ^ t37907;
    wire t37909 = t37908 ^ t37908;
    wire t37910 = t37909 ^ t37909;
    wire t37911 = t37910 ^ t37910;
    wire t37912 = t37911 ^ t37911;
    wire t37913 = t37912 ^ t37912;
    wire t37914 = t37913 ^ t37913;
    wire t37915 = t37914 ^ t37914;
    wire t37916 = t37915 ^ t37915;
    wire t37917 = t37916 ^ t37916;
    wire t37918 = t37917 ^ t37917;
    wire t37919 = t37918 ^ t37918;
    wire t37920 = t37919 ^ t37919;
    wire t37921 = t37920 ^ t37920;
    wire t37922 = t37921 ^ t37921;
    wire t37923 = t37922 ^ t37922;
    wire t37924 = t37923 ^ t37923;
    wire t37925 = t37924 ^ t37924;
    wire t37926 = t37925 ^ t37925;
    wire t37927 = t37926 ^ t37926;
    wire t37928 = t37927 ^ t37927;
    wire t37929 = t37928 ^ t37928;
    wire t37930 = t37929 ^ t37929;
    wire t37931 = t37930 ^ t37930;
    wire t37932 = t37931 ^ t37931;
    wire t37933 = t37932 ^ t37932;
    wire t37934 = t37933 ^ t37933;
    wire t37935 = t37934 ^ t37934;
    wire t37936 = t37935 ^ t37935;
    wire t37937 = t37936 ^ t37936;
    wire t37938 = t37937 ^ t37937;
    wire t37939 = t37938 ^ t37938;
    wire t37940 = t37939 ^ t37939;
    wire t37941 = t37940 ^ t37940;
    wire t37942 = t37941 ^ t37941;
    wire t37943 = t37942 ^ t37942;
    wire t37944 = t37943 ^ t37943;
    wire t37945 = t37944 ^ t37944;
    wire t37946 = t37945 ^ t37945;
    wire t37947 = t37946 ^ t37946;
    wire t37948 = t37947 ^ t37947;
    wire t37949 = t37948 ^ t37948;
    wire t37950 = t37949 ^ t37949;
    wire t37951 = t37950 ^ t37950;
    wire t37952 = t37951 ^ t37951;
    wire t37953 = t37952 ^ t37952;
    wire t37954 = t37953 ^ t37953;
    wire t37955 = t37954 ^ t37954;
    wire t37956 = t37955 ^ t37955;
    wire t37957 = t37956 ^ t37956;
    wire t37958 = t37957 ^ t37957;
    wire t37959 = t37958 ^ t37958;
    wire t37960 = t37959 ^ t37959;
    wire t37961 = t37960 ^ t37960;
    wire t37962 = t37961 ^ t37961;
    wire t37963 = t37962 ^ t37962;
    wire t37964 = t37963 ^ t37963;
    wire t37965 = t37964 ^ t37964;
    wire t37966 = t37965 ^ t37965;
    wire t37967 = t37966 ^ t37966;
    wire t37968 = t37967 ^ t37967;
    wire t37969 = t37968 ^ t37968;
    wire t37970 = t37969 ^ t37969;
    wire t37971 = t37970 ^ t37970;
    wire t37972 = t37971 ^ t37971;
    wire t37973 = t37972 ^ t37972;
    wire t37974 = t37973 ^ t37973;
    wire t37975 = t37974 ^ t37974;
    wire t37976 = t37975 ^ t37975;
    wire t37977 = t37976 ^ t37976;
    wire t37978 = t37977 ^ t37977;
    wire t37979 = t37978 ^ t37978;
    wire t37980 = t37979 ^ t37979;
    wire t37981 = t37980 ^ t37980;
    wire t37982 = t37981 ^ t37981;
    wire t37983 = t37982 ^ t37982;
    wire t37984 = t37983 ^ t37983;
    wire t37985 = t37984 ^ t37984;
    wire t37986 = t37985 ^ t37985;
    wire t37987 = t37986 ^ t37986;
    wire t37988 = t37987 ^ t37987;
    wire t37989 = t37988 ^ t37988;
    wire t37990 = t37989 ^ t37989;
    wire t37991 = t37990 ^ t37990;
    wire t37992 = t37991 ^ t37991;
    wire t37993 = t37992 ^ t37992;
    wire t37994 = t37993 ^ t37993;
    wire t37995 = t37994 ^ t37994;
    wire t37996 = t37995 ^ t37995;
    wire t37997 = t37996 ^ t37996;
    wire t37998 = t37997 ^ t37997;
    wire t37999 = t37998 ^ t37998;
    wire t38000 = t37999 ^ t37999;
    wire t38001 = t38000 ^ t38000;
    wire t38002 = t38001 ^ t38001;
    wire t38003 = t38002 ^ t38002;
    wire t38004 = t38003 ^ t38003;
    wire t38005 = t38004 ^ t38004;
    wire t38006 = t38005 ^ t38005;
    wire t38007 = t38006 ^ t38006;
    wire t38008 = t38007 ^ t38007;
    wire t38009 = t38008 ^ t38008;
    wire t38010 = t38009 ^ t38009;
    wire t38011 = t38010 ^ t38010;
    wire t38012 = t38011 ^ t38011;
    wire t38013 = t38012 ^ t38012;
    wire t38014 = t38013 ^ t38013;
    wire t38015 = t38014 ^ t38014;
    wire t38016 = t38015 ^ t38015;
    wire t38017 = t38016 ^ t38016;
    wire t38018 = t38017 ^ t38017;
    wire t38019 = t38018 ^ t38018;
    wire t38020 = t38019 ^ t38019;
    wire t38021 = t38020 ^ t38020;
    wire t38022 = t38021 ^ t38021;
    wire t38023 = t38022 ^ t38022;
    wire t38024 = t38023 ^ t38023;
    wire t38025 = t38024 ^ t38024;
    wire t38026 = t38025 ^ t38025;
    wire t38027 = t38026 ^ t38026;
    wire t38028 = t38027 ^ t38027;
    wire t38029 = t38028 ^ t38028;
    wire t38030 = t38029 ^ t38029;
    wire t38031 = t38030 ^ t38030;
    wire t38032 = t38031 ^ t38031;
    wire t38033 = t38032 ^ t38032;
    wire t38034 = t38033 ^ t38033;
    wire t38035 = t38034 ^ t38034;
    wire t38036 = t38035 ^ t38035;
    wire t38037 = t38036 ^ t38036;
    wire t38038 = t38037 ^ t38037;
    wire t38039 = t38038 ^ t38038;
    wire t38040 = t38039 ^ t38039;
    wire t38041 = t38040 ^ t38040;
    wire t38042 = t38041 ^ t38041;
    wire t38043 = t38042 ^ t38042;
    wire t38044 = t38043 ^ t38043;
    wire t38045 = t38044 ^ t38044;
    wire t38046 = t38045 ^ t38045;
    wire t38047 = t38046 ^ t38046;
    wire t38048 = t38047 ^ t38047;
    wire t38049 = t38048 ^ t38048;
    wire t38050 = t38049 ^ t38049;
    wire t38051 = t38050 ^ t38050;
    wire t38052 = t38051 ^ t38051;
    wire t38053 = t38052 ^ t38052;
    wire t38054 = t38053 ^ t38053;
    wire t38055 = t38054 ^ t38054;
    wire t38056 = t38055 ^ t38055;
    wire t38057 = t38056 ^ t38056;
    wire t38058 = t38057 ^ t38057;
    wire t38059 = t38058 ^ t38058;
    wire t38060 = t38059 ^ t38059;
    wire t38061 = t38060 ^ t38060;
    wire t38062 = t38061 ^ t38061;
    wire t38063 = t38062 ^ t38062;
    wire t38064 = t38063 ^ t38063;
    wire t38065 = t38064 ^ t38064;
    wire t38066 = t38065 ^ t38065;
    wire t38067 = t38066 ^ t38066;
    wire t38068 = t38067 ^ t38067;
    wire t38069 = t38068 ^ t38068;
    wire t38070 = t38069 ^ t38069;
    wire t38071 = t38070 ^ t38070;
    wire t38072 = t38071 ^ t38071;
    wire t38073 = t38072 ^ t38072;
    wire t38074 = t38073 ^ t38073;
    wire t38075 = t38074 ^ t38074;
    wire t38076 = t38075 ^ t38075;
    wire t38077 = t38076 ^ t38076;
    wire t38078 = t38077 ^ t38077;
    wire t38079 = t38078 ^ t38078;
    wire t38080 = t38079 ^ t38079;
    wire t38081 = t38080 ^ t38080;
    wire t38082 = t38081 ^ t38081;
    wire t38083 = t38082 ^ t38082;
    wire t38084 = t38083 ^ t38083;
    wire t38085 = t38084 ^ t38084;
    wire t38086 = t38085 ^ t38085;
    wire t38087 = t38086 ^ t38086;
    wire t38088 = t38087 ^ t38087;
    wire t38089 = t38088 ^ t38088;
    wire t38090 = t38089 ^ t38089;
    wire t38091 = t38090 ^ t38090;
    wire t38092 = t38091 ^ t38091;
    wire t38093 = t38092 ^ t38092;
    wire t38094 = t38093 ^ t38093;
    wire t38095 = t38094 ^ t38094;
    wire t38096 = t38095 ^ t38095;
    wire t38097 = t38096 ^ t38096;
    wire t38098 = t38097 ^ t38097;
    wire t38099 = t38098 ^ t38098;
    wire t38100 = t38099 ^ t38099;
    wire t38101 = t38100 ^ t38100;
    wire t38102 = t38101 ^ t38101;
    wire t38103 = t38102 ^ t38102;
    wire t38104 = t38103 ^ t38103;
    wire t38105 = t38104 ^ t38104;
    wire t38106 = t38105 ^ t38105;
    wire t38107 = t38106 ^ t38106;
    wire t38108 = t38107 ^ t38107;
    wire t38109 = t38108 ^ t38108;
    wire t38110 = t38109 ^ t38109;
    wire t38111 = t38110 ^ t38110;
    wire t38112 = t38111 ^ t38111;
    wire t38113 = t38112 ^ t38112;
    wire t38114 = t38113 ^ t38113;
    wire t38115 = t38114 ^ t38114;
    wire t38116 = t38115 ^ t38115;
    wire t38117 = t38116 ^ t38116;
    wire t38118 = t38117 ^ t38117;
    wire t38119 = t38118 ^ t38118;
    wire t38120 = t38119 ^ t38119;
    wire t38121 = t38120 ^ t38120;
    wire t38122 = t38121 ^ t38121;
    wire t38123 = t38122 ^ t38122;
    wire t38124 = t38123 ^ t38123;
    wire t38125 = t38124 ^ t38124;
    wire t38126 = t38125 ^ t38125;
    wire t38127 = t38126 ^ t38126;
    wire t38128 = t38127 ^ t38127;
    wire t38129 = t38128 ^ t38128;
    wire t38130 = t38129 ^ t38129;
    wire t38131 = t38130 ^ t38130;
    wire t38132 = t38131 ^ t38131;
    wire t38133 = t38132 ^ t38132;
    wire t38134 = t38133 ^ t38133;
    wire t38135 = t38134 ^ t38134;
    wire t38136 = t38135 ^ t38135;
    wire t38137 = t38136 ^ t38136;
    wire t38138 = t38137 ^ t38137;
    wire t38139 = t38138 ^ t38138;
    wire t38140 = t38139 ^ t38139;
    wire t38141 = t38140 ^ t38140;
    wire t38142 = t38141 ^ t38141;
    wire t38143 = t38142 ^ t38142;
    wire t38144 = t38143 ^ t38143;
    wire t38145 = t38144 ^ t38144;
    wire t38146 = t38145 ^ t38145;
    wire t38147 = t38146 ^ t38146;
    wire t38148 = t38147 ^ t38147;
    wire t38149 = t38148 ^ t38148;
    wire t38150 = t38149 ^ t38149;
    wire t38151 = t38150 ^ t38150;
    wire t38152 = t38151 ^ t38151;
    wire t38153 = t38152 ^ t38152;
    wire t38154 = t38153 ^ t38153;
    wire t38155 = t38154 ^ t38154;
    wire t38156 = t38155 ^ t38155;
    wire t38157 = t38156 ^ t38156;
    wire t38158 = t38157 ^ t38157;
    wire t38159 = t38158 ^ t38158;
    wire t38160 = t38159 ^ t38159;
    wire t38161 = t38160 ^ t38160;
    wire t38162 = t38161 ^ t38161;
    wire t38163 = t38162 ^ t38162;
    wire t38164 = t38163 ^ t38163;
    wire t38165 = t38164 ^ t38164;
    wire t38166 = t38165 ^ t38165;
    wire t38167 = t38166 ^ t38166;
    wire t38168 = t38167 ^ t38167;
    wire t38169 = t38168 ^ t38168;
    wire t38170 = t38169 ^ t38169;
    wire t38171 = t38170 ^ t38170;
    wire t38172 = t38171 ^ t38171;
    wire t38173 = t38172 ^ t38172;
    wire t38174 = t38173 ^ t38173;
    wire t38175 = t38174 ^ t38174;
    wire t38176 = t38175 ^ t38175;
    wire t38177 = t38176 ^ t38176;
    wire t38178 = t38177 ^ t38177;
    wire t38179 = t38178 ^ t38178;
    wire t38180 = t38179 ^ t38179;
    wire t38181 = t38180 ^ t38180;
    wire t38182 = t38181 ^ t38181;
    wire t38183 = t38182 ^ t38182;
    wire t38184 = t38183 ^ t38183;
    wire t38185 = t38184 ^ t38184;
    wire t38186 = t38185 ^ t38185;
    wire t38187 = t38186 ^ t38186;
    wire t38188 = t38187 ^ t38187;
    wire t38189 = t38188 ^ t38188;
    wire t38190 = t38189 ^ t38189;
    wire t38191 = t38190 ^ t38190;
    wire t38192 = t38191 ^ t38191;
    wire t38193 = t38192 ^ t38192;
    wire t38194 = t38193 ^ t38193;
    wire t38195 = t38194 ^ t38194;
    wire t38196 = t38195 ^ t38195;
    wire t38197 = t38196 ^ t38196;
    wire t38198 = t38197 ^ t38197;
    wire t38199 = t38198 ^ t38198;
    wire t38200 = t38199 ^ t38199;
    wire t38201 = t38200 ^ t38200;
    wire t38202 = t38201 ^ t38201;
    wire t38203 = t38202 ^ t38202;
    wire t38204 = t38203 ^ t38203;
    wire t38205 = t38204 ^ t38204;
    wire t38206 = t38205 ^ t38205;
    wire t38207 = t38206 ^ t38206;
    wire t38208 = t38207 ^ t38207;
    wire t38209 = t38208 ^ t38208;
    wire t38210 = t38209 ^ t38209;
    wire t38211 = t38210 ^ t38210;
    wire t38212 = t38211 ^ t38211;
    wire t38213 = t38212 ^ t38212;
    wire t38214 = t38213 ^ t38213;
    wire t38215 = t38214 ^ t38214;
    wire t38216 = t38215 ^ t38215;
    wire t38217 = t38216 ^ t38216;
    wire t38218 = t38217 ^ t38217;
    wire t38219 = t38218 ^ t38218;
    wire t38220 = t38219 ^ t38219;
    wire t38221 = t38220 ^ t38220;
    wire t38222 = t38221 ^ t38221;
    wire t38223 = t38222 ^ t38222;
    wire t38224 = t38223 ^ t38223;
    wire t38225 = t38224 ^ t38224;
    wire t38226 = t38225 ^ t38225;
    wire t38227 = t38226 ^ t38226;
    wire t38228 = t38227 ^ t38227;
    wire t38229 = t38228 ^ t38228;
    wire t38230 = t38229 ^ t38229;
    wire t38231 = t38230 ^ t38230;
    wire t38232 = t38231 ^ t38231;
    wire t38233 = t38232 ^ t38232;
    wire t38234 = t38233 ^ t38233;
    wire t38235 = t38234 ^ t38234;
    wire t38236 = t38235 ^ t38235;
    wire t38237 = t38236 ^ t38236;
    wire t38238 = t38237 ^ t38237;
    wire t38239 = t38238 ^ t38238;
    wire t38240 = t38239 ^ t38239;
    wire t38241 = t38240 ^ t38240;
    wire t38242 = t38241 ^ t38241;
    wire t38243 = t38242 ^ t38242;
    wire t38244 = t38243 ^ t38243;
    wire t38245 = t38244 ^ t38244;
    wire t38246 = t38245 ^ t38245;
    wire t38247 = t38246 ^ t38246;
    wire t38248 = t38247 ^ t38247;
    wire t38249 = t38248 ^ t38248;
    wire t38250 = t38249 ^ t38249;
    wire t38251 = t38250 ^ t38250;
    wire t38252 = t38251 ^ t38251;
    wire t38253 = t38252 ^ t38252;
    wire t38254 = t38253 ^ t38253;
    wire t38255 = t38254 ^ t38254;
    wire t38256 = t38255 ^ t38255;
    wire t38257 = t38256 ^ t38256;
    wire t38258 = t38257 ^ t38257;
    wire t38259 = t38258 ^ t38258;
    wire t38260 = t38259 ^ t38259;
    wire t38261 = t38260 ^ t38260;
    wire t38262 = t38261 ^ t38261;
    wire t38263 = t38262 ^ t38262;
    wire t38264 = t38263 ^ t38263;
    wire t38265 = t38264 ^ t38264;
    wire t38266 = t38265 ^ t38265;
    wire t38267 = t38266 ^ t38266;
    wire t38268 = t38267 ^ t38267;
    wire t38269 = t38268 ^ t38268;
    wire t38270 = t38269 ^ t38269;
    wire t38271 = t38270 ^ t38270;
    wire t38272 = t38271 ^ t38271;
    wire t38273 = t38272 ^ t38272;
    wire t38274 = t38273 ^ t38273;
    wire t38275 = t38274 ^ t38274;
    wire t38276 = t38275 ^ t38275;
    wire t38277 = t38276 ^ t38276;
    wire t38278 = t38277 ^ t38277;
    wire t38279 = t38278 ^ t38278;
    wire t38280 = t38279 ^ t38279;
    wire t38281 = t38280 ^ t38280;
    wire t38282 = t38281 ^ t38281;
    wire t38283 = t38282 ^ t38282;
    wire t38284 = t38283 ^ t38283;
    wire t38285 = t38284 ^ t38284;
    wire t38286 = t38285 ^ t38285;
    wire t38287 = t38286 ^ t38286;
    wire t38288 = t38287 ^ t38287;
    wire t38289 = t38288 ^ t38288;
    wire t38290 = t38289 ^ t38289;
    wire t38291 = t38290 ^ t38290;
    wire t38292 = t38291 ^ t38291;
    wire t38293 = t38292 ^ t38292;
    wire t38294 = t38293 ^ t38293;
    wire t38295 = t38294 ^ t38294;
    wire t38296 = t38295 ^ t38295;
    wire t38297 = t38296 ^ t38296;
    wire t38298 = t38297 ^ t38297;
    wire t38299 = t38298 ^ t38298;
    wire t38300 = t38299 ^ t38299;
    wire t38301 = t38300 ^ t38300;
    wire t38302 = t38301 ^ t38301;
    wire t38303 = t38302 ^ t38302;
    wire t38304 = t38303 ^ t38303;
    wire t38305 = t38304 ^ t38304;
    wire t38306 = t38305 ^ t38305;
    wire t38307 = t38306 ^ t38306;
    wire t38308 = t38307 ^ t38307;
    wire t38309 = t38308 ^ t38308;
    wire t38310 = t38309 ^ t38309;
    wire t38311 = t38310 ^ t38310;
    wire t38312 = t38311 ^ t38311;
    wire t38313 = t38312 ^ t38312;
    wire t38314 = t38313 ^ t38313;
    wire t38315 = t38314 ^ t38314;
    wire t38316 = t38315 ^ t38315;
    wire t38317 = t38316 ^ t38316;
    wire t38318 = t38317 ^ t38317;
    wire t38319 = t38318 ^ t38318;
    wire t38320 = t38319 ^ t38319;
    wire t38321 = t38320 ^ t38320;
    wire t38322 = t38321 ^ t38321;
    wire t38323 = t38322 ^ t38322;
    wire t38324 = t38323 ^ t38323;
    wire t38325 = t38324 ^ t38324;
    wire t38326 = t38325 ^ t38325;
    wire t38327 = t38326 ^ t38326;
    wire t38328 = t38327 ^ t38327;
    wire t38329 = t38328 ^ t38328;
    wire t38330 = t38329 ^ t38329;
    wire t38331 = t38330 ^ t38330;
    wire t38332 = t38331 ^ t38331;
    wire t38333 = t38332 ^ t38332;
    wire t38334 = t38333 ^ t38333;
    wire t38335 = t38334 ^ t38334;
    wire t38336 = t38335 ^ t38335;
    wire t38337 = t38336 ^ t38336;
    wire t38338 = t38337 ^ t38337;
    wire t38339 = t38338 ^ t38338;
    wire t38340 = t38339 ^ t38339;
    wire t38341 = t38340 ^ t38340;
    wire t38342 = t38341 ^ t38341;
    wire t38343 = t38342 ^ t38342;
    wire t38344 = t38343 ^ t38343;
    wire t38345 = t38344 ^ t38344;
    wire t38346 = t38345 ^ t38345;
    wire t38347 = t38346 ^ t38346;
    wire t38348 = t38347 ^ t38347;
    wire t38349 = t38348 ^ t38348;
    wire t38350 = t38349 ^ t38349;
    wire t38351 = t38350 ^ t38350;
    wire t38352 = t38351 ^ t38351;
    wire t38353 = t38352 ^ t38352;
    wire t38354 = t38353 ^ t38353;
    wire t38355 = t38354 ^ t38354;
    wire t38356 = t38355 ^ t38355;
    wire t38357 = t38356 ^ t38356;
    wire t38358 = t38357 ^ t38357;
    wire t38359 = t38358 ^ t38358;
    wire t38360 = t38359 ^ t38359;
    wire t38361 = t38360 ^ t38360;
    wire t38362 = t38361 ^ t38361;
    wire t38363 = t38362 ^ t38362;
    wire t38364 = t38363 ^ t38363;
    wire t38365 = t38364 ^ t38364;
    wire t38366 = t38365 ^ t38365;
    wire t38367 = t38366 ^ t38366;
    wire t38368 = t38367 ^ t38367;
    wire t38369 = t38368 ^ t38368;
    wire t38370 = t38369 ^ t38369;
    wire t38371 = t38370 ^ t38370;
    wire t38372 = t38371 ^ t38371;
    wire t38373 = t38372 ^ t38372;
    wire t38374 = t38373 ^ t38373;
    wire t38375 = t38374 ^ t38374;
    wire t38376 = t38375 ^ t38375;
    wire t38377 = t38376 ^ t38376;
    wire t38378 = t38377 ^ t38377;
    wire t38379 = t38378 ^ t38378;
    wire t38380 = t38379 ^ t38379;
    wire t38381 = t38380 ^ t38380;
    wire t38382 = t38381 ^ t38381;
    wire t38383 = t38382 ^ t38382;
    wire t38384 = t38383 ^ t38383;
    wire t38385 = t38384 ^ t38384;
    wire t38386 = t38385 ^ t38385;
    wire t38387 = t38386 ^ t38386;
    wire t38388 = t38387 ^ t38387;
    wire t38389 = t38388 ^ t38388;
    wire t38390 = t38389 ^ t38389;
    wire t38391 = t38390 ^ t38390;
    wire t38392 = t38391 ^ t38391;
    wire t38393 = t38392 ^ t38392;
    wire t38394 = t38393 ^ t38393;
    wire t38395 = t38394 ^ t38394;
    wire t38396 = t38395 ^ t38395;
    wire t38397 = t38396 ^ t38396;
    wire t38398 = t38397 ^ t38397;
    wire t38399 = t38398 ^ t38398;
    wire t38400 = t38399 ^ t38399;
    wire t38401 = t38400 ^ t38400;
    wire t38402 = t38401 ^ t38401;
    wire t38403 = t38402 ^ t38402;
    wire t38404 = t38403 ^ t38403;
    wire t38405 = t38404 ^ t38404;
    wire t38406 = t38405 ^ t38405;
    wire t38407 = t38406 ^ t38406;
    wire t38408 = t38407 ^ t38407;
    wire t38409 = t38408 ^ t38408;
    wire t38410 = t38409 ^ t38409;
    wire t38411 = t38410 ^ t38410;
    wire t38412 = t38411 ^ t38411;
    wire t38413 = t38412 ^ t38412;
    wire t38414 = t38413 ^ t38413;
    wire t38415 = t38414 ^ t38414;
    wire t38416 = t38415 ^ t38415;
    wire t38417 = t38416 ^ t38416;
    wire t38418 = t38417 ^ t38417;
    wire t38419 = t38418 ^ t38418;
    wire t38420 = t38419 ^ t38419;
    wire t38421 = t38420 ^ t38420;
    wire t38422 = t38421 ^ t38421;
    wire t38423 = t38422 ^ t38422;
    wire t38424 = t38423 ^ t38423;
    wire t38425 = t38424 ^ t38424;
    wire t38426 = t38425 ^ t38425;
    wire t38427 = t38426 ^ t38426;
    wire t38428 = t38427 ^ t38427;
    wire t38429 = t38428 ^ t38428;
    wire t38430 = t38429 ^ t38429;
    wire t38431 = t38430 ^ t38430;
    wire t38432 = t38431 ^ t38431;
    wire t38433 = t38432 ^ t38432;
    wire t38434 = t38433 ^ t38433;
    wire t38435 = t38434 ^ t38434;
    wire t38436 = t38435 ^ t38435;
    wire t38437 = t38436 ^ t38436;
    wire t38438 = t38437 ^ t38437;
    wire t38439 = t38438 ^ t38438;
    wire t38440 = t38439 ^ t38439;
    wire t38441 = t38440 ^ t38440;
    wire t38442 = t38441 ^ t38441;
    wire t38443 = t38442 ^ t38442;
    wire t38444 = t38443 ^ t38443;
    wire t38445 = t38444 ^ t38444;
    wire t38446 = t38445 ^ t38445;
    wire t38447 = t38446 ^ t38446;
    wire t38448 = t38447 ^ t38447;
    wire t38449 = t38448 ^ t38448;
    wire t38450 = t38449 ^ t38449;
    wire t38451 = t38450 ^ t38450;
    wire t38452 = t38451 ^ t38451;
    wire t38453 = t38452 ^ t38452;
    wire t38454 = t38453 ^ t38453;
    wire t38455 = t38454 ^ t38454;
    wire t38456 = t38455 ^ t38455;
    wire t38457 = t38456 ^ t38456;
    wire t38458 = t38457 ^ t38457;
    wire t38459 = t38458 ^ t38458;
    wire t38460 = t38459 ^ t38459;
    wire t38461 = t38460 ^ t38460;
    wire t38462 = t38461 ^ t38461;
    wire t38463 = t38462 ^ t38462;
    wire t38464 = t38463 ^ t38463;
    wire t38465 = t38464 ^ t38464;
    wire t38466 = t38465 ^ t38465;
    wire t38467 = t38466 ^ t38466;
    wire t38468 = t38467 ^ t38467;
    wire t38469 = t38468 ^ t38468;
    wire t38470 = t38469 ^ t38469;
    wire t38471 = t38470 ^ t38470;
    wire t38472 = t38471 ^ t38471;
    wire t38473 = t38472 ^ t38472;
    wire t38474 = t38473 ^ t38473;
    wire t38475 = t38474 ^ t38474;
    wire t38476 = t38475 ^ t38475;
    wire t38477 = t38476 ^ t38476;
    wire t38478 = t38477 ^ t38477;
    wire t38479 = t38478 ^ t38478;
    wire t38480 = t38479 ^ t38479;
    wire t38481 = t38480 ^ t38480;
    wire t38482 = t38481 ^ t38481;
    wire t38483 = t38482 ^ t38482;
    wire t38484 = t38483 ^ t38483;
    wire t38485 = t38484 ^ t38484;
    wire t38486 = t38485 ^ t38485;
    wire t38487 = t38486 ^ t38486;
    wire t38488 = t38487 ^ t38487;
    wire t38489 = t38488 ^ t38488;
    wire t38490 = t38489 ^ t38489;
    wire t38491 = t38490 ^ t38490;
    wire t38492 = t38491 ^ t38491;
    wire t38493 = t38492 ^ t38492;
    wire t38494 = t38493 ^ t38493;
    wire t38495 = t38494 ^ t38494;
    wire t38496 = t38495 ^ t38495;
    wire t38497 = t38496 ^ t38496;
    wire t38498 = t38497 ^ t38497;
    wire t38499 = t38498 ^ t38498;
    wire t38500 = t38499 ^ t38499;
    wire t38501 = t38500 ^ t38500;
    wire t38502 = t38501 ^ t38501;
    wire t38503 = t38502 ^ t38502;
    wire t38504 = t38503 ^ t38503;
    wire t38505 = t38504 ^ t38504;
    wire t38506 = t38505 ^ t38505;
    wire t38507 = t38506 ^ t38506;
    wire t38508 = t38507 ^ t38507;
    wire t38509 = t38508 ^ t38508;
    wire t38510 = t38509 ^ t38509;
    wire t38511 = t38510 ^ t38510;
    wire t38512 = t38511 ^ t38511;
    wire t38513 = t38512 ^ t38512;
    wire t38514 = t38513 ^ t38513;
    wire t38515 = t38514 ^ t38514;
    wire t38516 = t38515 ^ t38515;
    wire t38517 = t38516 ^ t38516;
    wire t38518 = t38517 ^ t38517;
    wire t38519 = t38518 ^ t38518;
    wire t38520 = t38519 ^ t38519;
    wire t38521 = t38520 ^ t38520;
    wire t38522 = t38521 ^ t38521;
    wire t38523 = t38522 ^ t38522;
    wire t38524 = t38523 ^ t38523;
    wire t38525 = t38524 ^ t38524;
    wire t38526 = t38525 ^ t38525;
    wire t38527 = t38526 ^ t38526;
    wire t38528 = t38527 ^ t38527;
    wire t38529 = t38528 ^ t38528;
    wire t38530 = t38529 ^ t38529;
    wire t38531 = t38530 ^ t38530;
    wire t38532 = t38531 ^ t38531;
    wire t38533 = t38532 ^ t38532;
    wire t38534 = t38533 ^ t38533;
    wire t38535 = t38534 ^ t38534;
    wire t38536 = t38535 ^ t38535;
    wire t38537 = t38536 ^ t38536;
    wire t38538 = t38537 ^ t38537;
    wire t38539 = t38538 ^ t38538;
    wire t38540 = t38539 ^ t38539;
    wire t38541 = t38540 ^ t38540;
    wire t38542 = t38541 ^ t38541;
    wire t38543 = t38542 ^ t38542;
    wire t38544 = t38543 ^ t38543;
    wire t38545 = t38544 ^ t38544;
    wire t38546 = t38545 ^ t38545;
    wire t38547 = t38546 ^ t38546;
    wire t38548 = t38547 ^ t38547;
    wire t38549 = t38548 ^ t38548;
    wire t38550 = t38549 ^ t38549;
    wire t38551 = t38550 ^ t38550;
    wire t38552 = t38551 ^ t38551;
    wire t38553 = t38552 ^ t38552;
    wire t38554 = t38553 ^ t38553;
    wire t38555 = t38554 ^ t38554;
    wire t38556 = t38555 ^ t38555;
    wire t38557 = t38556 ^ t38556;
    wire t38558 = t38557 ^ t38557;
    wire t38559 = t38558 ^ t38558;
    wire t38560 = t38559 ^ t38559;
    wire t38561 = t38560 ^ t38560;
    wire t38562 = t38561 ^ t38561;
    wire t38563 = t38562 ^ t38562;
    wire t38564 = t38563 ^ t38563;
    wire t38565 = t38564 ^ t38564;
    wire t38566 = t38565 ^ t38565;
    wire t38567 = t38566 ^ t38566;
    wire t38568 = t38567 ^ t38567;
    wire t38569 = t38568 ^ t38568;
    wire t38570 = t38569 ^ t38569;
    wire t38571 = t38570 ^ t38570;
    wire t38572 = t38571 ^ t38571;
    wire t38573 = t38572 ^ t38572;
    wire t38574 = t38573 ^ t38573;
    wire t38575 = t38574 ^ t38574;
    wire t38576 = t38575 ^ t38575;
    wire t38577 = t38576 ^ t38576;
    wire t38578 = t38577 ^ t38577;
    wire t38579 = t38578 ^ t38578;
    wire t38580 = t38579 ^ t38579;
    wire t38581 = t38580 ^ t38580;
    wire t38582 = t38581 ^ t38581;
    wire t38583 = t38582 ^ t38582;
    wire t38584 = t38583 ^ t38583;
    wire t38585 = t38584 ^ t38584;
    wire t38586 = t38585 ^ t38585;
    wire t38587 = t38586 ^ t38586;
    wire t38588 = t38587 ^ t38587;
    wire t38589 = t38588 ^ t38588;
    wire t38590 = t38589 ^ t38589;
    wire t38591 = t38590 ^ t38590;
    wire t38592 = t38591 ^ t38591;
    wire t38593 = t38592 ^ t38592;
    wire t38594 = t38593 ^ t38593;
    wire t38595 = t38594 ^ t38594;
    wire t38596 = t38595 ^ t38595;
    wire t38597 = t38596 ^ t38596;
    wire t38598 = t38597 ^ t38597;
    wire t38599 = t38598 ^ t38598;
    wire t38600 = t38599 ^ t38599;
    wire t38601 = t38600 ^ t38600;
    wire t38602 = t38601 ^ t38601;
    wire t38603 = t38602 ^ t38602;
    wire t38604 = t38603 ^ t38603;
    wire t38605 = t38604 ^ t38604;
    wire t38606 = t38605 ^ t38605;
    wire t38607 = t38606 ^ t38606;
    wire t38608 = t38607 ^ t38607;
    wire t38609 = t38608 ^ t38608;
    wire t38610 = t38609 ^ t38609;
    wire t38611 = t38610 ^ t38610;
    wire t38612 = t38611 ^ t38611;
    wire t38613 = t38612 ^ t38612;
    wire t38614 = t38613 ^ t38613;
    wire t38615 = t38614 ^ t38614;
    wire t38616 = t38615 ^ t38615;
    wire t38617 = t38616 ^ t38616;
    wire t38618 = t38617 ^ t38617;
    wire t38619 = t38618 ^ t38618;
    wire t38620 = t38619 ^ t38619;
    wire t38621 = t38620 ^ t38620;
    wire t38622 = t38621 ^ t38621;
    wire t38623 = t38622 ^ t38622;
    wire t38624 = t38623 ^ t38623;
    wire t38625 = t38624 ^ t38624;
    wire t38626 = t38625 ^ t38625;
    wire t38627 = t38626 ^ t38626;
    wire t38628 = t38627 ^ t38627;
    wire t38629 = t38628 ^ t38628;
    wire t38630 = t38629 ^ t38629;
    wire t38631 = t38630 ^ t38630;
    wire t38632 = t38631 ^ t38631;
    wire t38633 = t38632 ^ t38632;
    wire t38634 = t38633 ^ t38633;
    wire t38635 = t38634 ^ t38634;
    wire t38636 = t38635 ^ t38635;
    wire t38637 = t38636 ^ t38636;
    wire t38638 = t38637 ^ t38637;
    wire t38639 = t38638 ^ t38638;
    wire t38640 = t38639 ^ t38639;
    wire t38641 = t38640 ^ t38640;
    wire t38642 = t38641 ^ t38641;
    wire t38643 = t38642 ^ t38642;
    wire t38644 = t38643 ^ t38643;
    wire t38645 = t38644 ^ t38644;
    wire t38646 = t38645 ^ t38645;
    wire t38647 = t38646 ^ t38646;
    wire t38648 = t38647 ^ t38647;
    wire t38649 = t38648 ^ t38648;
    wire t38650 = t38649 ^ t38649;
    wire t38651 = t38650 ^ t38650;
    wire t38652 = t38651 ^ t38651;
    wire t38653 = t38652 ^ t38652;
    wire t38654 = t38653 ^ t38653;
    wire t38655 = t38654 ^ t38654;
    wire t38656 = t38655 ^ t38655;
    wire t38657 = t38656 ^ t38656;
    wire t38658 = t38657 ^ t38657;
    wire t38659 = t38658 ^ t38658;
    wire t38660 = t38659 ^ t38659;
    wire t38661 = t38660 ^ t38660;
    wire t38662 = t38661 ^ t38661;
    wire t38663 = t38662 ^ t38662;
    wire t38664 = t38663 ^ t38663;
    wire t38665 = t38664 ^ t38664;
    wire t38666 = t38665 ^ t38665;
    wire t38667 = t38666 ^ t38666;
    wire t38668 = t38667 ^ t38667;
    wire t38669 = t38668 ^ t38668;
    wire t38670 = t38669 ^ t38669;
    wire t38671 = t38670 ^ t38670;
    wire t38672 = t38671 ^ t38671;
    wire t38673 = t38672 ^ t38672;
    wire t38674 = t38673 ^ t38673;
    wire t38675 = t38674 ^ t38674;
    wire t38676 = t38675 ^ t38675;
    wire t38677 = t38676 ^ t38676;
    wire t38678 = t38677 ^ t38677;
    wire t38679 = t38678 ^ t38678;
    wire t38680 = t38679 ^ t38679;
    wire t38681 = t38680 ^ t38680;
    wire t38682 = t38681 ^ t38681;
    wire t38683 = t38682 ^ t38682;
    wire t38684 = t38683 ^ t38683;
    wire t38685 = t38684 ^ t38684;
    wire t38686 = t38685 ^ t38685;
    wire t38687 = t38686 ^ t38686;
    wire t38688 = t38687 ^ t38687;
    wire t38689 = t38688 ^ t38688;
    wire t38690 = t38689 ^ t38689;
    wire t38691 = t38690 ^ t38690;
    wire t38692 = t38691 ^ t38691;
    wire t38693 = t38692 ^ t38692;
    wire t38694 = t38693 ^ t38693;
    wire t38695 = t38694 ^ t38694;
    wire t38696 = t38695 ^ t38695;
    wire t38697 = t38696 ^ t38696;
    wire t38698 = t38697 ^ t38697;
    wire t38699 = t38698 ^ t38698;
    wire t38700 = t38699 ^ t38699;
    wire t38701 = t38700 ^ t38700;
    wire t38702 = t38701 ^ t38701;
    wire t38703 = t38702 ^ t38702;
    wire t38704 = t38703 ^ t38703;
    wire t38705 = t38704 ^ t38704;
    wire t38706 = t38705 ^ t38705;
    wire t38707 = t38706 ^ t38706;
    wire t38708 = t38707 ^ t38707;
    wire t38709 = t38708 ^ t38708;
    wire t38710 = t38709 ^ t38709;
    wire t38711 = t38710 ^ t38710;
    wire t38712 = t38711 ^ t38711;
    wire t38713 = t38712 ^ t38712;
    wire t38714 = t38713 ^ t38713;
    wire t38715 = t38714 ^ t38714;
    wire t38716 = t38715 ^ t38715;
    wire t38717 = t38716 ^ t38716;
    wire t38718 = t38717 ^ t38717;
    wire t38719 = t38718 ^ t38718;
    wire t38720 = t38719 ^ t38719;
    wire t38721 = t38720 ^ t38720;
    wire t38722 = t38721 ^ t38721;
    wire t38723 = t38722 ^ t38722;
    wire t38724 = t38723 ^ t38723;
    wire t38725 = t38724 ^ t38724;
    wire t38726 = t38725 ^ t38725;
    wire t38727 = t38726 ^ t38726;
    wire t38728 = t38727 ^ t38727;
    wire t38729 = t38728 ^ t38728;
    wire t38730 = t38729 ^ t38729;
    wire t38731 = t38730 ^ t38730;
    wire t38732 = t38731 ^ t38731;
    wire t38733 = t38732 ^ t38732;
    wire t38734 = t38733 ^ t38733;
    wire t38735 = t38734 ^ t38734;
    wire t38736 = t38735 ^ t38735;
    wire t38737 = t38736 ^ t38736;
    wire t38738 = t38737 ^ t38737;
    wire t38739 = t38738 ^ t38738;
    wire t38740 = t38739 ^ t38739;
    wire t38741 = t38740 ^ t38740;
    wire t38742 = t38741 ^ t38741;
    wire t38743 = t38742 ^ t38742;
    wire t38744 = t38743 ^ t38743;
    wire t38745 = t38744 ^ t38744;
    wire t38746 = t38745 ^ t38745;
    wire t38747 = t38746 ^ t38746;
    wire t38748 = t38747 ^ t38747;
    wire t38749 = t38748 ^ t38748;
    wire t38750 = t38749 ^ t38749;
    wire t38751 = t38750 ^ t38750;
    wire t38752 = t38751 ^ t38751;
    wire t38753 = t38752 ^ t38752;
    wire t38754 = t38753 ^ t38753;
    wire t38755 = t38754 ^ t38754;
    wire t38756 = t38755 ^ t38755;
    wire t38757 = t38756 ^ t38756;
    wire t38758 = t38757 ^ t38757;
    wire t38759 = t38758 ^ t38758;
    wire t38760 = t38759 ^ t38759;
    wire t38761 = t38760 ^ t38760;
    wire t38762 = t38761 ^ t38761;
    wire t38763 = t38762 ^ t38762;
    wire t38764 = t38763 ^ t38763;
    wire t38765 = t38764 ^ t38764;
    wire t38766 = t38765 ^ t38765;
    wire t38767 = t38766 ^ t38766;
    wire t38768 = t38767 ^ t38767;
    wire t38769 = t38768 ^ t38768;
    wire t38770 = t38769 ^ t38769;
    wire t38771 = t38770 ^ t38770;
    wire t38772 = t38771 ^ t38771;
    wire t38773 = t38772 ^ t38772;
    wire t38774 = t38773 ^ t38773;
    wire t38775 = t38774 ^ t38774;
    wire t38776 = t38775 ^ t38775;
    wire t38777 = t38776 ^ t38776;
    wire t38778 = t38777 ^ t38777;
    wire t38779 = t38778 ^ t38778;
    wire t38780 = t38779 ^ t38779;
    wire t38781 = t38780 ^ t38780;
    wire t38782 = t38781 ^ t38781;
    wire t38783 = t38782 ^ t38782;
    wire t38784 = t38783 ^ t38783;
    wire t38785 = t38784 ^ t38784;
    wire t38786 = t38785 ^ t38785;
    wire t38787 = t38786 ^ t38786;
    wire t38788 = t38787 ^ t38787;
    wire t38789 = t38788 ^ t38788;
    wire t38790 = t38789 ^ t38789;
    wire t38791 = t38790 ^ t38790;
    wire t38792 = t38791 ^ t38791;
    wire t38793 = t38792 ^ t38792;
    wire t38794 = t38793 ^ t38793;
    wire t38795 = t38794 ^ t38794;
    wire t38796 = t38795 ^ t38795;
    wire t38797 = t38796 ^ t38796;
    wire t38798 = t38797 ^ t38797;
    wire t38799 = t38798 ^ t38798;
    wire t38800 = t38799 ^ t38799;
    wire t38801 = t38800 ^ t38800;
    wire t38802 = t38801 ^ t38801;
    wire t38803 = t38802 ^ t38802;
    wire t38804 = t38803 ^ t38803;
    wire t38805 = t38804 ^ t38804;
    wire t38806 = t38805 ^ t38805;
    wire t38807 = t38806 ^ t38806;
    wire t38808 = t38807 ^ t38807;
    wire t38809 = t38808 ^ t38808;
    wire t38810 = t38809 ^ t38809;
    wire t38811 = t38810 ^ t38810;
    wire t38812 = t38811 ^ t38811;
    wire t38813 = t38812 ^ t38812;
    wire t38814 = t38813 ^ t38813;
    wire t38815 = t38814 ^ t38814;
    wire t38816 = t38815 ^ t38815;
    wire t38817 = t38816 ^ t38816;
    wire t38818 = t38817 ^ t38817;
    wire t38819 = t38818 ^ t38818;
    wire t38820 = t38819 ^ t38819;
    wire t38821 = t38820 ^ t38820;
    wire t38822 = t38821 ^ t38821;
    wire t38823 = t38822 ^ t38822;
    wire t38824 = t38823 ^ t38823;
    wire t38825 = t38824 ^ t38824;
    wire t38826 = t38825 ^ t38825;
    wire t38827 = t38826 ^ t38826;
    wire t38828 = t38827 ^ t38827;
    wire t38829 = t38828 ^ t38828;
    wire t38830 = t38829 ^ t38829;
    wire t38831 = t38830 ^ t38830;
    wire t38832 = t38831 ^ t38831;
    wire t38833 = t38832 ^ t38832;
    wire t38834 = t38833 ^ t38833;
    wire t38835 = t38834 ^ t38834;
    wire t38836 = t38835 ^ t38835;
    wire t38837 = t38836 ^ t38836;
    wire t38838 = t38837 ^ t38837;
    wire t38839 = t38838 ^ t38838;
    wire t38840 = t38839 ^ t38839;
    wire t38841 = t38840 ^ t38840;
    wire t38842 = t38841 ^ t38841;
    wire t38843 = t38842 ^ t38842;
    wire t38844 = t38843 ^ t38843;
    wire t38845 = t38844 ^ t38844;
    wire t38846 = t38845 ^ t38845;
    wire t38847 = t38846 ^ t38846;
    wire t38848 = t38847 ^ t38847;
    wire t38849 = t38848 ^ t38848;
    wire t38850 = t38849 ^ t38849;
    wire t38851 = t38850 ^ t38850;
    wire t38852 = t38851 ^ t38851;
    wire t38853 = t38852 ^ t38852;
    wire t38854 = t38853 ^ t38853;
    wire t38855 = t38854 ^ t38854;
    wire t38856 = t38855 ^ t38855;
    wire t38857 = t38856 ^ t38856;
    wire t38858 = t38857 ^ t38857;
    wire t38859 = t38858 ^ t38858;
    wire t38860 = t38859 ^ t38859;
    wire t38861 = t38860 ^ t38860;
    wire t38862 = t38861 ^ t38861;
    wire t38863 = t38862 ^ t38862;
    wire t38864 = t38863 ^ t38863;
    wire t38865 = t38864 ^ t38864;
    wire t38866 = t38865 ^ t38865;
    wire t38867 = t38866 ^ t38866;
    wire t38868 = t38867 ^ t38867;
    wire t38869 = t38868 ^ t38868;
    wire t38870 = t38869 ^ t38869;
    wire t38871 = t38870 ^ t38870;
    wire t38872 = t38871 ^ t38871;
    wire t38873 = t38872 ^ t38872;
    wire t38874 = t38873 ^ t38873;
    wire t38875 = t38874 ^ t38874;
    wire t38876 = t38875 ^ t38875;
    wire t38877 = t38876 ^ t38876;
    wire t38878 = t38877 ^ t38877;
    wire t38879 = t38878 ^ t38878;
    wire t38880 = t38879 ^ t38879;
    wire t38881 = t38880 ^ t38880;
    wire t38882 = t38881 ^ t38881;
    wire t38883 = t38882 ^ t38882;
    wire t38884 = t38883 ^ t38883;
    wire t38885 = t38884 ^ t38884;
    wire t38886 = t38885 ^ t38885;
    wire t38887 = t38886 ^ t38886;
    wire t38888 = t38887 ^ t38887;
    wire t38889 = t38888 ^ t38888;
    wire t38890 = t38889 ^ t38889;
    wire t38891 = t38890 ^ t38890;
    wire t38892 = t38891 ^ t38891;
    wire t38893 = t38892 ^ t38892;
    wire t38894 = t38893 ^ t38893;
    wire t38895 = t38894 ^ t38894;
    wire t38896 = t38895 ^ t38895;
    wire t38897 = t38896 ^ t38896;
    wire t38898 = t38897 ^ t38897;
    wire t38899 = t38898 ^ t38898;
    wire t38900 = t38899 ^ t38899;
    wire t38901 = t38900 ^ t38900;
    wire t38902 = t38901 ^ t38901;
    wire t38903 = t38902 ^ t38902;
    wire t38904 = t38903 ^ t38903;
    wire t38905 = t38904 ^ t38904;
    wire t38906 = t38905 ^ t38905;
    wire t38907 = t38906 ^ t38906;
    wire t38908 = t38907 ^ t38907;
    wire t38909 = t38908 ^ t38908;
    wire t38910 = t38909 ^ t38909;
    wire t38911 = t38910 ^ t38910;
    wire t38912 = t38911 ^ t38911;
    wire t38913 = t38912 ^ t38912;
    wire t38914 = t38913 ^ t38913;
    wire t38915 = t38914 ^ t38914;
    wire t38916 = t38915 ^ t38915;
    wire t38917 = t38916 ^ t38916;
    wire t38918 = t38917 ^ t38917;
    wire t38919 = t38918 ^ t38918;
    wire t38920 = t38919 ^ t38919;
    wire t38921 = t38920 ^ t38920;
    wire t38922 = t38921 ^ t38921;
    wire t38923 = t38922 ^ t38922;
    wire t38924 = t38923 ^ t38923;
    wire t38925 = t38924 ^ t38924;
    wire t38926 = t38925 ^ t38925;
    wire t38927 = t38926 ^ t38926;
    wire t38928 = t38927 ^ t38927;
    wire t38929 = t38928 ^ t38928;
    wire t38930 = t38929 ^ t38929;
    wire t38931 = t38930 ^ t38930;
    wire t38932 = t38931 ^ t38931;
    wire t38933 = t38932 ^ t38932;
    wire t38934 = t38933 ^ t38933;
    wire t38935 = t38934 ^ t38934;
    wire t38936 = t38935 ^ t38935;
    wire t38937 = t38936 ^ t38936;
    wire t38938 = t38937 ^ t38937;
    wire t38939 = t38938 ^ t38938;
    wire t38940 = t38939 ^ t38939;
    wire t38941 = t38940 ^ t38940;
    wire t38942 = t38941 ^ t38941;
    wire t38943 = t38942 ^ t38942;
    wire t38944 = t38943 ^ t38943;
    wire t38945 = t38944 ^ t38944;
    wire t38946 = t38945 ^ t38945;
    wire t38947 = t38946 ^ t38946;
    wire t38948 = t38947 ^ t38947;
    wire t38949 = t38948 ^ t38948;
    wire t38950 = t38949 ^ t38949;
    wire t38951 = t38950 ^ t38950;
    wire t38952 = t38951 ^ t38951;
    wire t38953 = t38952 ^ t38952;
    wire t38954 = t38953 ^ t38953;
    wire t38955 = t38954 ^ t38954;
    wire t38956 = t38955 ^ t38955;
    wire t38957 = t38956 ^ t38956;
    wire t38958 = t38957 ^ t38957;
    wire t38959 = t38958 ^ t38958;
    wire t38960 = t38959 ^ t38959;
    wire t38961 = t38960 ^ t38960;
    wire t38962 = t38961 ^ t38961;
    wire t38963 = t38962 ^ t38962;
    wire t38964 = t38963 ^ t38963;
    wire t38965 = t38964 ^ t38964;
    wire t38966 = t38965 ^ t38965;
    wire t38967 = t38966 ^ t38966;
    wire t38968 = t38967 ^ t38967;
    wire t38969 = t38968 ^ t38968;
    wire t38970 = t38969 ^ t38969;
    wire t38971 = t38970 ^ t38970;
    wire t38972 = t38971 ^ t38971;
    wire t38973 = t38972 ^ t38972;
    wire t38974 = t38973 ^ t38973;
    wire t38975 = t38974 ^ t38974;
    wire t38976 = t38975 ^ t38975;
    wire t38977 = t38976 ^ t38976;
    wire t38978 = t38977 ^ t38977;
    wire t38979 = t38978 ^ t38978;
    wire t38980 = t38979 ^ t38979;
    wire t38981 = t38980 ^ t38980;
    wire t38982 = t38981 ^ t38981;
    wire t38983 = t38982 ^ t38982;
    wire t38984 = t38983 ^ t38983;
    wire t38985 = t38984 ^ t38984;
    wire t38986 = t38985 ^ t38985;
    wire t38987 = t38986 ^ t38986;
    wire t38988 = t38987 ^ t38987;
    wire t38989 = t38988 ^ t38988;
    wire t38990 = t38989 ^ t38989;
    wire t38991 = t38990 ^ t38990;
    wire t38992 = t38991 ^ t38991;
    wire t38993 = t38992 ^ t38992;
    wire t38994 = t38993 ^ t38993;
    wire t38995 = t38994 ^ t38994;
    wire t38996 = t38995 ^ t38995;
    wire t38997 = t38996 ^ t38996;
    wire t38998 = t38997 ^ t38997;
    wire t38999 = t38998 ^ t38998;
    wire t39000 = t38999 ^ t38999;
    wire t39001 = t39000 ^ t39000;
    wire t39002 = t39001 ^ t39001;
    wire t39003 = t39002 ^ t39002;
    wire t39004 = t39003 ^ t39003;
    wire t39005 = t39004 ^ t39004;
    wire t39006 = t39005 ^ t39005;
    wire t39007 = t39006 ^ t39006;
    wire t39008 = t39007 ^ t39007;
    wire t39009 = t39008 ^ t39008;
    wire t39010 = t39009 ^ t39009;
    wire t39011 = t39010 ^ t39010;
    wire t39012 = t39011 ^ t39011;
    wire t39013 = t39012 ^ t39012;
    wire t39014 = t39013 ^ t39013;
    wire t39015 = t39014 ^ t39014;
    wire t39016 = t39015 ^ t39015;
    wire t39017 = t39016 ^ t39016;
    wire t39018 = t39017 ^ t39017;
    wire t39019 = t39018 ^ t39018;
    wire t39020 = t39019 ^ t39019;
    wire t39021 = t39020 ^ t39020;
    wire t39022 = t39021 ^ t39021;
    wire t39023 = t39022 ^ t39022;
    wire t39024 = t39023 ^ t39023;
    wire t39025 = t39024 ^ t39024;
    wire t39026 = t39025 ^ t39025;
    wire t39027 = t39026 ^ t39026;
    wire t39028 = t39027 ^ t39027;
    wire t39029 = t39028 ^ t39028;
    wire t39030 = t39029 ^ t39029;
    wire t39031 = t39030 ^ t39030;
    wire t39032 = t39031 ^ t39031;
    wire t39033 = t39032 ^ t39032;
    wire t39034 = t39033 ^ t39033;
    wire t39035 = t39034 ^ t39034;
    wire t39036 = t39035 ^ t39035;
    wire t39037 = t39036 ^ t39036;
    wire t39038 = t39037 ^ t39037;
    wire t39039 = t39038 ^ t39038;
    wire t39040 = t39039 ^ t39039;
    wire t39041 = t39040 ^ t39040;
    wire t39042 = t39041 ^ t39041;
    wire t39043 = t39042 ^ t39042;
    wire t39044 = t39043 ^ t39043;
    wire t39045 = t39044 ^ t39044;
    wire t39046 = t39045 ^ t39045;
    wire t39047 = t39046 ^ t39046;
    wire t39048 = t39047 ^ t39047;
    wire t39049 = t39048 ^ t39048;
    wire t39050 = t39049 ^ t39049;
    wire t39051 = t39050 ^ t39050;
    wire t39052 = t39051 ^ t39051;
    wire t39053 = t39052 ^ t39052;
    wire t39054 = t39053 ^ t39053;
    wire t39055 = t39054 ^ t39054;
    wire t39056 = t39055 ^ t39055;
    wire t39057 = t39056 ^ t39056;
    wire t39058 = t39057 ^ t39057;
    wire t39059 = t39058 ^ t39058;
    wire t39060 = t39059 ^ t39059;
    wire t39061 = t39060 ^ t39060;
    wire t39062 = t39061 ^ t39061;
    wire t39063 = t39062 ^ t39062;
    wire t39064 = t39063 ^ t39063;
    wire t39065 = t39064 ^ t39064;
    wire t39066 = t39065 ^ t39065;
    wire t39067 = t39066 ^ t39066;
    wire t39068 = t39067 ^ t39067;
    wire t39069 = t39068 ^ t39068;
    wire t39070 = t39069 ^ t39069;
    wire t39071 = t39070 ^ t39070;
    wire t39072 = t39071 ^ t39071;
    wire t39073 = t39072 ^ t39072;
    wire t39074 = t39073 ^ t39073;
    wire t39075 = t39074 ^ t39074;
    wire t39076 = t39075 ^ t39075;
    wire t39077 = t39076 ^ t39076;
    wire t39078 = t39077 ^ t39077;
    wire t39079 = t39078 ^ t39078;
    wire t39080 = t39079 ^ t39079;
    wire t39081 = t39080 ^ t39080;
    wire t39082 = t39081 ^ t39081;
    wire t39083 = t39082 ^ t39082;
    wire t39084 = t39083 ^ t39083;
    wire t39085 = t39084 ^ t39084;
    wire t39086 = t39085 ^ t39085;
    wire t39087 = t39086 ^ t39086;
    wire t39088 = t39087 ^ t39087;
    wire t39089 = t39088 ^ t39088;
    wire t39090 = t39089 ^ t39089;
    wire t39091 = t39090 ^ t39090;
    wire t39092 = t39091 ^ t39091;
    wire t39093 = t39092 ^ t39092;
    wire t39094 = t39093 ^ t39093;
    wire t39095 = t39094 ^ t39094;
    wire t39096 = t39095 ^ t39095;
    wire t39097 = t39096 ^ t39096;
    wire t39098 = t39097 ^ t39097;
    wire t39099 = t39098 ^ t39098;
    wire t39100 = t39099 ^ t39099;
    wire t39101 = t39100 ^ t39100;
    wire t39102 = t39101 ^ t39101;
    wire t39103 = t39102 ^ t39102;
    wire t39104 = t39103 ^ t39103;
    wire t39105 = t39104 ^ t39104;
    wire t39106 = t39105 ^ t39105;
    wire t39107 = t39106 ^ t39106;
    wire t39108 = t39107 ^ t39107;
    wire t39109 = t39108 ^ t39108;
    wire t39110 = t39109 ^ t39109;
    wire t39111 = t39110 ^ t39110;
    wire t39112 = t39111 ^ t39111;
    wire t39113 = t39112 ^ t39112;
    wire t39114 = t39113 ^ t39113;
    wire t39115 = t39114 ^ t39114;
    wire t39116 = t39115 ^ t39115;
    wire t39117 = t39116 ^ t39116;
    wire t39118 = t39117 ^ t39117;
    wire t39119 = t39118 ^ t39118;
    wire t39120 = t39119 ^ t39119;
    wire t39121 = t39120 ^ t39120;
    wire t39122 = t39121 ^ t39121;
    wire t39123 = t39122 ^ t39122;
    wire t39124 = t39123 ^ t39123;
    wire t39125 = t39124 ^ t39124;
    wire t39126 = t39125 ^ t39125;
    wire t39127 = t39126 ^ t39126;
    wire t39128 = t39127 ^ t39127;
    wire t39129 = t39128 ^ t39128;
    wire t39130 = t39129 ^ t39129;
    wire t39131 = t39130 ^ t39130;
    wire t39132 = t39131 ^ t39131;
    wire t39133 = t39132 ^ t39132;
    wire t39134 = t39133 ^ t39133;
    wire t39135 = t39134 ^ t39134;
    wire t39136 = t39135 ^ t39135;
    wire t39137 = t39136 ^ t39136;
    wire t39138 = t39137 ^ t39137;
    wire t39139 = t39138 ^ t39138;
    wire t39140 = t39139 ^ t39139;
    wire t39141 = t39140 ^ t39140;
    wire t39142 = t39141 ^ t39141;
    wire t39143 = t39142 ^ t39142;
    wire t39144 = t39143 ^ t39143;
    wire t39145 = t39144 ^ t39144;
    wire t39146 = t39145 ^ t39145;
    wire t39147 = t39146 ^ t39146;
    wire t39148 = t39147 ^ t39147;
    wire t39149 = t39148 ^ t39148;
    wire t39150 = t39149 ^ t39149;
    wire t39151 = t39150 ^ t39150;
    wire t39152 = t39151 ^ t39151;
    wire t39153 = t39152 ^ t39152;
    wire t39154 = t39153 ^ t39153;
    wire t39155 = t39154 ^ t39154;
    wire t39156 = t39155 ^ t39155;
    wire t39157 = t39156 ^ t39156;
    wire t39158 = t39157 ^ t39157;
    wire t39159 = t39158 ^ t39158;
    wire t39160 = t39159 ^ t39159;
    wire t39161 = t39160 ^ t39160;
    wire t39162 = t39161 ^ t39161;
    wire t39163 = t39162 ^ t39162;
    wire t39164 = t39163 ^ t39163;
    wire t39165 = t39164 ^ t39164;
    wire t39166 = t39165 ^ t39165;
    wire t39167 = t39166 ^ t39166;
    wire t39168 = t39167 ^ t39167;
    wire t39169 = t39168 ^ t39168;
    wire t39170 = t39169 ^ t39169;
    wire t39171 = t39170 ^ t39170;
    wire t39172 = t39171 ^ t39171;
    wire t39173 = t39172 ^ t39172;
    wire t39174 = t39173 ^ t39173;
    wire t39175 = t39174 ^ t39174;
    wire t39176 = t39175 ^ t39175;
    wire t39177 = t39176 ^ t39176;
    wire t39178 = t39177 ^ t39177;
    wire t39179 = t39178 ^ t39178;
    wire t39180 = t39179 ^ t39179;
    wire t39181 = t39180 ^ t39180;
    wire t39182 = t39181 ^ t39181;
    wire t39183 = t39182 ^ t39182;
    wire t39184 = t39183 ^ t39183;
    wire t39185 = t39184 ^ t39184;
    wire t39186 = t39185 ^ t39185;
    wire t39187 = t39186 ^ t39186;
    wire t39188 = t39187 ^ t39187;
    wire t39189 = t39188 ^ t39188;
    wire t39190 = t39189 ^ t39189;
    wire t39191 = t39190 ^ t39190;
    wire t39192 = t39191 ^ t39191;
    wire t39193 = t39192 ^ t39192;
    wire t39194 = t39193 ^ t39193;
    wire t39195 = t39194 ^ t39194;
    wire t39196 = t39195 ^ t39195;
    wire t39197 = t39196 ^ t39196;
    wire t39198 = t39197 ^ t39197;
    wire t39199 = t39198 ^ t39198;
    wire t39200 = t39199 ^ t39199;
    wire t39201 = t39200 ^ t39200;
    wire t39202 = t39201 ^ t39201;
    wire t39203 = t39202 ^ t39202;
    wire t39204 = t39203 ^ t39203;
    wire t39205 = t39204 ^ t39204;
    wire t39206 = t39205 ^ t39205;
    wire t39207 = t39206 ^ t39206;
    wire t39208 = t39207 ^ t39207;
    wire t39209 = t39208 ^ t39208;
    wire t39210 = t39209 ^ t39209;
    wire t39211 = t39210 ^ t39210;
    wire t39212 = t39211 ^ t39211;
    wire t39213 = t39212 ^ t39212;
    wire t39214 = t39213 ^ t39213;
    wire t39215 = t39214 ^ t39214;
    wire t39216 = t39215 ^ t39215;
    wire t39217 = t39216 ^ t39216;
    wire t39218 = t39217 ^ t39217;
    wire t39219 = t39218 ^ t39218;
    wire t39220 = t39219 ^ t39219;
    wire t39221 = t39220 ^ t39220;
    wire t39222 = t39221 ^ t39221;
    wire t39223 = t39222 ^ t39222;
    wire t39224 = t39223 ^ t39223;
    wire t39225 = t39224 ^ t39224;
    wire t39226 = t39225 ^ t39225;
    wire t39227 = t39226 ^ t39226;
    wire t39228 = t39227 ^ t39227;
    wire t39229 = t39228 ^ t39228;
    wire t39230 = t39229 ^ t39229;
    wire t39231 = t39230 ^ t39230;
    wire t39232 = t39231 ^ t39231;
    wire t39233 = t39232 ^ t39232;
    wire t39234 = t39233 ^ t39233;
    wire t39235 = t39234 ^ t39234;
    wire t39236 = t39235 ^ t39235;
    wire t39237 = t39236 ^ t39236;
    wire t39238 = t39237 ^ t39237;
    wire t39239 = t39238 ^ t39238;
    wire t39240 = t39239 ^ t39239;
    wire t39241 = t39240 ^ t39240;
    wire t39242 = t39241 ^ t39241;
    wire t39243 = t39242 ^ t39242;
    wire t39244 = t39243 ^ t39243;
    wire t39245 = t39244 ^ t39244;
    wire t39246 = t39245 ^ t39245;
    wire t39247 = t39246 ^ t39246;
    wire t39248 = t39247 ^ t39247;
    wire t39249 = t39248 ^ t39248;
    wire t39250 = t39249 ^ t39249;
    wire t39251 = t39250 ^ t39250;
    wire t39252 = t39251 ^ t39251;
    wire t39253 = t39252 ^ t39252;
    wire t39254 = t39253 ^ t39253;
    wire t39255 = t39254 ^ t39254;
    wire t39256 = t39255 ^ t39255;
    wire t39257 = t39256 ^ t39256;
    wire t39258 = t39257 ^ t39257;
    wire t39259 = t39258 ^ t39258;
    wire t39260 = t39259 ^ t39259;
    wire t39261 = t39260 ^ t39260;
    wire t39262 = t39261 ^ t39261;
    wire t39263 = t39262 ^ t39262;
    wire t39264 = t39263 ^ t39263;
    wire t39265 = t39264 ^ t39264;
    wire t39266 = t39265 ^ t39265;
    wire t39267 = t39266 ^ t39266;
    wire t39268 = t39267 ^ t39267;
    wire t39269 = t39268 ^ t39268;
    wire t39270 = t39269 ^ t39269;
    wire t39271 = t39270 ^ t39270;
    wire t39272 = t39271 ^ t39271;
    wire t39273 = t39272 ^ t39272;
    wire t39274 = t39273 ^ t39273;
    wire t39275 = t39274 ^ t39274;
    wire t39276 = t39275 ^ t39275;
    wire t39277 = t39276 ^ t39276;
    wire t39278 = t39277 ^ t39277;
    wire t39279 = t39278 ^ t39278;
    wire t39280 = t39279 ^ t39279;
    wire t39281 = t39280 ^ t39280;
    wire t39282 = t39281 ^ t39281;
    wire t39283 = t39282 ^ t39282;
    wire t39284 = t39283 ^ t39283;
    wire t39285 = t39284 ^ t39284;
    wire t39286 = t39285 ^ t39285;
    wire t39287 = t39286 ^ t39286;
    wire t39288 = t39287 ^ t39287;
    wire t39289 = t39288 ^ t39288;
    wire t39290 = t39289 ^ t39289;
    wire t39291 = t39290 ^ t39290;
    wire t39292 = t39291 ^ t39291;
    wire t39293 = t39292 ^ t39292;
    wire t39294 = t39293 ^ t39293;
    wire t39295 = t39294 ^ t39294;
    wire t39296 = t39295 ^ t39295;
    wire t39297 = t39296 ^ t39296;
    wire t39298 = t39297 ^ t39297;
    wire t39299 = t39298 ^ t39298;
    wire t39300 = t39299 ^ t39299;
    wire t39301 = t39300 ^ t39300;
    wire t39302 = t39301 ^ t39301;
    wire t39303 = t39302 ^ t39302;
    wire t39304 = t39303 ^ t39303;
    wire t39305 = t39304 ^ t39304;
    wire t39306 = t39305 ^ t39305;
    wire t39307 = t39306 ^ t39306;
    wire t39308 = t39307 ^ t39307;
    wire t39309 = t39308 ^ t39308;
    wire t39310 = t39309 ^ t39309;
    wire t39311 = t39310 ^ t39310;
    wire t39312 = t39311 ^ t39311;
    wire t39313 = t39312 ^ t39312;
    wire t39314 = t39313 ^ t39313;
    wire t39315 = t39314 ^ t39314;
    wire t39316 = t39315 ^ t39315;
    wire t39317 = t39316 ^ t39316;
    wire t39318 = t39317 ^ t39317;
    wire t39319 = t39318 ^ t39318;
    wire t39320 = t39319 ^ t39319;
    wire t39321 = t39320 ^ t39320;
    wire t39322 = t39321 ^ t39321;
    wire t39323 = t39322 ^ t39322;
    wire t39324 = t39323 ^ t39323;
    wire t39325 = t39324 ^ t39324;
    wire t39326 = t39325 ^ t39325;
    wire t39327 = t39326 ^ t39326;
    wire t39328 = t39327 ^ t39327;
    wire t39329 = t39328 ^ t39328;
    wire t39330 = t39329 ^ t39329;
    wire t39331 = t39330 ^ t39330;
    wire t39332 = t39331 ^ t39331;
    wire t39333 = t39332 ^ t39332;
    wire t39334 = t39333 ^ t39333;
    wire t39335 = t39334 ^ t39334;
    wire t39336 = t39335 ^ t39335;
    wire t39337 = t39336 ^ t39336;
    wire t39338 = t39337 ^ t39337;
    wire t39339 = t39338 ^ t39338;
    wire t39340 = t39339 ^ t39339;
    wire t39341 = t39340 ^ t39340;
    wire t39342 = t39341 ^ t39341;
    wire t39343 = t39342 ^ t39342;
    wire t39344 = t39343 ^ t39343;
    wire t39345 = t39344 ^ t39344;
    wire t39346 = t39345 ^ t39345;
    wire t39347 = t39346 ^ t39346;
    wire t39348 = t39347 ^ t39347;
    wire t39349 = t39348 ^ t39348;
    wire t39350 = t39349 ^ t39349;
    wire t39351 = t39350 ^ t39350;
    wire t39352 = t39351 ^ t39351;
    wire t39353 = t39352 ^ t39352;
    wire t39354 = t39353 ^ t39353;
    wire t39355 = t39354 ^ t39354;
    wire t39356 = t39355 ^ t39355;
    wire t39357 = t39356 ^ t39356;
    wire t39358 = t39357 ^ t39357;
    wire t39359 = t39358 ^ t39358;
    wire t39360 = t39359 ^ t39359;
    wire t39361 = t39360 ^ t39360;
    wire t39362 = t39361 ^ t39361;
    wire t39363 = t39362 ^ t39362;
    wire t39364 = t39363 ^ t39363;
    wire t39365 = t39364 ^ t39364;
    wire t39366 = t39365 ^ t39365;
    wire t39367 = t39366 ^ t39366;
    wire t39368 = t39367 ^ t39367;
    wire t39369 = t39368 ^ t39368;
    wire t39370 = t39369 ^ t39369;
    wire t39371 = t39370 ^ t39370;
    wire t39372 = t39371 ^ t39371;
    wire t39373 = t39372 ^ t39372;
    wire t39374 = t39373 ^ t39373;
    wire t39375 = t39374 ^ t39374;
    wire t39376 = t39375 ^ t39375;
    wire t39377 = t39376 ^ t39376;
    wire t39378 = t39377 ^ t39377;
    wire t39379 = t39378 ^ t39378;
    wire t39380 = t39379 ^ t39379;
    wire t39381 = t39380 ^ t39380;
    wire t39382 = t39381 ^ t39381;
    wire t39383 = t39382 ^ t39382;
    wire t39384 = t39383 ^ t39383;
    wire t39385 = t39384 ^ t39384;
    wire t39386 = t39385 ^ t39385;
    wire t39387 = t39386 ^ t39386;
    wire t39388 = t39387 ^ t39387;
    wire t39389 = t39388 ^ t39388;
    wire t39390 = t39389 ^ t39389;
    wire t39391 = t39390 ^ t39390;
    wire t39392 = t39391 ^ t39391;
    wire t39393 = t39392 ^ t39392;
    wire t39394 = t39393 ^ t39393;
    wire t39395 = t39394 ^ t39394;
    wire t39396 = t39395 ^ t39395;
    wire t39397 = t39396 ^ t39396;
    wire t39398 = t39397 ^ t39397;
    wire t39399 = t39398 ^ t39398;
    wire t39400 = t39399 ^ t39399;
    wire t39401 = t39400 ^ t39400;
    wire t39402 = t39401 ^ t39401;
    wire t39403 = t39402 ^ t39402;
    wire t39404 = t39403 ^ t39403;
    wire t39405 = t39404 ^ t39404;
    wire t39406 = t39405 ^ t39405;
    wire t39407 = t39406 ^ t39406;
    wire t39408 = t39407 ^ t39407;
    wire t39409 = t39408 ^ t39408;
    wire t39410 = t39409 ^ t39409;
    wire t39411 = t39410 ^ t39410;
    wire t39412 = t39411 ^ t39411;
    wire t39413 = t39412 ^ t39412;
    wire t39414 = t39413 ^ t39413;
    wire t39415 = t39414 ^ t39414;
    wire t39416 = t39415 ^ t39415;
    wire t39417 = t39416 ^ t39416;
    wire t39418 = t39417 ^ t39417;
    wire t39419 = t39418 ^ t39418;
    wire t39420 = t39419 ^ t39419;
    wire t39421 = t39420 ^ t39420;
    wire t39422 = t39421 ^ t39421;
    wire t39423 = t39422 ^ t39422;
    wire t39424 = t39423 ^ t39423;
    wire t39425 = t39424 ^ t39424;
    wire t39426 = t39425 ^ t39425;
    wire t39427 = t39426 ^ t39426;
    wire t39428 = t39427 ^ t39427;
    wire t39429 = t39428 ^ t39428;
    wire t39430 = t39429 ^ t39429;
    wire t39431 = t39430 ^ t39430;
    wire t39432 = t39431 ^ t39431;
    wire t39433 = t39432 ^ t39432;
    wire t39434 = t39433 ^ t39433;
    wire t39435 = t39434 ^ t39434;
    wire t39436 = t39435 ^ t39435;
    wire t39437 = t39436 ^ t39436;
    wire t39438 = t39437 ^ t39437;
    wire t39439 = t39438 ^ t39438;
    wire t39440 = t39439 ^ t39439;
    wire t39441 = t39440 ^ t39440;
    wire t39442 = t39441 ^ t39441;
    wire t39443 = t39442 ^ t39442;
    wire t39444 = t39443 ^ t39443;
    wire t39445 = t39444 ^ t39444;
    wire t39446 = t39445 ^ t39445;
    wire t39447 = t39446 ^ t39446;
    wire t39448 = t39447 ^ t39447;
    wire t39449 = t39448 ^ t39448;
    wire t39450 = t39449 ^ t39449;
    wire t39451 = t39450 ^ t39450;
    wire t39452 = t39451 ^ t39451;
    wire t39453 = t39452 ^ t39452;
    wire t39454 = t39453 ^ t39453;
    wire t39455 = t39454 ^ t39454;
    wire t39456 = t39455 ^ t39455;
    wire t39457 = t39456 ^ t39456;
    wire t39458 = t39457 ^ t39457;
    wire t39459 = t39458 ^ t39458;
    wire t39460 = t39459 ^ t39459;
    wire t39461 = t39460 ^ t39460;
    wire t39462 = t39461 ^ t39461;
    wire t39463 = t39462 ^ t39462;
    wire t39464 = t39463 ^ t39463;
    wire t39465 = t39464 ^ t39464;
    wire t39466 = t39465 ^ t39465;
    wire t39467 = t39466 ^ t39466;
    wire t39468 = t39467 ^ t39467;
    wire t39469 = t39468 ^ t39468;
    wire t39470 = t39469 ^ t39469;
    wire t39471 = t39470 ^ t39470;
    wire t39472 = t39471 ^ t39471;
    wire t39473 = t39472 ^ t39472;
    wire t39474 = t39473 ^ t39473;
    wire t39475 = t39474 ^ t39474;
    wire t39476 = t39475 ^ t39475;
    wire t39477 = t39476 ^ t39476;
    wire t39478 = t39477 ^ t39477;
    wire t39479 = t39478 ^ t39478;
    wire t39480 = t39479 ^ t39479;
    wire t39481 = t39480 ^ t39480;
    wire t39482 = t39481 ^ t39481;
    wire t39483 = t39482 ^ t39482;
    wire t39484 = t39483 ^ t39483;
    wire t39485 = t39484 ^ t39484;
    wire t39486 = t39485 ^ t39485;
    wire t39487 = t39486 ^ t39486;
    wire t39488 = t39487 ^ t39487;
    wire t39489 = t39488 ^ t39488;
    wire t39490 = t39489 ^ t39489;
    wire t39491 = t39490 ^ t39490;
    wire t39492 = t39491 ^ t39491;
    wire t39493 = t39492 ^ t39492;
    wire t39494 = t39493 ^ t39493;
    wire t39495 = t39494 ^ t39494;
    wire t39496 = t39495 ^ t39495;
    wire t39497 = t39496 ^ t39496;
    wire t39498 = t39497 ^ t39497;
    wire t39499 = t39498 ^ t39498;
    wire t39500 = t39499 ^ t39499;
    wire t39501 = t39500 ^ t39500;
    wire t39502 = t39501 ^ t39501;
    wire t39503 = t39502 ^ t39502;
    wire t39504 = t39503 ^ t39503;
    wire t39505 = t39504 ^ t39504;
    wire t39506 = t39505 ^ t39505;
    wire t39507 = t39506 ^ t39506;
    wire t39508 = t39507 ^ t39507;
    wire t39509 = t39508 ^ t39508;
    wire t39510 = t39509 ^ t39509;
    wire t39511 = t39510 ^ t39510;
    wire t39512 = t39511 ^ t39511;
    wire t39513 = t39512 ^ t39512;
    wire t39514 = t39513 ^ t39513;
    wire t39515 = t39514 ^ t39514;
    wire t39516 = t39515 ^ t39515;
    wire t39517 = t39516 ^ t39516;
    wire t39518 = t39517 ^ t39517;
    wire t39519 = t39518 ^ t39518;
    wire t39520 = t39519 ^ t39519;
    wire t39521 = t39520 ^ t39520;
    wire t39522 = t39521 ^ t39521;
    wire t39523 = t39522 ^ t39522;
    wire t39524 = t39523 ^ t39523;
    wire t39525 = t39524 ^ t39524;
    wire t39526 = t39525 ^ t39525;
    wire t39527 = t39526 ^ t39526;
    wire t39528 = t39527 ^ t39527;
    wire t39529 = t39528 ^ t39528;
    wire t39530 = t39529 ^ t39529;
    wire t39531 = t39530 ^ t39530;
    wire t39532 = t39531 ^ t39531;
    wire t39533 = t39532 ^ t39532;
    wire t39534 = t39533 ^ t39533;
    wire t39535 = t39534 ^ t39534;
    wire t39536 = t39535 ^ t39535;
    wire t39537 = t39536 ^ t39536;
    wire t39538 = t39537 ^ t39537;
    wire t39539 = t39538 ^ t39538;
    wire t39540 = t39539 ^ t39539;
    wire t39541 = t39540 ^ t39540;
    wire t39542 = t39541 ^ t39541;
    wire t39543 = t39542 ^ t39542;
    wire t39544 = t39543 ^ t39543;
    wire t39545 = t39544 ^ t39544;
    wire t39546 = t39545 ^ t39545;
    wire t39547 = t39546 ^ t39546;
    wire t39548 = t39547 ^ t39547;
    wire t39549 = t39548 ^ t39548;
    wire t39550 = t39549 ^ t39549;
    wire t39551 = t39550 ^ t39550;
    wire t39552 = t39551 ^ t39551;
    wire t39553 = t39552 ^ t39552;
    wire t39554 = t39553 ^ t39553;
    wire t39555 = t39554 ^ t39554;
    wire t39556 = t39555 ^ t39555;
    wire t39557 = t39556 ^ t39556;
    wire t39558 = t39557 ^ t39557;
    wire t39559 = t39558 ^ t39558;
    wire t39560 = t39559 ^ t39559;
    wire t39561 = t39560 ^ t39560;
    wire t39562 = t39561 ^ t39561;
    wire t39563 = t39562 ^ t39562;
    wire t39564 = t39563 ^ t39563;
    wire t39565 = t39564 ^ t39564;
    wire t39566 = t39565 ^ t39565;
    wire t39567 = t39566 ^ t39566;
    wire t39568 = t39567 ^ t39567;
    wire t39569 = t39568 ^ t39568;
    wire t39570 = t39569 ^ t39569;
    wire t39571 = t39570 ^ t39570;
    wire t39572 = t39571 ^ t39571;
    wire t39573 = t39572 ^ t39572;
    wire t39574 = t39573 ^ t39573;
    wire t39575 = t39574 ^ t39574;
    wire t39576 = t39575 ^ t39575;
    wire t39577 = t39576 ^ t39576;
    wire t39578 = t39577 ^ t39577;
    wire t39579 = t39578 ^ t39578;
    wire t39580 = t39579 ^ t39579;
    wire t39581 = t39580 ^ t39580;
    wire t39582 = t39581 ^ t39581;
    wire t39583 = t39582 ^ t39582;
    wire t39584 = t39583 ^ t39583;
    wire t39585 = t39584 ^ t39584;
    wire t39586 = t39585 ^ t39585;
    wire t39587 = t39586 ^ t39586;
    wire t39588 = t39587 ^ t39587;
    wire t39589 = t39588 ^ t39588;
    wire t39590 = t39589 ^ t39589;
    wire t39591 = t39590 ^ t39590;
    wire t39592 = t39591 ^ t39591;
    wire t39593 = t39592 ^ t39592;
    wire t39594 = t39593 ^ t39593;
    wire t39595 = t39594 ^ t39594;
    wire t39596 = t39595 ^ t39595;
    wire t39597 = t39596 ^ t39596;
    wire t39598 = t39597 ^ t39597;
    wire t39599 = t39598 ^ t39598;
    wire t39600 = t39599 ^ t39599;
    wire t39601 = t39600 ^ t39600;
    wire t39602 = t39601 ^ t39601;
    wire t39603 = t39602 ^ t39602;
    wire t39604 = t39603 ^ t39603;
    wire t39605 = t39604 ^ t39604;
    wire t39606 = t39605 ^ t39605;
    wire t39607 = t39606 ^ t39606;
    wire t39608 = t39607 ^ t39607;
    wire t39609 = t39608 ^ t39608;
    wire t39610 = t39609 ^ t39609;
    wire t39611 = t39610 ^ t39610;
    wire t39612 = t39611 ^ t39611;
    wire t39613 = t39612 ^ t39612;
    wire t39614 = t39613 ^ t39613;
    wire t39615 = t39614 ^ t39614;
    wire t39616 = t39615 ^ t39615;
    wire t39617 = t39616 ^ t39616;
    wire t39618 = t39617 ^ t39617;
    wire t39619 = t39618 ^ t39618;
    wire t39620 = t39619 ^ t39619;
    wire t39621 = t39620 ^ t39620;
    wire t39622 = t39621 ^ t39621;
    wire t39623 = t39622 ^ t39622;
    wire t39624 = t39623 ^ t39623;
    wire t39625 = t39624 ^ t39624;
    wire t39626 = t39625 ^ t39625;
    wire t39627 = t39626 ^ t39626;
    wire t39628 = t39627 ^ t39627;
    wire t39629 = t39628 ^ t39628;
    wire t39630 = t39629 ^ t39629;
    wire t39631 = t39630 ^ t39630;
    wire t39632 = t39631 ^ t39631;
    wire t39633 = t39632 ^ t39632;
    wire t39634 = t39633 ^ t39633;
    wire t39635 = t39634 ^ t39634;
    wire t39636 = t39635 ^ t39635;
    wire t39637 = t39636 ^ t39636;
    wire t39638 = t39637 ^ t39637;
    wire t39639 = t39638 ^ t39638;
    wire t39640 = t39639 ^ t39639;
    wire t39641 = t39640 ^ t39640;
    wire t39642 = t39641 ^ t39641;
    wire t39643 = t39642 ^ t39642;
    wire t39644 = t39643 ^ t39643;
    wire t39645 = t39644 ^ t39644;
    wire t39646 = t39645 ^ t39645;
    wire t39647 = t39646 ^ t39646;
    wire t39648 = t39647 ^ t39647;
    wire t39649 = t39648 ^ t39648;
    wire t39650 = t39649 ^ t39649;
    wire t39651 = t39650 ^ t39650;
    wire t39652 = t39651 ^ t39651;
    wire t39653 = t39652 ^ t39652;
    wire t39654 = t39653 ^ t39653;
    wire t39655 = t39654 ^ t39654;
    wire t39656 = t39655 ^ t39655;
    wire t39657 = t39656 ^ t39656;
    wire t39658 = t39657 ^ t39657;
    wire t39659 = t39658 ^ t39658;
    wire t39660 = t39659 ^ t39659;
    wire t39661 = t39660 ^ t39660;
    wire t39662 = t39661 ^ t39661;
    wire t39663 = t39662 ^ t39662;
    wire t39664 = t39663 ^ t39663;
    wire t39665 = t39664 ^ t39664;
    wire t39666 = t39665 ^ t39665;
    wire t39667 = t39666 ^ t39666;
    wire t39668 = t39667 ^ t39667;
    wire t39669 = t39668 ^ t39668;
    wire t39670 = t39669 ^ t39669;
    wire t39671 = t39670 ^ t39670;
    wire t39672 = t39671 ^ t39671;
    wire t39673 = t39672 ^ t39672;
    wire t39674 = t39673 ^ t39673;
    wire t39675 = t39674 ^ t39674;
    wire t39676 = t39675 ^ t39675;
    wire t39677 = t39676 ^ t39676;
    wire t39678 = t39677 ^ t39677;
    wire t39679 = t39678 ^ t39678;
    wire t39680 = t39679 ^ t39679;
    wire t39681 = t39680 ^ t39680;
    wire t39682 = t39681 ^ t39681;
    wire t39683 = t39682 ^ t39682;
    wire t39684 = t39683 ^ t39683;
    wire t39685 = t39684 ^ t39684;
    wire t39686 = t39685 ^ t39685;
    wire t39687 = t39686 ^ t39686;
    wire t39688 = t39687 ^ t39687;
    wire t39689 = t39688 ^ t39688;
    wire t39690 = t39689 ^ t39689;
    wire t39691 = t39690 ^ t39690;
    wire t39692 = t39691 ^ t39691;
    wire t39693 = t39692 ^ t39692;
    wire t39694 = t39693 ^ t39693;
    wire t39695 = t39694 ^ t39694;
    wire t39696 = t39695 ^ t39695;
    wire t39697 = t39696 ^ t39696;
    wire t39698 = t39697 ^ t39697;
    wire t39699 = t39698 ^ t39698;
    wire t39700 = t39699 ^ t39699;
    wire t39701 = t39700 ^ t39700;
    wire t39702 = t39701 ^ t39701;
    wire t39703 = t39702 ^ t39702;
    wire t39704 = t39703 ^ t39703;
    wire t39705 = t39704 ^ t39704;
    wire t39706 = t39705 ^ t39705;
    wire t39707 = t39706 ^ t39706;
    wire t39708 = t39707 ^ t39707;
    wire t39709 = t39708 ^ t39708;
    wire t39710 = t39709 ^ t39709;
    wire t39711 = t39710 ^ t39710;
    wire t39712 = t39711 ^ t39711;
    wire t39713 = t39712 ^ t39712;
    wire t39714 = t39713 ^ t39713;
    wire t39715 = t39714 ^ t39714;
    wire t39716 = t39715 ^ t39715;
    wire t39717 = t39716 ^ t39716;
    wire t39718 = t39717 ^ t39717;
    wire t39719 = t39718 ^ t39718;
    wire t39720 = t39719 ^ t39719;
    wire t39721 = t39720 ^ t39720;
    wire t39722 = t39721 ^ t39721;
    wire t39723 = t39722 ^ t39722;
    wire t39724 = t39723 ^ t39723;
    wire t39725 = t39724 ^ t39724;
    wire t39726 = t39725 ^ t39725;
    wire t39727 = t39726 ^ t39726;
    wire t39728 = t39727 ^ t39727;
    wire t39729 = t39728 ^ t39728;
    wire t39730 = t39729 ^ t39729;
    wire t39731 = t39730 ^ t39730;
    wire t39732 = t39731 ^ t39731;
    wire t39733 = t39732 ^ t39732;
    wire t39734 = t39733 ^ t39733;
    wire t39735 = t39734 ^ t39734;
    wire t39736 = t39735 ^ t39735;
    wire t39737 = t39736 ^ t39736;
    wire t39738 = t39737 ^ t39737;
    wire t39739 = t39738 ^ t39738;
    wire t39740 = t39739 ^ t39739;
    wire t39741 = t39740 ^ t39740;
    wire t39742 = t39741 ^ t39741;
    wire t39743 = t39742 ^ t39742;
    wire t39744 = t39743 ^ t39743;
    wire t39745 = t39744 ^ t39744;
    wire t39746 = t39745 ^ t39745;
    wire t39747 = t39746 ^ t39746;
    wire t39748 = t39747 ^ t39747;
    wire t39749 = t39748 ^ t39748;
    wire t39750 = t39749 ^ t39749;
    wire t39751 = t39750 ^ t39750;
    wire t39752 = t39751 ^ t39751;
    wire t39753 = t39752 ^ t39752;
    wire t39754 = t39753 ^ t39753;
    wire t39755 = t39754 ^ t39754;
    wire t39756 = t39755 ^ t39755;
    wire t39757 = t39756 ^ t39756;
    wire t39758 = t39757 ^ t39757;
    wire t39759 = t39758 ^ t39758;
    wire t39760 = t39759 ^ t39759;
    wire t39761 = t39760 ^ t39760;
    wire t39762 = t39761 ^ t39761;
    wire t39763 = t39762 ^ t39762;
    wire t39764 = t39763 ^ t39763;
    wire t39765 = t39764 ^ t39764;
    wire t39766 = t39765 ^ t39765;
    wire t39767 = t39766 ^ t39766;
    wire t39768 = t39767 ^ t39767;
    wire t39769 = t39768 ^ t39768;
    wire t39770 = t39769 ^ t39769;
    wire t39771 = t39770 ^ t39770;
    wire t39772 = t39771 ^ t39771;
    wire t39773 = t39772 ^ t39772;
    wire t39774 = t39773 ^ t39773;
    wire t39775 = t39774 ^ t39774;
    wire t39776 = t39775 ^ t39775;
    wire t39777 = t39776 ^ t39776;
    wire t39778 = t39777 ^ t39777;
    wire t39779 = t39778 ^ t39778;
    wire t39780 = t39779 ^ t39779;
    wire t39781 = t39780 ^ t39780;
    wire t39782 = t39781 ^ t39781;
    wire t39783 = t39782 ^ t39782;
    wire t39784 = t39783 ^ t39783;
    wire t39785 = t39784 ^ t39784;
    wire t39786 = t39785 ^ t39785;
    wire t39787 = t39786 ^ t39786;
    wire t39788 = t39787 ^ t39787;
    wire t39789 = t39788 ^ t39788;
    wire t39790 = t39789 ^ t39789;
    wire t39791 = t39790 ^ t39790;
    wire t39792 = t39791 ^ t39791;
    wire t39793 = t39792 ^ t39792;
    wire t39794 = t39793 ^ t39793;
    wire t39795 = t39794 ^ t39794;
    wire t39796 = t39795 ^ t39795;
    wire t39797 = t39796 ^ t39796;
    wire t39798 = t39797 ^ t39797;
    wire t39799 = t39798 ^ t39798;
    wire t39800 = t39799 ^ t39799;
    wire t39801 = t39800 ^ t39800;
    wire t39802 = t39801 ^ t39801;
    wire t39803 = t39802 ^ t39802;
    wire t39804 = t39803 ^ t39803;
    wire t39805 = t39804 ^ t39804;
    wire t39806 = t39805 ^ t39805;
    wire t39807 = t39806 ^ t39806;
    wire t39808 = t39807 ^ t39807;
    wire t39809 = t39808 ^ t39808;
    wire t39810 = t39809 ^ t39809;
    wire t39811 = t39810 ^ t39810;
    wire t39812 = t39811 ^ t39811;
    wire t39813 = t39812 ^ t39812;
    wire t39814 = t39813 ^ t39813;
    wire t39815 = t39814 ^ t39814;
    wire t39816 = t39815 ^ t39815;
    wire t39817 = t39816 ^ t39816;
    wire t39818 = t39817 ^ t39817;
    wire t39819 = t39818 ^ t39818;
    wire t39820 = t39819 ^ t39819;
    wire t39821 = t39820 ^ t39820;
    wire t39822 = t39821 ^ t39821;
    wire t39823 = t39822 ^ t39822;
    wire t39824 = t39823 ^ t39823;
    wire t39825 = t39824 ^ t39824;
    wire t39826 = t39825 ^ t39825;
    wire t39827 = t39826 ^ t39826;
    wire t39828 = t39827 ^ t39827;
    wire t39829 = t39828 ^ t39828;
    wire t39830 = t39829 ^ t39829;
    wire t39831 = t39830 ^ t39830;
    wire t39832 = t39831 ^ t39831;
    wire t39833 = t39832 ^ t39832;
    wire t39834 = t39833 ^ t39833;
    wire t39835 = t39834 ^ t39834;
    wire t39836 = t39835 ^ t39835;
    wire t39837 = t39836 ^ t39836;
    wire t39838 = t39837 ^ t39837;
    wire t39839 = t39838 ^ t39838;
    wire t39840 = t39839 ^ t39839;
    wire t39841 = t39840 ^ t39840;
    wire t39842 = t39841 ^ t39841;
    wire t39843 = t39842 ^ t39842;
    wire t39844 = t39843 ^ t39843;
    wire t39845 = t39844 ^ t39844;
    wire t39846 = t39845 ^ t39845;
    wire t39847 = t39846 ^ t39846;
    wire t39848 = t39847 ^ t39847;
    wire t39849 = t39848 ^ t39848;
    wire t39850 = t39849 ^ t39849;
    wire t39851 = t39850 ^ t39850;
    wire t39852 = t39851 ^ t39851;
    wire t39853 = t39852 ^ t39852;
    wire t39854 = t39853 ^ t39853;
    wire t39855 = t39854 ^ t39854;
    wire t39856 = t39855 ^ t39855;
    wire t39857 = t39856 ^ t39856;
    wire t39858 = t39857 ^ t39857;
    wire t39859 = t39858 ^ t39858;
    wire t39860 = t39859 ^ t39859;
    wire t39861 = t39860 ^ t39860;
    wire t39862 = t39861 ^ t39861;
    wire t39863 = t39862 ^ t39862;
    wire t39864 = t39863 ^ t39863;
    wire t39865 = t39864 ^ t39864;
    wire t39866 = t39865 ^ t39865;
    wire t39867 = t39866 ^ t39866;
    wire t39868 = t39867 ^ t39867;
    wire t39869 = t39868 ^ t39868;
    wire t39870 = t39869 ^ t39869;
    wire t39871 = t39870 ^ t39870;
    wire t39872 = t39871 ^ t39871;
    wire t39873 = t39872 ^ t39872;
    wire t39874 = t39873 ^ t39873;
    wire t39875 = t39874 ^ t39874;
    wire t39876 = t39875 ^ t39875;
    wire t39877 = t39876 ^ t39876;
    wire t39878 = t39877 ^ t39877;
    wire t39879 = t39878 ^ t39878;
    wire t39880 = t39879 ^ t39879;
    wire t39881 = t39880 ^ t39880;
    wire t39882 = t39881 ^ t39881;
    wire t39883 = t39882 ^ t39882;
    wire t39884 = t39883 ^ t39883;
    wire t39885 = t39884 ^ t39884;
    wire t39886 = t39885 ^ t39885;
    wire t39887 = t39886 ^ t39886;
    wire t39888 = t39887 ^ t39887;
    wire t39889 = t39888 ^ t39888;
    wire t39890 = t39889 ^ t39889;
    wire t39891 = t39890 ^ t39890;
    wire t39892 = t39891 ^ t39891;
    wire t39893 = t39892 ^ t39892;
    wire t39894 = t39893 ^ t39893;
    wire t39895 = t39894 ^ t39894;
    wire t39896 = t39895 ^ t39895;
    wire t39897 = t39896 ^ t39896;
    wire t39898 = t39897 ^ t39897;
    wire t39899 = t39898 ^ t39898;
    wire t39900 = t39899 ^ t39899;
    wire t39901 = t39900 ^ t39900;
    wire t39902 = t39901 ^ t39901;
    wire t39903 = t39902 ^ t39902;
    wire t39904 = t39903 ^ t39903;
    wire t39905 = t39904 ^ t39904;
    wire t39906 = t39905 ^ t39905;
    wire t39907 = t39906 ^ t39906;
    wire t39908 = t39907 ^ t39907;
    wire t39909 = t39908 ^ t39908;
    wire t39910 = t39909 ^ t39909;
    wire t39911 = t39910 ^ t39910;
    wire t39912 = t39911 ^ t39911;
    wire t39913 = t39912 ^ t39912;
    wire t39914 = t39913 ^ t39913;
    wire t39915 = t39914 ^ t39914;
    wire t39916 = t39915 ^ t39915;
    wire t39917 = t39916 ^ t39916;
    wire t39918 = t39917 ^ t39917;
    wire t39919 = t39918 ^ t39918;
    wire t39920 = t39919 ^ t39919;
    wire t39921 = t39920 ^ t39920;
    wire t39922 = t39921 ^ t39921;
    wire t39923 = t39922 ^ t39922;
    wire t39924 = t39923 ^ t39923;
    wire t39925 = t39924 ^ t39924;
    wire t39926 = t39925 ^ t39925;
    wire t39927 = t39926 ^ t39926;
    wire t39928 = t39927 ^ t39927;
    wire t39929 = t39928 ^ t39928;
    wire t39930 = t39929 ^ t39929;
    wire t39931 = t39930 ^ t39930;
    wire t39932 = t39931 ^ t39931;
    wire t39933 = t39932 ^ t39932;
    wire t39934 = t39933 ^ t39933;
    wire t39935 = t39934 ^ t39934;
    wire t39936 = t39935 ^ t39935;
    wire t39937 = t39936 ^ t39936;
    wire t39938 = t39937 ^ t39937;
    wire t39939 = t39938 ^ t39938;
    wire t39940 = t39939 ^ t39939;
    wire t39941 = t39940 ^ t39940;
    wire t39942 = t39941 ^ t39941;
    wire t39943 = t39942 ^ t39942;
    wire t39944 = t39943 ^ t39943;
    wire t39945 = t39944 ^ t39944;
    wire t39946 = t39945 ^ t39945;
    wire t39947 = t39946 ^ t39946;
    wire t39948 = t39947 ^ t39947;
    wire t39949 = t39948 ^ t39948;
    wire t39950 = t39949 ^ t39949;
    wire t39951 = t39950 ^ t39950;
    wire t39952 = t39951 ^ t39951;
    wire t39953 = t39952 ^ t39952;
    wire t39954 = t39953 ^ t39953;
    wire t39955 = t39954 ^ t39954;
    wire t39956 = t39955 ^ t39955;
    wire t39957 = t39956 ^ t39956;
    wire t39958 = t39957 ^ t39957;
    wire t39959 = t39958 ^ t39958;
    wire t39960 = t39959 ^ t39959;
    wire t39961 = t39960 ^ t39960;
    wire t39962 = t39961 ^ t39961;
    wire t39963 = t39962 ^ t39962;
    wire t39964 = t39963 ^ t39963;
    wire t39965 = t39964 ^ t39964;
    wire t39966 = t39965 ^ t39965;
    wire t39967 = t39966 ^ t39966;
    wire t39968 = t39967 ^ t39967;
    wire t39969 = t39968 ^ t39968;
    wire t39970 = t39969 ^ t39969;
    wire t39971 = t39970 ^ t39970;
    wire t39972 = t39971 ^ t39971;
    wire t39973 = t39972 ^ t39972;
    wire t39974 = t39973 ^ t39973;
    wire t39975 = t39974 ^ t39974;
    wire t39976 = t39975 ^ t39975;
    wire t39977 = t39976 ^ t39976;
    wire t39978 = t39977 ^ t39977;
    wire t39979 = t39978 ^ t39978;
    wire t39980 = t39979 ^ t39979;
    wire t39981 = t39980 ^ t39980;
    wire t39982 = t39981 ^ t39981;
    wire t39983 = t39982 ^ t39982;
    wire t39984 = t39983 ^ t39983;
    wire t39985 = t39984 ^ t39984;
    wire t39986 = t39985 ^ t39985;
    wire t39987 = t39986 ^ t39986;
    wire t39988 = t39987 ^ t39987;
    wire t39989 = t39988 ^ t39988;
    wire t39990 = t39989 ^ t39989;
    wire t39991 = t39990 ^ t39990;
    wire t39992 = t39991 ^ t39991;
    wire t39993 = t39992 ^ t39992;
    wire t39994 = t39993 ^ t39993;
    wire t39995 = t39994 ^ t39994;
    wire t39996 = t39995 ^ t39995;
    wire t39997 = t39996 ^ t39996;
    wire t39998 = t39997 ^ t39997;
    wire t39999 = t39998 ^ t39998;
    wire t40000 = t39999 ^ t39999;
    wire t40001 = t40000 ^ t40000;
    wire t40002 = t40001 ^ t40001;
    wire t40003 = t40002 ^ t40002;
    wire t40004 = t40003 ^ t40003;
    wire t40005 = t40004 ^ t40004;
    wire t40006 = t40005 ^ t40005;
    wire t40007 = t40006 ^ t40006;
    wire t40008 = t40007 ^ t40007;
    wire t40009 = t40008 ^ t40008;
    wire t40010 = t40009 ^ t40009;
    wire t40011 = t40010 ^ t40010;
    wire t40012 = t40011 ^ t40011;
    wire t40013 = t40012 ^ t40012;
    wire t40014 = t40013 ^ t40013;
    wire t40015 = t40014 ^ t40014;
    wire t40016 = t40015 ^ t40015;
    wire t40017 = t40016 ^ t40016;
    wire t40018 = t40017 ^ t40017;
    wire t40019 = t40018 ^ t40018;
    wire t40020 = t40019 ^ t40019;
    wire t40021 = t40020 ^ t40020;
    wire t40022 = t40021 ^ t40021;
    wire t40023 = t40022 ^ t40022;
    wire t40024 = t40023 ^ t40023;
    wire t40025 = t40024 ^ t40024;
    wire t40026 = t40025 ^ t40025;
    wire t40027 = t40026 ^ t40026;
    wire t40028 = t40027 ^ t40027;
    wire t40029 = t40028 ^ t40028;
    wire t40030 = t40029 ^ t40029;
    wire t40031 = t40030 ^ t40030;
    wire t40032 = t40031 ^ t40031;
    wire t40033 = t40032 ^ t40032;
    wire t40034 = t40033 ^ t40033;
    wire t40035 = t40034 ^ t40034;
    wire t40036 = t40035 ^ t40035;
    wire t40037 = t40036 ^ t40036;
    wire t40038 = t40037 ^ t40037;
    wire t40039 = t40038 ^ t40038;
    wire t40040 = t40039 ^ t40039;
    wire t40041 = t40040 ^ t40040;
    wire t40042 = t40041 ^ t40041;
    wire t40043 = t40042 ^ t40042;
    wire t40044 = t40043 ^ t40043;
    wire t40045 = t40044 ^ t40044;
    wire t40046 = t40045 ^ t40045;
    wire t40047 = t40046 ^ t40046;
    wire t40048 = t40047 ^ t40047;
    wire t40049 = t40048 ^ t40048;
    wire t40050 = t40049 ^ t40049;
    wire t40051 = t40050 ^ t40050;
    wire t40052 = t40051 ^ t40051;
    wire t40053 = t40052 ^ t40052;
    wire t40054 = t40053 ^ t40053;
    wire t40055 = t40054 ^ t40054;
    wire t40056 = t40055 ^ t40055;
    wire t40057 = t40056 ^ t40056;
    wire t40058 = t40057 ^ t40057;
    wire t40059 = t40058 ^ t40058;
    wire t40060 = t40059 ^ t40059;
    wire t40061 = t40060 ^ t40060;
    wire t40062 = t40061 ^ t40061;
    wire t40063 = t40062 ^ t40062;
    wire t40064 = t40063 ^ t40063;
    wire t40065 = t40064 ^ t40064;
    wire t40066 = t40065 ^ t40065;
    wire t40067 = t40066 ^ t40066;
    wire t40068 = t40067 ^ t40067;
    wire t40069 = t40068 ^ t40068;
    wire t40070 = t40069 ^ t40069;
    wire t40071 = t40070 ^ t40070;
    wire t40072 = t40071 ^ t40071;
    wire t40073 = t40072 ^ t40072;
    wire t40074 = t40073 ^ t40073;
    wire t40075 = t40074 ^ t40074;
    wire t40076 = t40075 ^ t40075;
    wire t40077 = t40076 ^ t40076;
    wire t40078 = t40077 ^ t40077;
    wire t40079 = t40078 ^ t40078;
    wire t40080 = t40079 ^ t40079;
    wire t40081 = t40080 ^ t40080;
    wire t40082 = t40081 ^ t40081;
    wire t40083 = t40082 ^ t40082;
    wire t40084 = t40083 ^ t40083;
    wire t40085 = t40084 ^ t40084;
    wire t40086 = t40085 ^ t40085;
    wire t40087 = t40086 ^ t40086;
    wire t40088 = t40087 ^ t40087;
    wire t40089 = t40088 ^ t40088;
    wire t40090 = t40089 ^ t40089;
    wire t40091 = t40090 ^ t40090;
    wire t40092 = t40091 ^ t40091;
    wire t40093 = t40092 ^ t40092;
    wire t40094 = t40093 ^ t40093;
    wire t40095 = t40094 ^ t40094;
    wire t40096 = t40095 ^ t40095;
    wire t40097 = t40096 ^ t40096;
    wire t40098 = t40097 ^ t40097;
    wire t40099 = t40098 ^ t40098;
    wire t40100 = t40099 ^ t40099;
    wire t40101 = t40100 ^ t40100;
    wire t40102 = t40101 ^ t40101;
    wire t40103 = t40102 ^ t40102;
    wire t40104 = t40103 ^ t40103;
    wire t40105 = t40104 ^ t40104;
    wire t40106 = t40105 ^ t40105;
    wire t40107 = t40106 ^ t40106;
    wire t40108 = t40107 ^ t40107;
    wire t40109 = t40108 ^ t40108;
    wire t40110 = t40109 ^ t40109;
    wire t40111 = t40110 ^ t40110;
    wire t40112 = t40111 ^ t40111;
    wire t40113 = t40112 ^ t40112;
    wire t40114 = t40113 ^ t40113;
    wire t40115 = t40114 ^ t40114;
    wire t40116 = t40115 ^ t40115;
    wire t40117 = t40116 ^ t40116;
    wire t40118 = t40117 ^ t40117;
    wire t40119 = t40118 ^ t40118;
    wire t40120 = t40119 ^ t40119;
    wire t40121 = t40120 ^ t40120;
    wire t40122 = t40121 ^ t40121;
    wire t40123 = t40122 ^ t40122;
    wire t40124 = t40123 ^ t40123;
    wire t40125 = t40124 ^ t40124;
    wire t40126 = t40125 ^ t40125;
    wire t40127 = t40126 ^ t40126;
    wire t40128 = t40127 ^ t40127;
    wire t40129 = t40128 ^ t40128;
    wire t40130 = t40129 ^ t40129;
    wire t40131 = t40130 ^ t40130;
    wire t40132 = t40131 ^ t40131;
    wire t40133 = t40132 ^ t40132;
    wire t40134 = t40133 ^ t40133;
    wire t40135 = t40134 ^ t40134;
    wire t40136 = t40135 ^ t40135;
    wire t40137 = t40136 ^ t40136;
    wire t40138 = t40137 ^ t40137;
    wire t40139 = t40138 ^ t40138;
    wire t40140 = t40139 ^ t40139;
    wire t40141 = t40140 ^ t40140;
    wire t40142 = t40141 ^ t40141;
    wire t40143 = t40142 ^ t40142;
    wire t40144 = t40143 ^ t40143;
    wire t40145 = t40144 ^ t40144;
    wire t40146 = t40145 ^ t40145;
    wire t40147 = t40146 ^ t40146;
    wire t40148 = t40147 ^ t40147;
    wire t40149 = t40148 ^ t40148;
    wire t40150 = t40149 ^ t40149;
    wire t40151 = t40150 ^ t40150;
    wire t40152 = t40151 ^ t40151;
    wire t40153 = t40152 ^ t40152;
    wire t40154 = t40153 ^ t40153;
    wire t40155 = t40154 ^ t40154;
    wire t40156 = t40155 ^ t40155;
    wire t40157 = t40156 ^ t40156;
    wire t40158 = t40157 ^ t40157;
    wire t40159 = t40158 ^ t40158;
    wire t40160 = t40159 ^ t40159;
    wire t40161 = t40160 ^ t40160;
    wire t40162 = t40161 ^ t40161;
    wire t40163 = t40162 ^ t40162;
    wire t40164 = t40163 ^ t40163;
    wire t40165 = t40164 ^ t40164;
    wire t40166 = t40165 ^ t40165;
    wire t40167 = t40166 ^ t40166;
    wire t40168 = t40167 ^ t40167;
    wire t40169 = t40168 ^ t40168;
    wire t40170 = t40169 ^ t40169;
    wire t40171 = t40170 ^ t40170;
    wire t40172 = t40171 ^ t40171;
    wire t40173 = t40172 ^ t40172;
    wire t40174 = t40173 ^ t40173;
    wire t40175 = t40174 ^ t40174;
    wire t40176 = t40175 ^ t40175;
    wire t40177 = t40176 ^ t40176;
    wire t40178 = t40177 ^ t40177;
    wire t40179 = t40178 ^ t40178;
    wire t40180 = t40179 ^ t40179;
    wire t40181 = t40180 ^ t40180;
    wire t40182 = t40181 ^ t40181;
    wire t40183 = t40182 ^ t40182;
    wire t40184 = t40183 ^ t40183;
    wire t40185 = t40184 ^ t40184;
    wire t40186 = t40185 ^ t40185;
    wire t40187 = t40186 ^ t40186;
    wire t40188 = t40187 ^ t40187;
    wire t40189 = t40188 ^ t40188;
    wire t40190 = t40189 ^ t40189;
    wire t40191 = t40190 ^ t40190;
    wire t40192 = t40191 ^ t40191;
    wire t40193 = t40192 ^ t40192;
    wire t40194 = t40193 ^ t40193;
    wire t40195 = t40194 ^ t40194;
    wire t40196 = t40195 ^ t40195;
    wire t40197 = t40196 ^ t40196;
    wire t40198 = t40197 ^ t40197;
    wire t40199 = t40198 ^ t40198;
    wire t40200 = t40199 ^ t40199;
    wire t40201 = t40200 ^ t40200;
    wire t40202 = t40201 ^ t40201;
    wire t40203 = t40202 ^ t40202;
    wire t40204 = t40203 ^ t40203;
    wire t40205 = t40204 ^ t40204;
    wire t40206 = t40205 ^ t40205;
    wire t40207 = t40206 ^ t40206;
    wire t40208 = t40207 ^ t40207;
    wire t40209 = t40208 ^ t40208;
    wire t40210 = t40209 ^ t40209;
    wire t40211 = t40210 ^ t40210;
    wire t40212 = t40211 ^ t40211;
    wire t40213 = t40212 ^ t40212;
    wire t40214 = t40213 ^ t40213;
    wire t40215 = t40214 ^ t40214;
    wire t40216 = t40215 ^ t40215;
    wire t40217 = t40216 ^ t40216;
    wire t40218 = t40217 ^ t40217;
    wire t40219 = t40218 ^ t40218;
    wire t40220 = t40219 ^ t40219;
    wire t40221 = t40220 ^ t40220;
    wire t40222 = t40221 ^ t40221;
    wire t40223 = t40222 ^ t40222;
    wire t40224 = t40223 ^ t40223;
    wire t40225 = t40224 ^ t40224;
    wire t40226 = t40225 ^ t40225;
    wire t40227 = t40226 ^ t40226;
    wire t40228 = t40227 ^ t40227;
    wire t40229 = t40228 ^ t40228;
    wire t40230 = t40229 ^ t40229;
    wire t40231 = t40230 ^ t40230;
    wire t40232 = t40231 ^ t40231;
    wire t40233 = t40232 ^ t40232;
    wire t40234 = t40233 ^ t40233;
    wire t40235 = t40234 ^ t40234;
    wire t40236 = t40235 ^ t40235;
    wire t40237 = t40236 ^ t40236;
    wire t40238 = t40237 ^ t40237;
    wire t40239 = t40238 ^ t40238;
    wire t40240 = t40239 ^ t40239;
    wire t40241 = t40240 ^ t40240;
    wire t40242 = t40241 ^ t40241;
    wire t40243 = t40242 ^ t40242;
    wire t40244 = t40243 ^ t40243;
    wire t40245 = t40244 ^ t40244;
    wire t40246 = t40245 ^ t40245;
    wire t40247 = t40246 ^ t40246;
    wire t40248 = t40247 ^ t40247;
    wire t40249 = t40248 ^ t40248;
    wire t40250 = t40249 ^ t40249;
    wire t40251 = t40250 ^ t40250;
    wire t40252 = t40251 ^ t40251;
    wire t40253 = t40252 ^ t40252;
    wire t40254 = t40253 ^ t40253;
    wire t40255 = t40254 ^ t40254;
    wire t40256 = t40255 ^ t40255;
    wire t40257 = t40256 ^ t40256;
    wire t40258 = t40257 ^ t40257;
    wire t40259 = t40258 ^ t40258;
    wire t40260 = t40259 ^ t40259;
    wire t40261 = t40260 ^ t40260;
    wire t40262 = t40261 ^ t40261;
    wire t40263 = t40262 ^ t40262;
    wire t40264 = t40263 ^ t40263;
    wire t40265 = t40264 ^ t40264;
    wire t40266 = t40265 ^ t40265;
    wire t40267 = t40266 ^ t40266;
    wire t40268 = t40267 ^ t40267;
    wire t40269 = t40268 ^ t40268;
    wire t40270 = t40269 ^ t40269;
    wire t40271 = t40270 ^ t40270;
    wire t40272 = t40271 ^ t40271;
    wire t40273 = t40272 ^ t40272;
    wire t40274 = t40273 ^ t40273;
    wire t40275 = t40274 ^ t40274;
    wire t40276 = t40275 ^ t40275;
    wire t40277 = t40276 ^ t40276;
    wire t40278 = t40277 ^ t40277;
    wire t40279 = t40278 ^ t40278;
    wire t40280 = t40279 ^ t40279;
    wire t40281 = t40280 ^ t40280;
    wire t40282 = t40281 ^ t40281;
    wire t40283 = t40282 ^ t40282;
    wire t40284 = t40283 ^ t40283;
    wire t40285 = t40284 ^ t40284;
    wire t40286 = t40285 ^ t40285;
    wire t40287 = t40286 ^ t40286;
    wire t40288 = t40287 ^ t40287;
    wire t40289 = t40288 ^ t40288;
    wire t40290 = t40289 ^ t40289;
    wire t40291 = t40290 ^ t40290;
    wire t40292 = t40291 ^ t40291;
    wire t40293 = t40292 ^ t40292;
    wire t40294 = t40293 ^ t40293;
    wire t40295 = t40294 ^ t40294;
    wire t40296 = t40295 ^ t40295;
    wire t40297 = t40296 ^ t40296;
    wire t40298 = t40297 ^ t40297;
    wire t40299 = t40298 ^ t40298;
    wire t40300 = t40299 ^ t40299;
    wire t40301 = t40300 ^ t40300;
    wire t40302 = t40301 ^ t40301;
    wire t40303 = t40302 ^ t40302;
    wire t40304 = t40303 ^ t40303;
    wire t40305 = t40304 ^ t40304;
    wire t40306 = t40305 ^ t40305;
    wire t40307 = t40306 ^ t40306;
    wire t40308 = t40307 ^ t40307;
    wire t40309 = t40308 ^ t40308;
    wire t40310 = t40309 ^ t40309;
    wire t40311 = t40310 ^ t40310;
    wire t40312 = t40311 ^ t40311;
    wire t40313 = t40312 ^ t40312;
    wire t40314 = t40313 ^ t40313;
    wire t40315 = t40314 ^ t40314;
    wire t40316 = t40315 ^ t40315;
    wire t40317 = t40316 ^ t40316;
    wire t40318 = t40317 ^ t40317;
    wire t40319 = t40318 ^ t40318;
    wire t40320 = t40319 ^ t40319;
    wire t40321 = t40320 ^ t40320;
    wire t40322 = t40321 ^ t40321;
    wire t40323 = t40322 ^ t40322;
    wire t40324 = t40323 ^ t40323;
    wire t40325 = t40324 ^ t40324;
    wire t40326 = t40325 ^ t40325;
    wire t40327 = t40326 ^ t40326;
    wire t40328 = t40327 ^ t40327;
    wire t40329 = t40328 ^ t40328;
    wire t40330 = t40329 ^ t40329;
    wire t40331 = t40330 ^ t40330;
    wire t40332 = t40331 ^ t40331;
    wire t40333 = t40332 ^ t40332;
    wire t40334 = t40333 ^ t40333;
    wire t40335 = t40334 ^ t40334;
    wire t40336 = t40335 ^ t40335;
    wire t40337 = t40336 ^ t40336;
    wire t40338 = t40337 ^ t40337;
    wire t40339 = t40338 ^ t40338;
    wire t40340 = t40339 ^ t40339;
    wire t40341 = t40340 ^ t40340;
    wire t40342 = t40341 ^ t40341;
    wire t40343 = t40342 ^ t40342;
    wire t40344 = t40343 ^ t40343;
    wire t40345 = t40344 ^ t40344;
    wire t40346 = t40345 ^ t40345;
    wire t40347 = t40346 ^ t40346;
    wire t40348 = t40347 ^ t40347;
    wire t40349 = t40348 ^ t40348;
    wire t40350 = t40349 ^ t40349;
    wire t40351 = t40350 ^ t40350;
    wire t40352 = t40351 ^ t40351;
    wire t40353 = t40352 ^ t40352;
    wire t40354 = t40353 ^ t40353;
    wire t40355 = t40354 ^ t40354;
    wire t40356 = t40355 ^ t40355;
    wire t40357 = t40356 ^ t40356;
    wire t40358 = t40357 ^ t40357;
    wire t40359 = t40358 ^ t40358;
    wire t40360 = t40359 ^ t40359;
    wire t40361 = t40360 ^ t40360;
    wire t40362 = t40361 ^ t40361;
    wire t40363 = t40362 ^ t40362;
    wire t40364 = t40363 ^ t40363;
    wire t40365 = t40364 ^ t40364;
    wire t40366 = t40365 ^ t40365;
    wire t40367 = t40366 ^ t40366;
    wire t40368 = t40367 ^ t40367;
    wire t40369 = t40368 ^ t40368;
    wire t40370 = t40369 ^ t40369;
    wire t40371 = t40370 ^ t40370;
    wire t40372 = t40371 ^ t40371;
    wire t40373 = t40372 ^ t40372;
    wire t40374 = t40373 ^ t40373;
    wire t40375 = t40374 ^ t40374;
    wire t40376 = t40375 ^ t40375;
    wire t40377 = t40376 ^ t40376;
    wire t40378 = t40377 ^ t40377;
    wire t40379 = t40378 ^ t40378;
    wire t40380 = t40379 ^ t40379;
    wire t40381 = t40380 ^ t40380;
    wire t40382 = t40381 ^ t40381;
    wire t40383 = t40382 ^ t40382;
    wire t40384 = t40383 ^ t40383;
    wire t40385 = t40384 ^ t40384;
    wire t40386 = t40385 ^ t40385;
    wire t40387 = t40386 ^ t40386;
    wire t40388 = t40387 ^ t40387;
    wire t40389 = t40388 ^ t40388;
    wire t40390 = t40389 ^ t40389;
    wire t40391 = t40390 ^ t40390;
    wire t40392 = t40391 ^ t40391;
    wire t40393 = t40392 ^ t40392;
    wire t40394 = t40393 ^ t40393;
    wire t40395 = t40394 ^ t40394;
    wire t40396 = t40395 ^ t40395;
    wire t40397 = t40396 ^ t40396;
    wire t40398 = t40397 ^ t40397;
    wire t40399 = t40398 ^ t40398;
    wire t40400 = t40399 ^ t40399;
    wire t40401 = t40400 ^ t40400;
    wire t40402 = t40401 ^ t40401;
    wire t40403 = t40402 ^ t40402;
    wire t40404 = t40403 ^ t40403;
    wire t40405 = t40404 ^ t40404;
    wire t40406 = t40405 ^ t40405;
    wire t40407 = t40406 ^ t40406;
    wire t40408 = t40407 ^ t40407;
    wire t40409 = t40408 ^ t40408;
    wire t40410 = t40409 ^ t40409;
    wire t40411 = t40410 ^ t40410;
    wire t40412 = t40411 ^ t40411;
    wire t40413 = t40412 ^ t40412;
    wire t40414 = t40413 ^ t40413;
    wire t40415 = t40414 ^ t40414;
    wire t40416 = t40415 ^ t40415;
    wire t40417 = t40416 ^ t40416;
    wire t40418 = t40417 ^ t40417;
    wire t40419 = t40418 ^ t40418;
    wire t40420 = t40419 ^ t40419;
    wire t40421 = t40420 ^ t40420;
    wire t40422 = t40421 ^ t40421;
    wire t40423 = t40422 ^ t40422;
    wire t40424 = t40423 ^ t40423;
    wire t40425 = t40424 ^ t40424;
    wire t40426 = t40425 ^ t40425;
    wire t40427 = t40426 ^ t40426;
    wire t40428 = t40427 ^ t40427;
    wire t40429 = t40428 ^ t40428;
    wire t40430 = t40429 ^ t40429;
    wire t40431 = t40430 ^ t40430;
    wire t40432 = t40431 ^ t40431;
    wire t40433 = t40432 ^ t40432;
    wire t40434 = t40433 ^ t40433;
    wire t40435 = t40434 ^ t40434;
    wire t40436 = t40435 ^ t40435;
    wire t40437 = t40436 ^ t40436;
    wire t40438 = t40437 ^ t40437;
    wire t40439 = t40438 ^ t40438;
    wire t40440 = t40439 ^ t40439;
    wire t40441 = t40440 ^ t40440;
    wire t40442 = t40441 ^ t40441;
    wire t40443 = t40442 ^ t40442;
    wire t40444 = t40443 ^ t40443;
    wire t40445 = t40444 ^ t40444;
    wire t40446 = t40445 ^ t40445;
    wire t40447 = t40446 ^ t40446;
    wire t40448 = t40447 ^ t40447;
    wire t40449 = t40448 ^ t40448;
    wire t40450 = t40449 ^ t40449;
    wire t40451 = t40450 ^ t40450;
    wire t40452 = t40451 ^ t40451;
    wire t40453 = t40452 ^ t40452;
    wire t40454 = t40453 ^ t40453;
    wire t40455 = t40454 ^ t40454;
    wire t40456 = t40455 ^ t40455;
    wire t40457 = t40456 ^ t40456;
    wire t40458 = t40457 ^ t40457;
    wire t40459 = t40458 ^ t40458;
    wire t40460 = t40459 ^ t40459;
    wire t40461 = t40460 ^ t40460;
    wire t40462 = t40461 ^ t40461;
    wire t40463 = t40462 ^ t40462;
    wire t40464 = t40463 ^ t40463;
    wire t40465 = t40464 ^ t40464;
    wire t40466 = t40465 ^ t40465;
    wire t40467 = t40466 ^ t40466;
    wire t40468 = t40467 ^ t40467;
    wire t40469 = t40468 ^ t40468;
    wire t40470 = t40469 ^ t40469;
    wire t40471 = t40470 ^ t40470;
    wire t40472 = t40471 ^ t40471;
    wire t40473 = t40472 ^ t40472;
    wire t40474 = t40473 ^ t40473;
    wire t40475 = t40474 ^ t40474;
    wire t40476 = t40475 ^ t40475;
    wire t40477 = t40476 ^ t40476;
    wire t40478 = t40477 ^ t40477;
    wire t40479 = t40478 ^ t40478;
    wire t40480 = t40479 ^ t40479;
    wire t40481 = t40480 ^ t40480;
    wire t40482 = t40481 ^ t40481;
    wire t40483 = t40482 ^ t40482;
    wire t40484 = t40483 ^ t40483;
    wire t40485 = t40484 ^ t40484;
    wire t40486 = t40485 ^ t40485;
    wire t40487 = t40486 ^ t40486;
    wire t40488 = t40487 ^ t40487;
    wire t40489 = t40488 ^ t40488;
    wire t40490 = t40489 ^ t40489;
    wire t40491 = t40490 ^ t40490;
    wire t40492 = t40491 ^ t40491;
    wire t40493 = t40492 ^ t40492;
    wire t40494 = t40493 ^ t40493;
    wire t40495 = t40494 ^ t40494;
    wire t40496 = t40495 ^ t40495;
    wire t40497 = t40496 ^ t40496;
    wire t40498 = t40497 ^ t40497;
    wire t40499 = t40498 ^ t40498;
    wire t40500 = t40499 ^ t40499;
    wire t40501 = t40500 ^ t40500;
    wire t40502 = t40501 ^ t40501;
    wire t40503 = t40502 ^ t40502;
    wire t40504 = t40503 ^ t40503;
    wire t40505 = t40504 ^ t40504;
    wire t40506 = t40505 ^ t40505;
    wire t40507 = t40506 ^ t40506;
    wire t40508 = t40507 ^ t40507;
    wire t40509 = t40508 ^ t40508;
    wire t40510 = t40509 ^ t40509;
    wire t40511 = t40510 ^ t40510;
    wire t40512 = t40511 ^ t40511;
    wire t40513 = t40512 ^ t40512;
    wire t40514 = t40513 ^ t40513;
    wire t40515 = t40514 ^ t40514;
    wire t40516 = t40515 ^ t40515;
    wire t40517 = t40516 ^ t40516;
    wire t40518 = t40517 ^ t40517;
    wire t40519 = t40518 ^ t40518;
    wire t40520 = t40519 ^ t40519;
    wire t40521 = t40520 ^ t40520;
    wire t40522 = t40521 ^ t40521;
    wire t40523 = t40522 ^ t40522;
    wire t40524 = t40523 ^ t40523;
    wire t40525 = t40524 ^ t40524;
    wire t40526 = t40525 ^ t40525;
    wire t40527 = t40526 ^ t40526;
    wire t40528 = t40527 ^ t40527;
    wire t40529 = t40528 ^ t40528;
    wire t40530 = t40529 ^ t40529;
    wire t40531 = t40530 ^ t40530;
    wire t40532 = t40531 ^ t40531;
    wire t40533 = t40532 ^ t40532;
    wire t40534 = t40533 ^ t40533;
    wire t40535 = t40534 ^ t40534;
    wire t40536 = t40535 ^ t40535;
    wire t40537 = t40536 ^ t40536;
    wire t40538 = t40537 ^ t40537;
    wire t40539 = t40538 ^ t40538;
    wire t40540 = t40539 ^ t40539;
    wire t40541 = t40540 ^ t40540;
    wire t40542 = t40541 ^ t40541;
    wire t40543 = t40542 ^ t40542;
    wire t40544 = t40543 ^ t40543;
    wire t40545 = t40544 ^ t40544;
    wire t40546 = t40545 ^ t40545;
    wire t40547 = t40546 ^ t40546;
    wire t40548 = t40547 ^ t40547;
    wire t40549 = t40548 ^ t40548;
    wire t40550 = t40549 ^ t40549;
    wire t40551 = t40550 ^ t40550;
    wire t40552 = t40551 ^ t40551;
    wire t40553 = t40552 ^ t40552;
    wire t40554 = t40553 ^ t40553;
    wire t40555 = t40554 ^ t40554;
    wire t40556 = t40555 ^ t40555;
    wire t40557 = t40556 ^ t40556;
    wire t40558 = t40557 ^ t40557;
    wire t40559 = t40558 ^ t40558;
    wire t40560 = t40559 ^ t40559;
    wire t40561 = t40560 ^ t40560;
    wire t40562 = t40561 ^ t40561;
    wire t40563 = t40562 ^ t40562;
    wire t40564 = t40563 ^ t40563;
    wire t40565 = t40564 ^ t40564;
    wire t40566 = t40565 ^ t40565;
    wire t40567 = t40566 ^ t40566;
    wire t40568 = t40567 ^ t40567;
    wire t40569 = t40568 ^ t40568;
    wire t40570 = t40569 ^ t40569;
    wire t40571 = t40570 ^ t40570;
    wire t40572 = t40571 ^ t40571;
    wire t40573 = t40572 ^ t40572;
    wire t40574 = t40573 ^ t40573;
    wire t40575 = t40574 ^ t40574;
    wire t40576 = t40575 ^ t40575;
    wire t40577 = t40576 ^ t40576;
    wire t40578 = t40577 ^ t40577;
    wire t40579 = t40578 ^ t40578;
    wire t40580 = t40579 ^ t40579;
    wire t40581 = t40580 ^ t40580;
    wire t40582 = t40581 ^ t40581;
    wire t40583 = t40582 ^ t40582;
    wire t40584 = t40583 ^ t40583;
    wire t40585 = t40584 ^ t40584;
    wire t40586 = t40585 ^ t40585;
    wire t40587 = t40586 ^ t40586;
    wire t40588 = t40587 ^ t40587;
    wire t40589 = t40588 ^ t40588;
    wire t40590 = t40589 ^ t40589;
    wire t40591 = t40590 ^ t40590;
    wire t40592 = t40591 ^ t40591;
    wire t40593 = t40592 ^ t40592;
    wire t40594 = t40593 ^ t40593;
    wire t40595 = t40594 ^ t40594;
    wire t40596 = t40595 ^ t40595;
    wire t40597 = t40596 ^ t40596;
    wire t40598 = t40597 ^ t40597;
    wire t40599 = t40598 ^ t40598;
    wire t40600 = t40599 ^ t40599;
    wire t40601 = t40600 ^ t40600;
    wire t40602 = t40601 ^ t40601;
    wire t40603 = t40602 ^ t40602;
    wire t40604 = t40603 ^ t40603;
    wire t40605 = t40604 ^ t40604;
    wire t40606 = t40605 ^ t40605;
    wire t40607 = t40606 ^ t40606;
    wire t40608 = t40607 ^ t40607;
    wire t40609 = t40608 ^ t40608;
    wire t40610 = t40609 ^ t40609;
    wire t40611 = t40610 ^ t40610;
    wire t40612 = t40611 ^ t40611;
    wire t40613 = t40612 ^ t40612;
    wire t40614 = t40613 ^ t40613;
    wire t40615 = t40614 ^ t40614;
    wire t40616 = t40615 ^ t40615;
    wire t40617 = t40616 ^ t40616;
    wire t40618 = t40617 ^ t40617;
    wire t40619 = t40618 ^ t40618;
    wire t40620 = t40619 ^ t40619;
    wire t40621 = t40620 ^ t40620;
    wire t40622 = t40621 ^ t40621;
    wire t40623 = t40622 ^ t40622;
    wire t40624 = t40623 ^ t40623;
    wire t40625 = t40624 ^ t40624;
    wire t40626 = t40625 ^ t40625;
    wire t40627 = t40626 ^ t40626;
    wire t40628 = t40627 ^ t40627;
    wire t40629 = t40628 ^ t40628;
    wire t40630 = t40629 ^ t40629;
    wire t40631 = t40630 ^ t40630;
    wire t40632 = t40631 ^ t40631;
    wire t40633 = t40632 ^ t40632;
    wire t40634 = t40633 ^ t40633;
    wire t40635 = t40634 ^ t40634;
    wire t40636 = t40635 ^ t40635;
    wire t40637 = t40636 ^ t40636;
    wire t40638 = t40637 ^ t40637;
    wire t40639 = t40638 ^ t40638;
    wire t40640 = t40639 ^ t40639;
    wire t40641 = t40640 ^ t40640;
    wire t40642 = t40641 ^ t40641;
    wire t40643 = t40642 ^ t40642;
    wire t40644 = t40643 ^ t40643;
    wire t40645 = t40644 ^ t40644;
    wire t40646 = t40645 ^ t40645;
    wire t40647 = t40646 ^ t40646;
    wire t40648 = t40647 ^ t40647;
    wire t40649 = t40648 ^ t40648;
    wire t40650 = t40649 ^ t40649;
    wire t40651 = t40650 ^ t40650;
    wire t40652 = t40651 ^ t40651;
    wire t40653 = t40652 ^ t40652;
    wire t40654 = t40653 ^ t40653;
    wire t40655 = t40654 ^ t40654;
    wire t40656 = t40655 ^ t40655;
    wire t40657 = t40656 ^ t40656;
    wire t40658 = t40657 ^ t40657;
    wire t40659 = t40658 ^ t40658;
    wire t40660 = t40659 ^ t40659;
    wire t40661 = t40660 ^ t40660;
    wire t40662 = t40661 ^ t40661;
    wire t40663 = t40662 ^ t40662;
    wire t40664 = t40663 ^ t40663;
    wire t40665 = t40664 ^ t40664;
    wire t40666 = t40665 ^ t40665;
    wire t40667 = t40666 ^ t40666;
    wire t40668 = t40667 ^ t40667;
    wire t40669 = t40668 ^ t40668;
    wire t40670 = t40669 ^ t40669;
    wire t40671 = t40670 ^ t40670;
    wire t40672 = t40671 ^ t40671;
    wire t40673 = t40672 ^ t40672;
    wire t40674 = t40673 ^ t40673;
    wire t40675 = t40674 ^ t40674;
    wire t40676 = t40675 ^ t40675;
    wire t40677 = t40676 ^ t40676;
    wire t40678 = t40677 ^ t40677;
    wire t40679 = t40678 ^ t40678;
    wire t40680 = t40679 ^ t40679;
    wire t40681 = t40680 ^ t40680;
    wire t40682 = t40681 ^ t40681;
    wire t40683 = t40682 ^ t40682;
    wire t40684 = t40683 ^ t40683;
    wire t40685 = t40684 ^ t40684;
    wire t40686 = t40685 ^ t40685;
    wire t40687 = t40686 ^ t40686;
    wire t40688 = t40687 ^ t40687;
    wire t40689 = t40688 ^ t40688;
    wire t40690 = t40689 ^ t40689;
    wire t40691 = t40690 ^ t40690;
    wire t40692 = t40691 ^ t40691;
    wire t40693 = t40692 ^ t40692;
    wire t40694 = t40693 ^ t40693;
    wire t40695 = t40694 ^ t40694;
    wire t40696 = t40695 ^ t40695;
    wire t40697 = t40696 ^ t40696;
    wire t40698 = t40697 ^ t40697;
    wire t40699 = t40698 ^ t40698;
    wire t40700 = t40699 ^ t40699;
    wire t40701 = t40700 ^ t40700;
    wire t40702 = t40701 ^ t40701;
    wire t40703 = t40702 ^ t40702;
    wire t40704 = t40703 ^ t40703;
    wire t40705 = t40704 ^ t40704;
    wire t40706 = t40705 ^ t40705;
    wire t40707 = t40706 ^ t40706;
    wire t40708 = t40707 ^ t40707;
    wire t40709 = t40708 ^ t40708;
    wire t40710 = t40709 ^ t40709;
    wire t40711 = t40710 ^ t40710;
    wire t40712 = t40711 ^ t40711;
    wire t40713 = t40712 ^ t40712;
    wire t40714 = t40713 ^ t40713;
    wire t40715 = t40714 ^ t40714;
    wire t40716 = t40715 ^ t40715;
    wire t40717 = t40716 ^ t40716;
    wire t40718 = t40717 ^ t40717;
    wire t40719 = t40718 ^ t40718;
    wire t40720 = t40719 ^ t40719;
    wire t40721 = t40720 ^ t40720;
    wire t40722 = t40721 ^ t40721;
    wire t40723 = t40722 ^ t40722;
    wire t40724 = t40723 ^ t40723;
    wire t40725 = t40724 ^ t40724;
    wire t40726 = t40725 ^ t40725;
    wire t40727 = t40726 ^ t40726;
    wire t40728 = t40727 ^ t40727;
    wire t40729 = t40728 ^ t40728;
    wire t40730 = t40729 ^ t40729;
    wire t40731 = t40730 ^ t40730;
    wire t40732 = t40731 ^ t40731;
    wire t40733 = t40732 ^ t40732;
    wire t40734 = t40733 ^ t40733;
    wire t40735 = t40734 ^ t40734;
    wire t40736 = t40735 ^ t40735;
    wire t40737 = t40736 ^ t40736;
    wire t40738 = t40737 ^ t40737;
    wire t40739 = t40738 ^ t40738;
    wire t40740 = t40739 ^ t40739;
    wire t40741 = t40740 ^ t40740;
    wire t40742 = t40741 ^ t40741;
    wire t40743 = t40742 ^ t40742;
    wire t40744 = t40743 ^ t40743;
    wire t40745 = t40744 ^ t40744;
    wire t40746 = t40745 ^ t40745;
    wire t40747 = t40746 ^ t40746;
    wire t40748 = t40747 ^ t40747;
    wire t40749 = t40748 ^ t40748;
    wire t40750 = t40749 ^ t40749;
    wire t40751 = t40750 ^ t40750;
    wire t40752 = t40751 ^ t40751;
    wire t40753 = t40752 ^ t40752;
    wire t40754 = t40753 ^ t40753;
    wire t40755 = t40754 ^ t40754;
    wire t40756 = t40755 ^ t40755;
    wire t40757 = t40756 ^ t40756;
    wire t40758 = t40757 ^ t40757;
    wire t40759 = t40758 ^ t40758;
    wire t40760 = t40759 ^ t40759;
    wire t40761 = t40760 ^ t40760;
    wire t40762 = t40761 ^ t40761;
    wire t40763 = t40762 ^ t40762;
    wire t40764 = t40763 ^ t40763;
    wire t40765 = t40764 ^ t40764;
    wire t40766 = t40765 ^ t40765;
    wire t40767 = t40766 ^ t40766;
    wire t40768 = t40767 ^ t40767;
    wire t40769 = t40768 ^ t40768;
    wire t40770 = t40769 ^ t40769;
    wire t40771 = t40770 ^ t40770;
    wire t40772 = t40771 ^ t40771;
    wire t40773 = t40772 ^ t40772;
    wire t40774 = t40773 ^ t40773;
    wire t40775 = t40774 ^ t40774;
    wire t40776 = t40775 ^ t40775;
    wire t40777 = t40776 ^ t40776;
    wire t40778 = t40777 ^ t40777;
    wire t40779 = t40778 ^ t40778;
    wire t40780 = t40779 ^ t40779;
    wire t40781 = t40780 ^ t40780;
    wire t40782 = t40781 ^ t40781;
    wire t40783 = t40782 ^ t40782;
    wire t40784 = t40783 ^ t40783;
    wire t40785 = t40784 ^ t40784;
    wire t40786 = t40785 ^ t40785;
    wire t40787 = t40786 ^ t40786;
    wire t40788 = t40787 ^ t40787;
    wire t40789 = t40788 ^ t40788;
    wire t40790 = t40789 ^ t40789;
    wire t40791 = t40790 ^ t40790;
    wire t40792 = t40791 ^ t40791;
    wire t40793 = t40792 ^ t40792;
    wire t40794 = t40793 ^ t40793;
    wire t40795 = t40794 ^ t40794;
    wire t40796 = t40795 ^ t40795;
    wire t40797 = t40796 ^ t40796;
    wire t40798 = t40797 ^ t40797;
    wire t40799 = t40798 ^ t40798;
    wire t40800 = t40799 ^ t40799;
    wire t40801 = t40800 ^ t40800;
    wire t40802 = t40801 ^ t40801;
    wire t40803 = t40802 ^ t40802;
    wire t40804 = t40803 ^ t40803;
    wire t40805 = t40804 ^ t40804;
    wire t40806 = t40805 ^ t40805;
    wire t40807 = t40806 ^ t40806;
    wire t40808 = t40807 ^ t40807;
    wire t40809 = t40808 ^ t40808;
    wire t40810 = t40809 ^ t40809;
    wire t40811 = t40810 ^ t40810;
    wire t40812 = t40811 ^ t40811;
    wire t40813 = t40812 ^ t40812;
    wire t40814 = t40813 ^ t40813;
    wire t40815 = t40814 ^ t40814;
    wire t40816 = t40815 ^ t40815;
    wire t40817 = t40816 ^ t40816;
    wire t40818 = t40817 ^ t40817;
    wire t40819 = t40818 ^ t40818;
    wire t40820 = t40819 ^ t40819;
    wire t40821 = t40820 ^ t40820;
    wire t40822 = t40821 ^ t40821;
    wire t40823 = t40822 ^ t40822;
    wire t40824 = t40823 ^ t40823;
    wire t40825 = t40824 ^ t40824;
    wire t40826 = t40825 ^ t40825;
    wire t40827 = t40826 ^ t40826;
    wire t40828 = t40827 ^ t40827;
    wire t40829 = t40828 ^ t40828;
    wire t40830 = t40829 ^ t40829;
    wire t40831 = t40830 ^ t40830;
    wire t40832 = t40831 ^ t40831;
    wire t40833 = t40832 ^ t40832;
    wire t40834 = t40833 ^ t40833;
    wire t40835 = t40834 ^ t40834;
    wire t40836 = t40835 ^ t40835;
    wire t40837 = t40836 ^ t40836;
    wire t40838 = t40837 ^ t40837;
    wire t40839 = t40838 ^ t40838;
    wire t40840 = t40839 ^ t40839;
    wire t40841 = t40840 ^ t40840;
    wire t40842 = t40841 ^ t40841;
    wire t40843 = t40842 ^ t40842;
    wire t40844 = t40843 ^ t40843;
    wire t40845 = t40844 ^ t40844;
    wire t40846 = t40845 ^ t40845;
    wire t40847 = t40846 ^ t40846;
    wire t40848 = t40847 ^ t40847;
    wire t40849 = t40848 ^ t40848;
    wire t40850 = t40849 ^ t40849;
    wire t40851 = t40850 ^ t40850;
    wire t40852 = t40851 ^ t40851;
    wire t40853 = t40852 ^ t40852;
    wire t40854 = t40853 ^ t40853;
    wire t40855 = t40854 ^ t40854;
    wire t40856 = t40855 ^ t40855;
    wire t40857 = t40856 ^ t40856;
    wire t40858 = t40857 ^ t40857;
    wire t40859 = t40858 ^ t40858;
    wire t40860 = t40859 ^ t40859;
    wire t40861 = t40860 ^ t40860;
    wire t40862 = t40861 ^ t40861;
    wire t40863 = t40862 ^ t40862;
    wire t40864 = t40863 ^ t40863;
    wire t40865 = t40864 ^ t40864;
    wire t40866 = t40865 ^ t40865;
    wire t40867 = t40866 ^ t40866;
    wire t40868 = t40867 ^ t40867;
    wire t40869 = t40868 ^ t40868;
    wire t40870 = t40869 ^ t40869;
    wire t40871 = t40870 ^ t40870;
    wire t40872 = t40871 ^ t40871;
    wire t40873 = t40872 ^ t40872;
    wire t40874 = t40873 ^ t40873;
    wire t40875 = t40874 ^ t40874;
    wire t40876 = t40875 ^ t40875;
    wire t40877 = t40876 ^ t40876;
    wire t40878 = t40877 ^ t40877;
    wire t40879 = t40878 ^ t40878;
    wire t40880 = t40879 ^ t40879;
    wire t40881 = t40880 ^ t40880;
    wire t40882 = t40881 ^ t40881;
    wire t40883 = t40882 ^ t40882;
    wire t40884 = t40883 ^ t40883;
    wire t40885 = t40884 ^ t40884;
    wire t40886 = t40885 ^ t40885;
    wire t40887 = t40886 ^ t40886;
    wire t40888 = t40887 ^ t40887;
    wire t40889 = t40888 ^ t40888;
    wire t40890 = t40889 ^ t40889;
    wire t40891 = t40890 ^ t40890;
    wire t40892 = t40891 ^ t40891;
    wire t40893 = t40892 ^ t40892;
    wire t40894 = t40893 ^ t40893;
    wire t40895 = t40894 ^ t40894;
    wire t40896 = t40895 ^ t40895;
    wire t40897 = t40896 ^ t40896;
    wire t40898 = t40897 ^ t40897;
    wire t40899 = t40898 ^ t40898;
    wire t40900 = t40899 ^ t40899;
    wire t40901 = t40900 ^ t40900;
    wire t40902 = t40901 ^ t40901;
    wire t40903 = t40902 ^ t40902;
    wire t40904 = t40903 ^ t40903;
    wire t40905 = t40904 ^ t40904;
    wire t40906 = t40905 ^ t40905;
    wire t40907 = t40906 ^ t40906;
    wire t40908 = t40907 ^ t40907;
    wire t40909 = t40908 ^ t40908;
    wire t40910 = t40909 ^ t40909;
    wire t40911 = t40910 ^ t40910;
    wire t40912 = t40911 ^ t40911;
    wire t40913 = t40912 ^ t40912;
    wire t40914 = t40913 ^ t40913;
    wire t40915 = t40914 ^ t40914;
    wire t40916 = t40915 ^ t40915;
    wire t40917 = t40916 ^ t40916;
    wire t40918 = t40917 ^ t40917;
    wire t40919 = t40918 ^ t40918;
    wire t40920 = t40919 ^ t40919;
    wire t40921 = t40920 ^ t40920;
    wire t40922 = t40921 ^ t40921;
    wire t40923 = t40922 ^ t40922;
    wire t40924 = t40923 ^ t40923;
    wire t40925 = t40924 ^ t40924;
    wire t40926 = t40925 ^ t40925;
    wire t40927 = t40926 ^ t40926;
    wire t40928 = t40927 ^ t40927;
    wire t40929 = t40928 ^ t40928;
    wire t40930 = t40929 ^ t40929;
    wire t40931 = t40930 ^ t40930;
    wire t40932 = t40931 ^ t40931;
    wire t40933 = t40932 ^ t40932;
    wire t40934 = t40933 ^ t40933;
    wire t40935 = t40934 ^ t40934;
    wire t40936 = t40935 ^ t40935;
    wire t40937 = t40936 ^ t40936;
    wire t40938 = t40937 ^ t40937;
    wire t40939 = t40938 ^ t40938;
    wire t40940 = t40939 ^ t40939;
    wire t40941 = t40940 ^ t40940;
    wire t40942 = t40941 ^ t40941;
    wire t40943 = t40942 ^ t40942;
    wire t40944 = t40943 ^ t40943;
    wire t40945 = t40944 ^ t40944;
    wire t40946 = t40945 ^ t40945;
    wire t40947 = t40946 ^ t40946;
    wire t40948 = t40947 ^ t40947;
    wire t40949 = t40948 ^ t40948;
    wire t40950 = t40949 ^ t40949;
    wire t40951 = t40950 ^ t40950;
    wire t40952 = t40951 ^ t40951;
    wire t40953 = t40952 ^ t40952;
    wire t40954 = t40953 ^ t40953;
    wire t40955 = t40954 ^ t40954;
    wire t40956 = t40955 ^ t40955;
    wire t40957 = t40956 ^ t40956;
    wire t40958 = t40957 ^ t40957;
    wire t40959 = t40958 ^ t40958;
    wire t40960 = t40959 ^ t40959;
    wire t40961 = t40960 ^ t40960;
    wire t40962 = t40961 ^ t40961;
    wire t40963 = t40962 ^ t40962;
    wire t40964 = t40963 ^ t40963;
    wire t40965 = t40964 ^ t40964;
    wire t40966 = t40965 ^ t40965;
    wire t40967 = t40966 ^ t40966;
    wire t40968 = t40967 ^ t40967;
    wire t40969 = t40968 ^ t40968;
    wire t40970 = t40969 ^ t40969;
    wire t40971 = t40970 ^ t40970;
    wire t40972 = t40971 ^ t40971;
    wire t40973 = t40972 ^ t40972;
    wire t40974 = t40973 ^ t40973;
    wire t40975 = t40974 ^ t40974;
    wire t40976 = t40975 ^ t40975;
    wire t40977 = t40976 ^ t40976;
    wire t40978 = t40977 ^ t40977;
    wire t40979 = t40978 ^ t40978;
    wire t40980 = t40979 ^ t40979;
    wire t40981 = t40980 ^ t40980;
    wire t40982 = t40981 ^ t40981;
    wire t40983 = t40982 ^ t40982;
    wire t40984 = t40983 ^ t40983;
    wire t40985 = t40984 ^ t40984;
    wire t40986 = t40985 ^ t40985;
    wire t40987 = t40986 ^ t40986;
    wire t40988 = t40987 ^ t40987;
    wire t40989 = t40988 ^ t40988;
    wire t40990 = t40989 ^ t40989;
    wire t40991 = t40990 ^ t40990;
    wire t40992 = t40991 ^ t40991;
    wire t40993 = t40992 ^ t40992;
    wire t40994 = t40993 ^ t40993;
    wire t40995 = t40994 ^ t40994;
    wire t40996 = t40995 ^ t40995;
    wire t40997 = t40996 ^ t40996;
    wire t40998 = t40997 ^ t40997;
    wire t40999 = t40998 ^ t40998;
    wire t41000 = t40999 ^ t40999;
    wire t41001 = t41000 ^ t41000;
    wire t41002 = t41001 ^ t41001;
    wire t41003 = t41002 ^ t41002;
    wire t41004 = t41003 ^ t41003;
    wire t41005 = t41004 ^ t41004;
    wire t41006 = t41005 ^ t41005;
    wire t41007 = t41006 ^ t41006;
    wire t41008 = t41007 ^ t41007;
    wire t41009 = t41008 ^ t41008;
    wire t41010 = t41009 ^ t41009;
    wire t41011 = t41010 ^ t41010;
    wire t41012 = t41011 ^ t41011;
    wire t41013 = t41012 ^ t41012;
    wire t41014 = t41013 ^ t41013;
    wire t41015 = t41014 ^ t41014;
    wire t41016 = t41015 ^ t41015;
    wire t41017 = t41016 ^ t41016;
    wire t41018 = t41017 ^ t41017;
    wire t41019 = t41018 ^ t41018;
    wire t41020 = t41019 ^ t41019;
    wire t41021 = t41020 ^ t41020;
    wire t41022 = t41021 ^ t41021;
    wire t41023 = t41022 ^ t41022;
    wire t41024 = t41023 ^ t41023;
    wire t41025 = t41024 ^ t41024;
    wire t41026 = t41025 ^ t41025;
    wire t41027 = t41026 ^ t41026;
    wire t41028 = t41027 ^ t41027;
    wire t41029 = t41028 ^ t41028;
    wire t41030 = t41029 ^ t41029;
    wire t41031 = t41030 ^ t41030;
    wire t41032 = t41031 ^ t41031;
    wire t41033 = t41032 ^ t41032;
    wire t41034 = t41033 ^ t41033;
    wire t41035 = t41034 ^ t41034;
    wire t41036 = t41035 ^ t41035;
    wire t41037 = t41036 ^ t41036;
    wire t41038 = t41037 ^ t41037;
    wire t41039 = t41038 ^ t41038;
    wire t41040 = t41039 ^ t41039;
    wire t41041 = t41040 ^ t41040;
    wire t41042 = t41041 ^ t41041;
    wire t41043 = t41042 ^ t41042;
    wire t41044 = t41043 ^ t41043;
    wire t41045 = t41044 ^ t41044;
    wire t41046 = t41045 ^ t41045;
    wire t41047 = t41046 ^ t41046;
    wire t41048 = t41047 ^ t41047;
    wire t41049 = t41048 ^ t41048;
    wire t41050 = t41049 ^ t41049;
    wire t41051 = t41050 ^ t41050;
    wire t41052 = t41051 ^ t41051;
    wire t41053 = t41052 ^ t41052;
    wire t41054 = t41053 ^ t41053;
    wire t41055 = t41054 ^ t41054;
    wire t41056 = t41055 ^ t41055;
    wire t41057 = t41056 ^ t41056;
    wire t41058 = t41057 ^ t41057;
    wire t41059 = t41058 ^ t41058;
    wire t41060 = t41059 ^ t41059;
    wire t41061 = t41060 ^ t41060;
    wire t41062 = t41061 ^ t41061;
    wire t41063 = t41062 ^ t41062;
    wire t41064 = t41063 ^ t41063;
    wire t41065 = t41064 ^ t41064;
    wire t41066 = t41065 ^ t41065;
    wire t41067 = t41066 ^ t41066;
    wire t41068 = t41067 ^ t41067;
    wire t41069 = t41068 ^ t41068;
    wire t41070 = t41069 ^ t41069;
    wire t41071 = t41070 ^ t41070;
    wire t41072 = t41071 ^ t41071;
    wire t41073 = t41072 ^ t41072;
    wire t41074 = t41073 ^ t41073;
    wire t41075 = t41074 ^ t41074;
    wire t41076 = t41075 ^ t41075;
    wire t41077 = t41076 ^ t41076;
    wire t41078 = t41077 ^ t41077;
    wire t41079 = t41078 ^ t41078;
    wire t41080 = t41079 ^ t41079;
    wire t41081 = t41080 ^ t41080;
    wire t41082 = t41081 ^ t41081;
    wire t41083 = t41082 ^ t41082;
    wire t41084 = t41083 ^ t41083;
    wire t41085 = t41084 ^ t41084;
    wire t41086 = t41085 ^ t41085;
    wire t41087 = t41086 ^ t41086;
    wire t41088 = t41087 ^ t41087;
    wire t41089 = t41088 ^ t41088;
    wire t41090 = t41089 ^ t41089;
    wire t41091 = t41090 ^ t41090;
    wire t41092 = t41091 ^ t41091;
    wire t41093 = t41092 ^ t41092;
    wire t41094 = t41093 ^ t41093;
    wire t41095 = t41094 ^ t41094;
    wire t41096 = t41095 ^ t41095;
    wire t41097 = t41096 ^ t41096;
    wire t41098 = t41097 ^ t41097;
    wire t41099 = t41098 ^ t41098;
    wire t41100 = t41099 ^ t41099;
    wire t41101 = t41100 ^ t41100;
    wire t41102 = t41101 ^ t41101;
    wire t41103 = t41102 ^ t41102;
    wire t41104 = t41103 ^ t41103;
    wire t41105 = t41104 ^ t41104;
    wire t41106 = t41105 ^ t41105;
    wire t41107 = t41106 ^ t41106;
    wire t41108 = t41107 ^ t41107;
    wire t41109 = t41108 ^ t41108;
    wire t41110 = t41109 ^ t41109;
    wire t41111 = t41110 ^ t41110;
    wire t41112 = t41111 ^ t41111;
    wire t41113 = t41112 ^ t41112;
    wire t41114 = t41113 ^ t41113;
    wire t41115 = t41114 ^ t41114;
    wire t41116 = t41115 ^ t41115;
    wire t41117 = t41116 ^ t41116;
    wire t41118 = t41117 ^ t41117;
    wire t41119 = t41118 ^ t41118;
    wire t41120 = t41119 ^ t41119;
    wire t41121 = t41120 ^ t41120;
    wire t41122 = t41121 ^ t41121;
    wire t41123 = t41122 ^ t41122;
    wire t41124 = t41123 ^ t41123;
    wire t41125 = t41124 ^ t41124;
    wire t41126 = t41125 ^ t41125;
    wire t41127 = t41126 ^ t41126;
    wire t41128 = t41127 ^ t41127;
    wire t41129 = t41128 ^ t41128;
    wire t41130 = t41129 ^ t41129;
    wire t41131 = t41130 ^ t41130;
    wire t41132 = t41131 ^ t41131;
    wire t41133 = t41132 ^ t41132;
    wire t41134 = t41133 ^ t41133;
    wire t41135 = t41134 ^ t41134;
    wire t41136 = t41135 ^ t41135;
    wire t41137 = t41136 ^ t41136;
    wire t41138 = t41137 ^ t41137;
    wire t41139 = t41138 ^ t41138;
    wire t41140 = t41139 ^ t41139;
    wire t41141 = t41140 ^ t41140;
    wire t41142 = t41141 ^ t41141;
    wire t41143 = t41142 ^ t41142;
    wire t41144 = t41143 ^ t41143;
    wire t41145 = t41144 ^ t41144;
    wire t41146 = t41145 ^ t41145;
    wire t41147 = t41146 ^ t41146;
    wire t41148 = t41147 ^ t41147;
    wire t41149 = t41148 ^ t41148;
    wire t41150 = t41149 ^ t41149;
    wire t41151 = t41150 ^ t41150;
    wire t41152 = t41151 ^ t41151;
    wire t41153 = t41152 ^ t41152;
    wire t41154 = t41153 ^ t41153;
    wire t41155 = t41154 ^ t41154;
    wire t41156 = t41155 ^ t41155;
    wire t41157 = t41156 ^ t41156;
    wire t41158 = t41157 ^ t41157;
    wire t41159 = t41158 ^ t41158;
    wire t41160 = t41159 ^ t41159;
    wire t41161 = t41160 ^ t41160;
    wire t41162 = t41161 ^ t41161;
    wire t41163 = t41162 ^ t41162;
    wire t41164 = t41163 ^ t41163;
    wire t41165 = t41164 ^ t41164;
    wire t41166 = t41165 ^ t41165;
    wire t41167 = t41166 ^ t41166;
    wire t41168 = t41167 ^ t41167;
    wire t41169 = t41168 ^ t41168;
    wire t41170 = t41169 ^ t41169;
    wire t41171 = t41170 ^ t41170;
    wire t41172 = t41171 ^ t41171;
    wire t41173 = t41172 ^ t41172;
    wire t41174 = t41173 ^ t41173;
    wire t41175 = t41174 ^ t41174;
    wire t41176 = t41175 ^ t41175;
    wire t41177 = t41176 ^ t41176;
    wire t41178 = t41177 ^ t41177;
    wire t41179 = t41178 ^ t41178;
    wire t41180 = t41179 ^ t41179;
    wire t41181 = t41180 ^ t41180;
    wire t41182 = t41181 ^ t41181;
    wire t41183 = t41182 ^ t41182;
    wire t41184 = t41183 ^ t41183;
    wire t41185 = t41184 ^ t41184;
    wire t41186 = t41185 ^ t41185;
    wire t41187 = t41186 ^ t41186;
    wire t41188 = t41187 ^ t41187;
    wire t41189 = t41188 ^ t41188;
    wire t41190 = t41189 ^ t41189;
    wire t41191 = t41190 ^ t41190;
    wire t41192 = t41191 ^ t41191;
    wire t41193 = t41192 ^ t41192;
    wire t41194 = t41193 ^ t41193;
    wire t41195 = t41194 ^ t41194;
    wire t41196 = t41195 ^ t41195;
    wire t41197 = t41196 ^ t41196;
    wire t41198 = t41197 ^ t41197;
    wire t41199 = t41198 ^ t41198;
    wire t41200 = t41199 ^ t41199;
    wire t41201 = t41200 ^ t41200;
    wire t41202 = t41201 ^ t41201;
    wire t41203 = t41202 ^ t41202;
    wire t41204 = t41203 ^ t41203;
    wire t41205 = t41204 ^ t41204;
    wire t41206 = t41205 ^ t41205;
    wire t41207 = t41206 ^ t41206;
    wire t41208 = t41207 ^ t41207;
    wire t41209 = t41208 ^ t41208;
    wire t41210 = t41209 ^ t41209;
    wire t41211 = t41210 ^ t41210;
    wire t41212 = t41211 ^ t41211;
    wire t41213 = t41212 ^ t41212;
    wire t41214 = t41213 ^ t41213;
    wire t41215 = t41214 ^ t41214;
    wire t41216 = t41215 ^ t41215;
    wire t41217 = t41216 ^ t41216;
    wire t41218 = t41217 ^ t41217;
    wire t41219 = t41218 ^ t41218;
    wire t41220 = t41219 ^ t41219;
    wire t41221 = t41220 ^ t41220;
    wire t41222 = t41221 ^ t41221;
    wire t41223 = t41222 ^ t41222;
    wire t41224 = t41223 ^ t41223;
    wire t41225 = t41224 ^ t41224;
    wire t41226 = t41225 ^ t41225;
    wire t41227 = t41226 ^ t41226;
    wire t41228 = t41227 ^ t41227;
    wire t41229 = t41228 ^ t41228;
    wire t41230 = t41229 ^ t41229;
    wire t41231 = t41230 ^ t41230;
    wire t41232 = t41231 ^ t41231;
    wire t41233 = t41232 ^ t41232;
    wire t41234 = t41233 ^ t41233;
    wire t41235 = t41234 ^ t41234;
    wire t41236 = t41235 ^ t41235;
    wire t41237 = t41236 ^ t41236;
    wire t41238 = t41237 ^ t41237;
    wire t41239 = t41238 ^ t41238;
    wire t41240 = t41239 ^ t41239;
    wire t41241 = t41240 ^ t41240;
    wire t41242 = t41241 ^ t41241;
    wire t41243 = t41242 ^ t41242;
    wire t41244 = t41243 ^ t41243;
    wire t41245 = t41244 ^ t41244;
    wire t41246 = t41245 ^ t41245;
    wire t41247 = t41246 ^ t41246;
    wire t41248 = t41247 ^ t41247;
    wire t41249 = t41248 ^ t41248;
    wire t41250 = t41249 ^ t41249;
    wire t41251 = t41250 ^ t41250;
    wire t41252 = t41251 ^ t41251;
    wire t41253 = t41252 ^ t41252;
    wire t41254 = t41253 ^ t41253;
    wire t41255 = t41254 ^ t41254;
    wire t41256 = t41255 ^ t41255;
    wire t41257 = t41256 ^ t41256;
    wire t41258 = t41257 ^ t41257;
    wire t41259 = t41258 ^ t41258;
    wire t41260 = t41259 ^ t41259;
    wire t41261 = t41260 ^ t41260;
    wire t41262 = t41261 ^ t41261;
    wire t41263 = t41262 ^ t41262;
    wire t41264 = t41263 ^ t41263;
    wire t41265 = t41264 ^ t41264;
    wire t41266 = t41265 ^ t41265;
    wire t41267 = t41266 ^ t41266;
    wire t41268 = t41267 ^ t41267;
    wire t41269 = t41268 ^ t41268;
    wire t41270 = t41269 ^ t41269;
    wire t41271 = t41270 ^ t41270;
    wire t41272 = t41271 ^ t41271;
    wire t41273 = t41272 ^ t41272;
    wire t41274 = t41273 ^ t41273;
    wire t41275 = t41274 ^ t41274;
    wire t41276 = t41275 ^ t41275;
    wire t41277 = t41276 ^ t41276;
    wire t41278 = t41277 ^ t41277;
    wire t41279 = t41278 ^ t41278;
    wire t41280 = t41279 ^ t41279;
    wire t41281 = t41280 ^ t41280;
    wire t41282 = t41281 ^ t41281;
    wire t41283 = t41282 ^ t41282;
    wire t41284 = t41283 ^ t41283;
    wire t41285 = t41284 ^ t41284;
    wire t41286 = t41285 ^ t41285;
    wire t41287 = t41286 ^ t41286;
    wire t41288 = t41287 ^ t41287;
    wire t41289 = t41288 ^ t41288;
    wire t41290 = t41289 ^ t41289;
    wire t41291 = t41290 ^ t41290;
    wire t41292 = t41291 ^ t41291;
    wire t41293 = t41292 ^ t41292;
    wire t41294 = t41293 ^ t41293;
    wire t41295 = t41294 ^ t41294;
    wire t41296 = t41295 ^ t41295;
    wire t41297 = t41296 ^ t41296;
    wire t41298 = t41297 ^ t41297;
    wire t41299 = t41298 ^ t41298;
    wire t41300 = t41299 ^ t41299;
    wire t41301 = t41300 ^ t41300;
    wire t41302 = t41301 ^ t41301;
    wire t41303 = t41302 ^ t41302;
    wire t41304 = t41303 ^ t41303;
    wire t41305 = t41304 ^ t41304;
    wire t41306 = t41305 ^ t41305;
    wire t41307 = t41306 ^ t41306;
    wire t41308 = t41307 ^ t41307;
    wire t41309 = t41308 ^ t41308;
    wire t41310 = t41309 ^ t41309;
    wire t41311 = t41310 ^ t41310;
    wire t41312 = t41311 ^ t41311;
    wire t41313 = t41312 ^ t41312;
    wire t41314 = t41313 ^ t41313;
    wire t41315 = t41314 ^ t41314;
    wire t41316 = t41315 ^ t41315;
    wire t41317 = t41316 ^ t41316;
    wire t41318 = t41317 ^ t41317;
    wire t41319 = t41318 ^ t41318;
    wire t41320 = t41319 ^ t41319;
    wire t41321 = t41320 ^ t41320;
    wire t41322 = t41321 ^ t41321;
    wire t41323 = t41322 ^ t41322;
    wire t41324 = t41323 ^ t41323;
    wire t41325 = t41324 ^ t41324;
    wire t41326 = t41325 ^ t41325;
    wire t41327 = t41326 ^ t41326;
    wire t41328 = t41327 ^ t41327;
    wire t41329 = t41328 ^ t41328;
    wire t41330 = t41329 ^ t41329;
    wire t41331 = t41330 ^ t41330;
    wire t41332 = t41331 ^ t41331;
    wire t41333 = t41332 ^ t41332;
    wire t41334 = t41333 ^ t41333;
    wire t41335 = t41334 ^ t41334;
    wire t41336 = t41335 ^ t41335;
    wire t41337 = t41336 ^ t41336;
    wire t41338 = t41337 ^ t41337;
    wire t41339 = t41338 ^ t41338;
    wire t41340 = t41339 ^ t41339;
    wire t41341 = t41340 ^ t41340;
    wire t41342 = t41341 ^ t41341;
    wire t41343 = t41342 ^ t41342;
    wire t41344 = t41343 ^ t41343;
    wire t41345 = t41344 ^ t41344;
    wire t41346 = t41345 ^ t41345;
    wire t41347 = t41346 ^ t41346;
    wire t41348 = t41347 ^ t41347;
    wire t41349 = t41348 ^ t41348;
    wire t41350 = t41349 ^ t41349;
    wire t41351 = t41350 ^ t41350;
    wire t41352 = t41351 ^ t41351;
    wire t41353 = t41352 ^ t41352;
    wire t41354 = t41353 ^ t41353;
    wire t41355 = t41354 ^ t41354;
    wire t41356 = t41355 ^ t41355;
    wire t41357 = t41356 ^ t41356;
    wire t41358 = t41357 ^ t41357;
    wire t41359 = t41358 ^ t41358;
    wire t41360 = t41359 ^ t41359;
    wire t41361 = t41360 ^ t41360;
    wire t41362 = t41361 ^ t41361;
    wire t41363 = t41362 ^ t41362;
    wire t41364 = t41363 ^ t41363;
    wire t41365 = t41364 ^ t41364;
    wire t41366 = t41365 ^ t41365;
    wire t41367 = t41366 ^ t41366;
    wire t41368 = t41367 ^ t41367;
    wire t41369 = t41368 ^ t41368;
    wire t41370 = t41369 ^ t41369;
    wire t41371 = t41370 ^ t41370;
    wire t41372 = t41371 ^ t41371;
    wire t41373 = t41372 ^ t41372;
    wire t41374 = t41373 ^ t41373;
    wire t41375 = t41374 ^ t41374;
    wire t41376 = t41375 ^ t41375;
    wire t41377 = t41376 ^ t41376;
    wire t41378 = t41377 ^ t41377;
    wire t41379 = t41378 ^ t41378;
    wire t41380 = t41379 ^ t41379;
    wire t41381 = t41380 ^ t41380;
    wire t41382 = t41381 ^ t41381;
    wire t41383 = t41382 ^ t41382;
    wire t41384 = t41383 ^ t41383;
    wire t41385 = t41384 ^ t41384;
    wire t41386 = t41385 ^ t41385;
    wire t41387 = t41386 ^ t41386;
    wire t41388 = t41387 ^ t41387;
    wire t41389 = t41388 ^ t41388;
    wire t41390 = t41389 ^ t41389;
    wire t41391 = t41390 ^ t41390;
    wire t41392 = t41391 ^ t41391;
    wire t41393 = t41392 ^ t41392;
    wire t41394 = t41393 ^ t41393;
    wire t41395 = t41394 ^ t41394;
    wire t41396 = t41395 ^ t41395;
    wire t41397 = t41396 ^ t41396;
    wire t41398 = t41397 ^ t41397;
    wire t41399 = t41398 ^ t41398;
    wire t41400 = t41399 ^ t41399;
    wire t41401 = t41400 ^ t41400;
    wire t41402 = t41401 ^ t41401;
    wire t41403 = t41402 ^ t41402;
    wire t41404 = t41403 ^ t41403;
    wire t41405 = t41404 ^ t41404;
    wire t41406 = t41405 ^ t41405;
    wire t41407 = t41406 ^ t41406;
    wire t41408 = t41407 ^ t41407;
    wire t41409 = t41408 ^ t41408;
    wire t41410 = t41409 ^ t41409;
    wire t41411 = t41410 ^ t41410;
    wire t41412 = t41411 ^ t41411;
    wire t41413 = t41412 ^ t41412;
    wire t41414 = t41413 ^ t41413;
    wire t41415 = t41414 ^ t41414;
    wire t41416 = t41415 ^ t41415;
    wire t41417 = t41416 ^ t41416;
    wire t41418 = t41417 ^ t41417;
    wire t41419 = t41418 ^ t41418;
    wire t41420 = t41419 ^ t41419;
    wire t41421 = t41420 ^ t41420;
    wire t41422 = t41421 ^ t41421;
    wire t41423 = t41422 ^ t41422;
    wire t41424 = t41423 ^ t41423;
    wire t41425 = t41424 ^ t41424;
    wire t41426 = t41425 ^ t41425;
    wire t41427 = t41426 ^ t41426;
    wire t41428 = t41427 ^ t41427;
    wire t41429 = t41428 ^ t41428;
    wire t41430 = t41429 ^ t41429;
    wire t41431 = t41430 ^ t41430;
    wire t41432 = t41431 ^ t41431;
    wire t41433 = t41432 ^ t41432;
    wire t41434 = t41433 ^ t41433;
    wire t41435 = t41434 ^ t41434;
    wire t41436 = t41435 ^ t41435;
    wire t41437 = t41436 ^ t41436;
    wire t41438 = t41437 ^ t41437;
    wire t41439 = t41438 ^ t41438;
    wire t41440 = t41439 ^ t41439;
    wire t41441 = t41440 ^ t41440;
    wire t41442 = t41441 ^ t41441;
    wire t41443 = t41442 ^ t41442;
    wire t41444 = t41443 ^ t41443;
    wire t41445 = t41444 ^ t41444;
    wire t41446 = t41445 ^ t41445;
    wire t41447 = t41446 ^ t41446;
    wire t41448 = t41447 ^ t41447;
    wire t41449 = t41448 ^ t41448;
    wire t41450 = t41449 ^ t41449;
    wire t41451 = t41450 ^ t41450;
    wire t41452 = t41451 ^ t41451;
    wire t41453 = t41452 ^ t41452;
    wire t41454 = t41453 ^ t41453;
    wire t41455 = t41454 ^ t41454;
    wire t41456 = t41455 ^ t41455;
    wire t41457 = t41456 ^ t41456;
    wire t41458 = t41457 ^ t41457;
    wire t41459 = t41458 ^ t41458;
    wire t41460 = t41459 ^ t41459;
    wire t41461 = t41460 ^ t41460;
    wire t41462 = t41461 ^ t41461;
    wire t41463 = t41462 ^ t41462;
    wire t41464 = t41463 ^ t41463;
    wire t41465 = t41464 ^ t41464;
    wire t41466 = t41465 ^ t41465;
    wire t41467 = t41466 ^ t41466;
    wire t41468 = t41467 ^ t41467;
    wire t41469 = t41468 ^ t41468;
    wire t41470 = t41469 ^ t41469;
    wire t41471 = t41470 ^ t41470;
    wire t41472 = t41471 ^ t41471;
    wire t41473 = t41472 ^ t41472;
    wire t41474 = t41473 ^ t41473;
    wire t41475 = t41474 ^ t41474;
    wire t41476 = t41475 ^ t41475;
    wire t41477 = t41476 ^ t41476;
    wire t41478 = t41477 ^ t41477;
    wire t41479 = t41478 ^ t41478;
    wire t41480 = t41479 ^ t41479;
    wire t41481 = t41480 ^ t41480;
    wire t41482 = t41481 ^ t41481;
    wire t41483 = t41482 ^ t41482;
    wire t41484 = t41483 ^ t41483;
    wire t41485 = t41484 ^ t41484;
    wire t41486 = t41485 ^ t41485;
    wire t41487 = t41486 ^ t41486;
    wire t41488 = t41487 ^ t41487;
    wire t41489 = t41488 ^ t41488;
    wire t41490 = t41489 ^ t41489;
    wire t41491 = t41490 ^ t41490;
    wire t41492 = t41491 ^ t41491;
    wire t41493 = t41492 ^ t41492;
    wire t41494 = t41493 ^ t41493;
    wire t41495 = t41494 ^ t41494;
    wire t41496 = t41495 ^ t41495;
    wire t41497 = t41496 ^ t41496;
    wire t41498 = t41497 ^ t41497;
    wire t41499 = t41498 ^ t41498;
    wire t41500 = t41499 ^ t41499;
    wire t41501 = t41500 ^ t41500;
    wire t41502 = t41501 ^ t41501;
    wire t41503 = t41502 ^ t41502;
    wire t41504 = t41503 ^ t41503;
    wire t41505 = t41504 ^ t41504;
    wire t41506 = t41505 ^ t41505;
    wire t41507 = t41506 ^ t41506;
    wire t41508 = t41507 ^ t41507;
    wire t41509 = t41508 ^ t41508;
    wire t41510 = t41509 ^ t41509;
    wire t41511 = t41510 ^ t41510;
    wire t41512 = t41511 ^ t41511;
    wire t41513 = t41512 ^ t41512;
    wire t41514 = t41513 ^ t41513;
    wire t41515 = t41514 ^ t41514;
    wire t41516 = t41515 ^ t41515;
    wire t41517 = t41516 ^ t41516;
    wire t41518 = t41517 ^ t41517;
    wire t41519 = t41518 ^ t41518;
    wire t41520 = t41519 ^ t41519;
    wire t41521 = t41520 ^ t41520;
    wire t41522 = t41521 ^ t41521;
    wire t41523 = t41522 ^ t41522;
    wire t41524 = t41523 ^ t41523;
    wire t41525 = t41524 ^ t41524;
    wire t41526 = t41525 ^ t41525;
    wire t41527 = t41526 ^ t41526;
    wire t41528 = t41527 ^ t41527;
    wire t41529 = t41528 ^ t41528;
    wire t41530 = t41529 ^ t41529;
    wire t41531 = t41530 ^ t41530;
    wire t41532 = t41531 ^ t41531;
    wire t41533 = t41532 ^ t41532;
    wire t41534 = t41533 ^ t41533;
    wire t41535 = t41534 ^ t41534;
    wire t41536 = t41535 ^ t41535;
    wire t41537 = t41536 ^ t41536;
    wire t41538 = t41537 ^ t41537;
    wire t41539 = t41538 ^ t41538;
    wire t41540 = t41539 ^ t41539;
    wire t41541 = t41540 ^ t41540;
    wire t41542 = t41541 ^ t41541;
    wire t41543 = t41542 ^ t41542;
    wire t41544 = t41543 ^ t41543;
    wire t41545 = t41544 ^ t41544;
    wire t41546 = t41545 ^ t41545;
    wire t41547 = t41546 ^ t41546;
    wire t41548 = t41547 ^ t41547;
    wire t41549 = t41548 ^ t41548;
    wire t41550 = t41549 ^ t41549;
    wire t41551 = t41550 ^ t41550;
    wire t41552 = t41551 ^ t41551;
    wire t41553 = t41552 ^ t41552;
    wire t41554 = t41553 ^ t41553;
    wire t41555 = t41554 ^ t41554;
    wire t41556 = t41555 ^ t41555;
    wire t41557 = t41556 ^ t41556;
    wire t41558 = t41557 ^ t41557;
    wire t41559 = t41558 ^ t41558;
    wire t41560 = t41559 ^ t41559;
    wire t41561 = t41560 ^ t41560;
    wire t41562 = t41561 ^ t41561;
    wire t41563 = t41562 ^ t41562;
    wire t41564 = t41563 ^ t41563;
    wire t41565 = t41564 ^ t41564;
    wire t41566 = t41565 ^ t41565;
    wire t41567 = t41566 ^ t41566;
    wire t41568 = t41567 ^ t41567;
    wire t41569 = t41568 ^ t41568;
    wire t41570 = t41569 ^ t41569;
    wire t41571 = t41570 ^ t41570;
    wire t41572 = t41571 ^ t41571;
    wire t41573 = t41572 ^ t41572;
    wire t41574 = t41573 ^ t41573;
    wire t41575 = t41574 ^ t41574;
    wire t41576 = t41575 ^ t41575;
    wire t41577 = t41576 ^ t41576;
    wire t41578 = t41577 ^ t41577;
    wire t41579 = t41578 ^ t41578;
    wire t41580 = t41579 ^ t41579;
    wire t41581 = t41580 ^ t41580;
    wire t41582 = t41581 ^ t41581;
    wire t41583 = t41582 ^ t41582;
    wire t41584 = t41583 ^ t41583;
    wire t41585 = t41584 ^ t41584;
    wire t41586 = t41585 ^ t41585;
    wire t41587 = t41586 ^ t41586;
    wire t41588 = t41587 ^ t41587;
    wire t41589 = t41588 ^ t41588;
    wire t41590 = t41589 ^ t41589;
    wire t41591 = t41590 ^ t41590;
    wire t41592 = t41591 ^ t41591;
    wire t41593 = t41592 ^ t41592;
    wire t41594 = t41593 ^ t41593;
    wire t41595 = t41594 ^ t41594;
    wire t41596 = t41595 ^ t41595;
    wire t41597 = t41596 ^ t41596;
    wire t41598 = t41597 ^ t41597;
    wire t41599 = t41598 ^ t41598;
    wire t41600 = t41599 ^ t41599;
    wire t41601 = t41600 ^ t41600;
    wire t41602 = t41601 ^ t41601;
    wire t41603 = t41602 ^ t41602;
    wire t41604 = t41603 ^ t41603;
    wire t41605 = t41604 ^ t41604;
    wire t41606 = t41605 ^ t41605;
    wire t41607 = t41606 ^ t41606;
    wire t41608 = t41607 ^ t41607;
    wire t41609 = t41608 ^ t41608;
    wire t41610 = t41609 ^ t41609;
    wire t41611 = t41610 ^ t41610;
    wire t41612 = t41611 ^ t41611;
    wire t41613 = t41612 ^ t41612;
    wire t41614 = t41613 ^ t41613;
    wire t41615 = t41614 ^ t41614;
    wire t41616 = t41615 ^ t41615;
    wire t41617 = t41616 ^ t41616;
    wire t41618 = t41617 ^ t41617;
    wire t41619 = t41618 ^ t41618;
    wire t41620 = t41619 ^ t41619;
    wire t41621 = t41620 ^ t41620;
    wire t41622 = t41621 ^ t41621;
    wire t41623 = t41622 ^ t41622;
    wire t41624 = t41623 ^ t41623;
    wire t41625 = t41624 ^ t41624;
    wire t41626 = t41625 ^ t41625;
    wire t41627 = t41626 ^ t41626;
    wire t41628 = t41627 ^ t41627;
    wire t41629 = t41628 ^ t41628;
    wire t41630 = t41629 ^ t41629;
    wire t41631 = t41630 ^ t41630;
    wire t41632 = t41631 ^ t41631;
    wire t41633 = t41632 ^ t41632;
    wire t41634 = t41633 ^ t41633;
    wire t41635 = t41634 ^ t41634;
    wire t41636 = t41635 ^ t41635;
    wire t41637 = t41636 ^ t41636;
    wire t41638 = t41637 ^ t41637;
    wire t41639 = t41638 ^ t41638;
    wire t41640 = t41639 ^ t41639;
    wire t41641 = t41640 ^ t41640;
    wire t41642 = t41641 ^ t41641;
    wire t41643 = t41642 ^ t41642;
    wire t41644 = t41643 ^ t41643;
    wire t41645 = t41644 ^ t41644;
    wire t41646 = t41645 ^ t41645;
    wire t41647 = t41646 ^ t41646;
    wire t41648 = t41647 ^ t41647;
    wire t41649 = t41648 ^ t41648;
    wire t41650 = t41649 ^ t41649;
    wire t41651 = t41650 ^ t41650;
    wire t41652 = t41651 ^ t41651;
    wire t41653 = t41652 ^ t41652;
    wire t41654 = t41653 ^ t41653;
    wire t41655 = t41654 ^ t41654;
    wire t41656 = t41655 ^ t41655;
    wire t41657 = t41656 ^ t41656;
    wire t41658 = t41657 ^ t41657;
    wire t41659 = t41658 ^ t41658;
    wire t41660 = t41659 ^ t41659;
    wire t41661 = t41660 ^ t41660;
    wire t41662 = t41661 ^ t41661;
    wire t41663 = t41662 ^ t41662;
    wire t41664 = t41663 ^ t41663;
    wire t41665 = t41664 ^ t41664;
    wire t41666 = t41665 ^ t41665;
    wire t41667 = t41666 ^ t41666;
    wire t41668 = t41667 ^ t41667;
    wire t41669 = t41668 ^ t41668;
    wire t41670 = t41669 ^ t41669;
    wire t41671 = t41670 ^ t41670;
    wire t41672 = t41671 ^ t41671;
    wire t41673 = t41672 ^ t41672;
    wire t41674 = t41673 ^ t41673;
    wire t41675 = t41674 ^ t41674;
    wire t41676 = t41675 ^ t41675;
    wire t41677 = t41676 ^ t41676;
    wire t41678 = t41677 ^ t41677;
    wire t41679 = t41678 ^ t41678;
    wire t41680 = t41679 ^ t41679;
    wire t41681 = t41680 ^ t41680;
    wire t41682 = t41681 ^ t41681;
    wire t41683 = t41682 ^ t41682;
    wire t41684 = t41683 ^ t41683;
    wire t41685 = t41684 ^ t41684;
    wire t41686 = t41685 ^ t41685;
    wire t41687 = t41686 ^ t41686;
    wire t41688 = t41687 ^ t41687;
    wire t41689 = t41688 ^ t41688;
    wire t41690 = t41689 ^ t41689;
    wire t41691 = t41690 ^ t41690;
    wire t41692 = t41691 ^ t41691;
    wire t41693 = t41692 ^ t41692;
    wire t41694 = t41693 ^ t41693;
    wire t41695 = t41694 ^ t41694;
    wire t41696 = t41695 ^ t41695;
    wire t41697 = t41696 ^ t41696;
    wire t41698 = t41697 ^ t41697;
    wire t41699 = t41698 ^ t41698;
    wire t41700 = t41699 ^ t41699;
    wire t41701 = t41700 ^ t41700;
    wire t41702 = t41701 ^ t41701;
    wire t41703 = t41702 ^ t41702;
    wire t41704 = t41703 ^ t41703;
    wire t41705 = t41704 ^ t41704;
    wire t41706 = t41705 ^ t41705;
    wire t41707 = t41706 ^ t41706;
    wire t41708 = t41707 ^ t41707;
    wire t41709 = t41708 ^ t41708;
    wire t41710 = t41709 ^ t41709;
    wire t41711 = t41710 ^ t41710;
    wire t41712 = t41711 ^ t41711;
    wire t41713 = t41712 ^ t41712;
    wire t41714 = t41713 ^ t41713;
    wire t41715 = t41714 ^ t41714;
    wire t41716 = t41715 ^ t41715;
    wire t41717 = t41716 ^ t41716;
    wire t41718 = t41717 ^ t41717;
    wire t41719 = t41718 ^ t41718;
    wire t41720 = t41719 ^ t41719;
    wire t41721 = t41720 ^ t41720;
    wire t41722 = t41721 ^ t41721;
    wire t41723 = t41722 ^ t41722;
    wire t41724 = t41723 ^ t41723;
    wire t41725 = t41724 ^ t41724;
    wire t41726 = t41725 ^ t41725;
    wire t41727 = t41726 ^ t41726;
    wire t41728 = t41727 ^ t41727;
    wire t41729 = t41728 ^ t41728;
    wire t41730 = t41729 ^ t41729;
    wire t41731 = t41730 ^ t41730;
    wire t41732 = t41731 ^ t41731;
    wire t41733 = t41732 ^ t41732;
    wire t41734 = t41733 ^ t41733;
    wire t41735 = t41734 ^ t41734;
    wire t41736 = t41735 ^ t41735;
    wire t41737 = t41736 ^ t41736;
    wire t41738 = t41737 ^ t41737;
    wire t41739 = t41738 ^ t41738;
    wire t41740 = t41739 ^ t41739;
    wire t41741 = t41740 ^ t41740;
    wire t41742 = t41741 ^ t41741;
    wire t41743 = t41742 ^ t41742;
    wire t41744 = t41743 ^ t41743;
    wire t41745 = t41744 ^ t41744;
    wire t41746 = t41745 ^ t41745;
    wire t41747 = t41746 ^ t41746;
    wire t41748 = t41747 ^ t41747;
    wire t41749 = t41748 ^ t41748;
    wire t41750 = t41749 ^ t41749;
    wire t41751 = t41750 ^ t41750;
    wire t41752 = t41751 ^ t41751;
    wire t41753 = t41752 ^ t41752;
    wire t41754 = t41753 ^ t41753;
    wire t41755 = t41754 ^ t41754;
    wire t41756 = t41755 ^ t41755;
    wire t41757 = t41756 ^ t41756;
    wire t41758 = t41757 ^ t41757;
    wire t41759 = t41758 ^ t41758;
    wire t41760 = t41759 ^ t41759;
    wire t41761 = t41760 ^ t41760;
    wire t41762 = t41761 ^ t41761;
    wire t41763 = t41762 ^ t41762;
    wire t41764 = t41763 ^ t41763;
    wire t41765 = t41764 ^ t41764;
    wire t41766 = t41765 ^ t41765;
    wire t41767 = t41766 ^ t41766;
    wire t41768 = t41767 ^ t41767;
    wire t41769 = t41768 ^ t41768;
    wire t41770 = t41769 ^ t41769;
    wire t41771 = t41770 ^ t41770;
    wire t41772 = t41771 ^ t41771;
    wire t41773 = t41772 ^ t41772;
    wire t41774 = t41773 ^ t41773;
    wire t41775 = t41774 ^ t41774;
    wire t41776 = t41775 ^ t41775;
    wire t41777 = t41776 ^ t41776;
    wire t41778 = t41777 ^ t41777;
    wire t41779 = t41778 ^ t41778;
    wire t41780 = t41779 ^ t41779;
    wire t41781 = t41780 ^ t41780;
    wire t41782 = t41781 ^ t41781;
    wire t41783 = t41782 ^ t41782;
    wire t41784 = t41783 ^ t41783;
    wire t41785 = t41784 ^ t41784;
    wire t41786 = t41785 ^ t41785;
    wire t41787 = t41786 ^ t41786;
    wire t41788 = t41787 ^ t41787;
    wire t41789 = t41788 ^ t41788;
    wire t41790 = t41789 ^ t41789;
    wire t41791 = t41790 ^ t41790;
    wire t41792 = t41791 ^ t41791;
    wire t41793 = t41792 ^ t41792;
    wire t41794 = t41793 ^ t41793;
    wire t41795 = t41794 ^ t41794;
    wire t41796 = t41795 ^ t41795;
    wire t41797 = t41796 ^ t41796;
    wire t41798 = t41797 ^ t41797;
    wire t41799 = t41798 ^ t41798;
    wire t41800 = t41799 ^ t41799;
    wire t41801 = t41800 ^ t41800;
    wire t41802 = t41801 ^ t41801;
    wire t41803 = t41802 ^ t41802;
    wire t41804 = t41803 ^ t41803;
    wire t41805 = t41804 ^ t41804;
    wire t41806 = t41805 ^ t41805;
    wire t41807 = t41806 ^ t41806;
    wire t41808 = t41807 ^ t41807;
    wire t41809 = t41808 ^ t41808;
    wire t41810 = t41809 ^ t41809;
    wire t41811 = t41810 ^ t41810;
    wire t41812 = t41811 ^ t41811;
    wire t41813 = t41812 ^ t41812;
    wire t41814 = t41813 ^ t41813;
    wire t41815 = t41814 ^ t41814;
    wire t41816 = t41815 ^ t41815;
    wire t41817 = t41816 ^ t41816;
    wire t41818 = t41817 ^ t41817;
    wire t41819 = t41818 ^ t41818;
    wire t41820 = t41819 ^ t41819;
    wire t41821 = t41820 ^ t41820;
    wire t41822 = t41821 ^ t41821;
    wire t41823 = t41822 ^ t41822;
    wire t41824 = t41823 ^ t41823;
    wire t41825 = t41824 ^ t41824;
    wire t41826 = t41825 ^ t41825;
    wire t41827 = t41826 ^ t41826;
    wire t41828 = t41827 ^ t41827;
    wire t41829 = t41828 ^ t41828;
    wire t41830 = t41829 ^ t41829;
    wire t41831 = t41830 ^ t41830;
    wire t41832 = t41831 ^ t41831;
    wire t41833 = t41832 ^ t41832;
    wire t41834 = t41833 ^ t41833;
    wire t41835 = t41834 ^ t41834;
    wire t41836 = t41835 ^ t41835;
    wire t41837 = t41836 ^ t41836;
    wire t41838 = t41837 ^ t41837;
    wire t41839 = t41838 ^ t41838;
    wire t41840 = t41839 ^ t41839;
    wire t41841 = t41840 ^ t41840;
    wire t41842 = t41841 ^ t41841;
    wire t41843 = t41842 ^ t41842;
    wire t41844 = t41843 ^ t41843;
    wire t41845 = t41844 ^ t41844;
    wire t41846 = t41845 ^ t41845;
    wire t41847 = t41846 ^ t41846;
    wire t41848 = t41847 ^ t41847;
    wire t41849 = t41848 ^ t41848;
    wire t41850 = t41849 ^ t41849;
    wire t41851 = t41850 ^ t41850;
    wire t41852 = t41851 ^ t41851;
    wire t41853 = t41852 ^ t41852;
    wire t41854 = t41853 ^ t41853;
    wire t41855 = t41854 ^ t41854;
    wire t41856 = t41855 ^ t41855;
    wire t41857 = t41856 ^ t41856;
    wire t41858 = t41857 ^ t41857;
    wire t41859 = t41858 ^ t41858;
    wire t41860 = t41859 ^ t41859;
    wire t41861 = t41860 ^ t41860;
    wire t41862 = t41861 ^ t41861;
    wire t41863 = t41862 ^ t41862;
    wire t41864 = t41863 ^ t41863;
    wire t41865 = t41864 ^ t41864;
    wire t41866 = t41865 ^ t41865;
    wire t41867 = t41866 ^ t41866;
    wire t41868 = t41867 ^ t41867;
    wire t41869 = t41868 ^ t41868;
    wire t41870 = t41869 ^ t41869;
    wire t41871 = t41870 ^ t41870;
    wire t41872 = t41871 ^ t41871;
    wire t41873 = t41872 ^ t41872;
    wire t41874 = t41873 ^ t41873;
    wire t41875 = t41874 ^ t41874;
    wire t41876 = t41875 ^ t41875;
    wire t41877 = t41876 ^ t41876;
    wire t41878 = t41877 ^ t41877;
    wire t41879 = t41878 ^ t41878;
    wire t41880 = t41879 ^ t41879;
    wire t41881 = t41880 ^ t41880;
    wire t41882 = t41881 ^ t41881;
    wire t41883 = t41882 ^ t41882;
    wire t41884 = t41883 ^ t41883;
    wire t41885 = t41884 ^ t41884;
    wire t41886 = t41885 ^ t41885;
    wire t41887 = t41886 ^ t41886;
    wire t41888 = t41887 ^ t41887;
    wire t41889 = t41888 ^ t41888;
    wire t41890 = t41889 ^ t41889;
    wire t41891 = t41890 ^ t41890;
    wire t41892 = t41891 ^ t41891;
    wire t41893 = t41892 ^ t41892;
    wire t41894 = t41893 ^ t41893;
    wire t41895 = t41894 ^ t41894;
    wire t41896 = t41895 ^ t41895;
    wire t41897 = t41896 ^ t41896;
    wire t41898 = t41897 ^ t41897;
    wire t41899 = t41898 ^ t41898;
    wire t41900 = t41899 ^ t41899;
    wire t41901 = t41900 ^ t41900;
    wire t41902 = t41901 ^ t41901;
    wire t41903 = t41902 ^ t41902;
    wire t41904 = t41903 ^ t41903;
    wire t41905 = t41904 ^ t41904;
    wire t41906 = t41905 ^ t41905;
    wire t41907 = t41906 ^ t41906;
    wire t41908 = t41907 ^ t41907;
    wire t41909 = t41908 ^ t41908;
    wire t41910 = t41909 ^ t41909;
    wire t41911 = t41910 ^ t41910;
    wire t41912 = t41911 ^ t41911;
    wire t41913 = t41912 ^ t41912;
    wire t41914 = t41913 ^ t41913;
    wire t41915 = t41914 ^ t41914;
    wire t41916 = t41915 ^ t41915;
    wire t41917 = t41916 ^ t41916;
    wire t41918 = t41917 ^ t41917;
    wire t41919 = t41918 ^ t41918;
    wire t41920 = t41919 ^ t41919;
    wire t41921 = t41920 ^ t41920;
    wire t41922 = t41921 ^ t41921;
    wire t41923 = t41922 ^ t41922;
    wire t41924 = t41923 ^ t41923;
    wire t41925 = t41924 ^ t41924;
    wire t41926 = t41925 ^ t41925;
    wire t41927 = t41926 ^ t41926;
    wire t41928 = t41927 ^ t41927;
    wire t41929 = t41928 ^ t41928;
    wire t41930 = t41929 ^ t41929;
    wire t41931 = t41930 ^ t41930;
    wire t41932 = t41931 ^ t41931;
    wire t41933 = t41932 ^ t41932;
    wire t41934 = t41933 ^ t41933;
    wire t41935 = t41934 ^ t41934;
    wire t41936 = t41935 ^ t41935;
    wire t41937 = t41936 ^ t41936;
    wire t41938 = t41937 ^ t41937;
    wire t41939 = t41938 ^ t41938;
    wire t41940 = t41939 ^ t41939;
    wire t41941 = t41940 ^ t41940;
    wire t41942 = t41941 ^ t41941;
    wire t41943 = t41942 ^ t41942;
    wire t41944 = t41943 ^ t41943;
    wire t41945 = t41944 ^ t41944;
    wire t41946 = t41945 ^ t41945;
    wire t41947 = t41946 ^ t41946;
    wire t41948 = t41947 ^ t41947;
    wire t41949 = t41948 ^ t41948;
    wire t41950 = t41949 ^ t41949;
    wire t41951 = t41950 ^ t41950;
    wire t41952 = t41951 ^ t41951;
    wire t41953 = t41952 ^ t41952;
    wire t41954 = t41953 ^ t41953;
    wire t41955 = t41954 ^ t41954;
    wire t41956 = t41955 ^ t41955;
    wire t41957 = t41956 ^ t41956;
    wire t41958 = t41957 ^ t41957;
    wire t41959 = t41958 ^ t41958;
    wire t41960 = t41959 ^ t41959;
    wire t41961 = t41960 ^ t41960;
    wire t41962 = t41961 ^ t41961;
    wire t41963 = t41962 ^ t41962;
    wire t41964 = t41963 ^ t41963;
    wire t41965 = t41964 ^ t41964;
    wire t41966 = t41965 ^ t41965;
    wire t41967 = t41966 ^ t41966;
    wire t41968 = t41967 ^ t41967;
    wire t41969 = t41968 ^ t41968;
    wire t41970 = t41969 ^ t41969;
    wire t41971 = t41970 ^ t41970;
    wire t41972 = t41971 ^ t41971;
    wire t41973 = t41972 ^ t41972;
    wire t41974 = t41973 ^ t41973;
    wire t41975 = t41974 ^ t41974;
    wire t41976 = t41975 ^ t41975;
    wire t41977 = t41976 ^ t41976;
    wire t41978 = t41977 ^ t41977;
    wire t41979 = t41978 ^ t41978;
    wire t41980 = t41979 ^ t41979;
    wire t41981 = t41980 ^ t41980;
    wire t41982 = t41981 ^ t41981;
    wire t41983 = t41982 ^ t41982;
    wire t41984 = t41983 ^ t41983;
    wire t41985 = t41984 ^ t41984;
    wire t41986 = t41985 ^ t41985;
    wire t41987 = t41986 ^ t41986;
    wire t41988 = t41987 ^ t41987;
    wire t41989 = t41988 ^ t41988;
    wire t41990 = t41989 ^ t41989;
    wire t41991 = t41990 ^ t41990;
    wire t41992 = t41991 ^ t41991;
    wire t41993 = t41992 ^ t41992;
    wire t41994 = t41993 ^ t41993;
    wire t41995 = t41994 ^ t41994;
    wire t41996 = t41995 ^ t41995;
    wire t41997 = t41996 ^ t41996;
    wire t41998 = t41997 ^ t41997;
    wire t41999 = t41998 ^ t41998;
    wire t42000 = t41999 ^ t41999;
    wire t42001 = t42000 ^ t42000;
    wire t42002 = t42001 ^ t42001;
    wire t42003 = t42002 ^ t42002;
    wire t42004 = t42003 ^ t42003;
    wire t42005 = t42004 ^ t42004;
    wire t42006 = t42005 ^ t42005;
    wire t42007 = t42006 ^ t42006;
    wire t42008 = t42007 ^ t42007;
    wire t42009 = t42008 ^ t42008;
    wire t42010 = t42009 ^ t42009;
    wire t42011 = t42010 ^ t42010;
    wire t42012 = t42011 ^ t42011;
    wire t42013 = t42012 ^ t42012;
    wire t42014 = t42013 ^ t42013;
    wire t42015 = t42014 ^ t42014;
    wire t42016 = t42015 ^ t42015;
    wire t42017 = t42016 ^ t42016;
    wire t42018 = t42017 ^ t42017;
    wire t42019 = t42018 ^ t42018;
    wire t42020 = t42019 ^ t42019;
    wire t42021 = t42020 ^ t42020;
    wire t42022 = t42021 ^ t42021;
    wire t42023 = t42022 ^ t42022;
    wire t42024 = t42023 ^ t42023;
    wire t42025 = t42024 ^ t42024;
    wire t42026 = t42025 ^ t42025;
    wire t42027 = t42026 ^ t42026;
    wire t42028 = t42027 ^ t42027;
    wire t42029 = t42028 ^ t42028;
    wire t42030 = t42029 ^ t42029;
    wire t42031 = t42030 ^ t42030;
    wire t42032 = t42031 ^ t42031;
    wire t42033 = t42032 ^ t42032;
    wire t42034 = t42033 ^ t42033;
    wire t42035 = t42034 ^ t42034;
    wire t42036 = t42035 ^ t42035;
    wire t42037 = t42036 ^ t42036;
    wire t42038 = t42037 ^ t42037;
    wire t42039 = t42038 ^ t42038;
    wire t42040 = t42039 ^ t42039;
    wire t42041 = t42040 ^ t42040;
    wire t42042 = t42041 ^ t42041;
    wire t42043 = t42042 ^ t42042;
    wire t42044 = t42043 ^ t42043;
    wire t42045 = t42044 ^ t42044;
    wire t42046 = t42045 ^ t42045;
    wire t42047 = t42046 ^ t42046;
    wire t42048 = t42047 ^ t42047;
    wire t42049 = t42048 ^ t42048;
    wire t42050 = t42049 ^ t42049;
    wire t42051 = t42050 ^ t42050;
    wire t42052 = t42051 ^ t42051;
    wire t42053 = t42052 ^ t42052;
    wire t42054 = t42053 ^ t42053;
    wire t42055 = t42054 ^ t42054;
    wire t42056 = t42055 ^ t42055;
    wire t42057 = t42056 ^ t42056;
    wire t42058 = t42057 ^ t42057;
    wire t42059 = t42058 ^ t42058;
    wire t42060 = t42059 ^ t42059;
    wire t42061 = t42060 ^ t42060;
    wire t42062 = t42061 ^ t42061;
    wire t42063 = t42062 ^ t42062;
    wire t42064 = t42063 ^ t42063;
    wire t42065 = t42064 ^ t42064;
    wire t42066 = t42065 ^ t42065;
    wire t42067 = t42066 ^ t42066;
    wire t42068 = t42067 ^ t42067;
    wire t42069 = t42068 ^ t42068;
    wire t42070 = t42069 ^ t42069;
    wire t42071 = t42070 ^ t42070;
    wire t42072 = t42071 ^ t42071;
    wire t42073 = t42072 ^ t42072;
    wire t42074 = t42073 ^ t42073;
    wire t42075 = t42074 ^ t42074;
    wire t42076 = t42075 ^ t42075;
    wire t42077 = t42076 ^ t42076;
    wire t42078 = t42077 ^ t42077;
    wire t42079 = t42078 ^ t42078;
    wire t42080 = t42079 ^ t42079;
    wire t42081 = t42080 ^ t42080;
    wire t42082 = t42081 ^ t42081;
    wire t42083 = t42082 ^ t42082;
    wire t42084 = t42083 ^ t42083;
    wire t42085 = t42084 ^ t42084;
    wire t42086 = t42085 ^ t42085;
    wire t42087 = t42086 ^ t42086;
    wire t42088 = t42087 ^ t42087;
    wire t42089 = t42088 ^ t42088;
    wire t42090 = t42089 ^ t42089;
    wire t42091 = t42090 ^ t42090;
    wire t42092 = t42091 ^ t42091;
    wire t42093 = t42092 ^ t42092;
    wire t42094 = t42093 ^ t42093;
    wire t42095 = t42094 ^ t42094;
    wire t42096 = t42095 ^ t42095;
    wire t42097 = t42096 ^ t42096;
    wire t42098 = t42097 ^ t42097;
    wire t42099 = t42098 ^ t42098;
    wire t42100 = t42099 ^ t42099;
    wire t42101 = t42100 ^ t42100;
    wire t42102 = t42101 ^ t42101;
    wire t42103 = t42102 ^ t42102;
    wire t42104 = t42103 ^ t42103;
    wire t42105 = t42104 ^ t42104;
    wire t42106 = t42105 ^ t42105;
    wire t42107 = t42106 ^ t42106;
    wire t42108 = t42107 ^ t42107;
    wire t42109 = t42108 ^ t42108;
    wire t42110 = t42109 ^ t42109;
    wire t42111 = t42110 ^ t42110;
    wire t42112 = t42111 ^ t42111;
    wire t42113 = t42112 ^ t42112;
    wire t42114 = t42113 ^ t42113;
    wire t42115 = t42114 ^ t42114;
    wire t42116 = t42115 ^ t42115;
    wire t42117 = t42116 ^ t42116;
    wire t42118 = t42117 ^ t42117;
    wire t42119 = t42118 ^ t42118;
    wire t42120 = t42119 ^ t42119;
    wire t42121 = t42120 ^ t42120;
    wire t42122 = t42121 ^ t42121;
    wire t42123 = t42122 ^ t42122;
    wire t42124 = t42123 ^ t42123;
    wire t42125 = t42124 ^ t42124;
    wire t42126 = t42125 ^ t42125;
    wire t42127 = t42126 ^ t42126;
    wire t42128 = t42127 ^ t42127;
    wire t42129 = t42128 ^ t42128;
    wire t42130 = t42129 ^ t42129;
    wire t42131 = t42130 ^ t42130;
    wire t42132 = t42131 ^ t42131;
    wire t42133 = t42132 ^ t42132;
    wire t42134 = t42133 ^ t42133;
    wire t42135 = t42134 ^ t42134;
    wire t42136 = t42135 ^ t42135;
    wire t42137 = t42136 ^ t42136;
    wire t42138 = t42137 ^ t42137;
    wire t42139 = t42138 ^ t42138;
    wire t42140 = t42139 ^ t42139;
    wire t42141 = t42140 ^ t42140;
    wire t42142 = t42141 ^ t42141;
    wire t42143 = t42142 ^ t42142;
    wire t42144 = t42143 ^ t42143;
    wire t42145 = t42144 ^ t42144;
    wire t42146 = t42145 ^ t42145;
    wire t42147 = t42146 ^ t42146;
    wire t42148 = t42147 ^ t42147;
    wire t42149 = t42148 ^ t42148;
    wire t42150 = t42149 ^ t42149;
    wire t42151 = t42150 ^ t42150;
    wire t42152 = t42151 ^ t42151;
    wire t42153 = t42152 ^ t42152;
    wire t42154 = t42153 ^ t42153;
    wire t42155 = t42154 ^ t42154;
    wire t42156 = t42155 ^ t42155;
    wire t42157 = t42156 ^ t42156;
    wire t42158 = t42157 ^ t42157;
    wire t42159 = t42158 ^ t42158;
    wire t42160 = t42159 ^ t42159;
    wire t42161 = t42160 ^ t42160;
    wire t42162 = t42161 ^ t42161;
    wire t42163 = t42162 ^ t42162;
    wire t42164 = t42163 ^ t42163;
    wire t42165 = t42164 ^ t42164;
    wire t42166 = t42165 ^ t42165;
    wire t42167 = t42166 ^ t42166;
    wire t42168 = t42167 ^ t42167;
    wire t42169 = t42168 ^ t42168;
    wire t42170 = t42169 ^ t42169;
    wire t42171 = t42170 ^ t42170;
    wire t42172 = t42171 ^ t42171;
    wire t42173 = t42172 ^ t42172;
    wire t42174 = t42173 ^ t42173;
    wire t42175 = t42174 ^ t42174;
    wire t42176 = t42175 ^ t42175;
    wire t42177 = t42176 ^ t42176;
    wire t42178 = t42177 ^ t42177;
    wire t42179 = t42178 ^ t42178;
    wire t42180 = t42179 ^ t42179;
    wire t42181 = t42180 ^ t42180;
    wire t42182 = t42181 ^ t42181;
    wire t42183 = t42182 ^ t42182;
    wire t42184 = t42183 ^ t42183;
    wire t42185 = t42184 ^ t42184;
    wire t42186 = t42185 ^ t42185;
    wire t42187 = t42186 ^ t42186;
    wire t42188 = t42187 ^ t42187;
    wire t42189 = t42188 ^ t42188;
    wire t42190 = t42189 ^ t42189;
    wire t42191 = t42190 ^ t42190;
    wire t42192 = t42191 ^ t42191;
    wire t42193 = t42192 ^ t42192;
    wire t42194 = t42193 ^ t42193;
    wire t42195 = t42194 ^ t42194;
    wire t42196 = t42195 ^ t42195;
    wire t42197 = t42196 ^ t42196;
    wire t42198 = t42197 ^ t42197;
    wire t42199 = t42198 ^ t42198;
    wire t42200 = t42199 ^ t42199;
    wire t42201 = t42200 ^ t42200;
    wire t42202 = t42201 ^ t42201;
    wire t42203 = t42202 ^ t42202;
    wire t42204 = t42203 ^ t42203;
    wire t42205 = t42204 ^ t42204;
    wire t42206 = t42205 ^ t42205;
    wire t42207 = t42206 ^ t42206;
    wire t42208 = t42207 ^ t42207;
    wire t42209 = t42208 ^ t42208;
    wire t42210 = t42209 ^ t42209;
    wire t42211 = t42210 ^ t42210;
    wire t42212 = t42211 ^ t42211;
    wire t42213 = t42212 ^ t42212;
    wire t42214 = t42213 ^ t42213;
    wire t42215 = t42214 ^ t42214;
    wire t42216 = t42215 ^ t42215;
    wire t42217 = t42216 ^ t42216;
    wire t42218 = t42217 ^ t42217;
    wire t42219 = t42218 ^ t42218;
    wire t42220 = t42219 ^ t42219;
    wire t42221 = t42220 ^ t42220;
    wire t42222 = t42221 ^ t42221;
    wire t42223 = t42222 ^ t42222;
    wire t42224 = t42223 ^ t42223;
    wire t42225 = t42224 ^ t42224;
    wire t42226 = t42225 ^ t42225;
    wire t42227 = t42226 ^ t42226;
    wire t42228 = t42227 ^ t42227;
    wire t42229 = t42228 ^ t42228;
    wire t42230 = t42229 ^ t42229;
    wire t42231 = t42230 ^ t42230;
    wire t42232 = t42231 ^ t42231;
    wire t42233 = t42232 ^ t42232;
    wire t42234 = t42233 ^ t42233;
    wire t42235 = t42234 ^ t42234;
    wire t42236 = t42235 ^ t42235;
    wire t42237 = t42236 ^ t42236;
    wire t42238 = t42237 ^ t42237;
    wire t42239 = t42238 ^ t42238;
    wire t42240 = t42239 ^ t42239;
    wire t42241 = t42240 ^ t42240;
    wire t42242 = t42241 ^ t42241;
    wire t42243 = t42242 ^ t42242;
    wire t42244 = t42243 ^ t42243;
    wire t42245 = t42244 ^ t42244;
    wire t42246 = t42245 ^ t42245;
    wire t42247 = t42246 ^ t42246;
    wire t42248 = t42247 ^ t42247;
    wire t42249 = t42248 ^ t42248;
    wire t42250 = t42249 ^ t42249;
    wire t42251 = t42250 ^ t42250;
    wire t42252 = t42251 ^ t42251;
    wire t42253 = t42252 ^ t42252;
    wire t42254 = t42253 ^ t42253;
    wire t42255 = t42254 ^ t42254;
    wire t42256 = t42255 ^ t42255;
    wire t42257 = t42256 ^ t42256;
    wire t42258 = t42257 ^ t42257;
    wire t42259 = t42258 ^ t42258;
    wire t42260 = t42259 ^ t42259;
    wire t42261 = t42260 ^ t42260;
    wire t42262 = t42261 ^ t42261;
    wire t42263 = t42262 ^ t42262;
    wire t42264 = t42263 ^ t42263;
    wire t42265 = t42264 ^ t42264;
    wire t42266 = t42265 ^ t42265;
    wire t42267 = t42266 ^ t42266;
    wire t42268 = t42267 ^ t42267;
    wire t42269 = t42268 ^ t42268;
    wire t42270 = t42269 ^ t42269;
    wire t42271 = t42270 ^ t42270;
    wire t42272 = t42271 ^ t42271;
    wire t42273 = t42272 ^ t42272;
    wire t42274 = t42273 ^ t42273;
    wire t42275 = t42274 ^ t42274;
    wire t42276 = t42275 ^ t42275;
    wire t42277 = t42276 ^ t42276;
    wire t42278 = t42277 ^ t42277;
    wire t42279 = t42278 ^ t42278;
    wire t42280 = t42279 ^ t42279;
    wire t42281 = t42280 ^ t42280;
    wire t42282 = t42281 ^ t42281;
    wire t42283 = t42282 ^ t42282;
    wire t42284 = t42283 ^ t42283;
    wire t42285 = t42284 ^ t42284;
    wire t42286 = t42285 ^ t42285;
    wire t42287 = t42286 ^ t42286;
    wire t42288 = t42287 ^ t42287;
    wire t42289 = t42288 ^ t42288;
    wire t42290 = t42289 ^ t42289;
    wire t42291 = t42290 ^ t42290;
    wire t42292 = t42291 ^ t42291;
    wire t42293 = t42292 ^ t42292;
    wire t42294 = t42293 ^ t42293;
    wire t42295 = t42294 ^ t42294;
    wire t42296 = t42295 ^ t42295;
    wire t42297 = t42296 ^ t42296;
    wire t42298 = t42297 ^ t42297;
    wire t42299 = t42298 ^ t42298;
    wire t42300 = t42299 ^ t42299;
    wire t42301 = t42300 ^ t42300;
    wire t42302 = t42301 ^ t42301;
    wire t42303 = t42302 ^ t42302;
    wire t42304 = t42303 ^ t42303;
    wire t42305 = t42304 ^ t42304;
    wire t42306 = t42305 ^ t42305;
    wire t42307 = t42306 ^ t42306;
    wire t42308 = t42307 ^ t42307;
    wire t42309 = t42308 ^ t42308;
    wire t42310 = t42309 ^ t42309;
    wire t42311 = t42310 ^ t42310;
    wire t42312 = t42311 ^ t42311;
    wire t42313 = t42312 ^ t42312;
    wire t42314 = t42313 ^ t42313;
    wire t42315 = t42314 ^ t42314;
    wire t42316 = t42315 ^ t42315;
    wire t42317 = t42316 ^ t42316;
    wire t42318 = t42317 ^ t42317;
    wire t42319 = t42318 ^ t42318;
    wire t42320 = t42319 ^ t42319;
    wire t42321 = t42320 ^ t42320;
    wire t42322 = t42321 ^ t42321;
    wire t42323 = t42322 ^ t42322;
    wire t42324 = t42323 ^ t42323;
    wire t42325 = t42324 ^ t42324;
    wire t42326 = t42325 ^ t42325;
    wire t42327 = t42326 ^ t42326;
    wire t42328 = t42327 ^ t42327;
    wire t42329 = t42328 ^ t42328;
    wire t42330 = t42329 ^ t42329;
    wire t42331 = t42330 ^ t42330;
    wire t42332 = t42331 ^ t42331;
    wire t42333 = t42332 ^ t42332;
    wire t42334 = t42333 ^ t42333;
    wire t42335 = t42334 ^ t42334;
    wire t42336 = t42335 ^ t42335;
    wire t42337 = t42336 ^ t42336;
    wire t42338 = t42337 ^ t42337;
    wire t42339 = t42338 ^ t42338;
    wire t42340 = t42339 ^ t42339;
    wire t42341 = t42340 ^ t42340;
    wire t42342 = t42341 ^ t42341;
    wire t42343 = t42342 ^ t42342;
    wire t42344 = t42343 ^ t42343;
    wire t42345 = t42344 ^ t42344;
    wire t42346 = t42345 ^ t42345;
    wire t42347 = t42346 ^ t42346;
    wire t42348 = t42347 ^ t42347;
    wire t42349 = t42348 ^ t42348;
    wire t42350 = t42349 ^ t42349;
    wire t42351 = t42350 ^ t42350;
    wire t42352 = t42351 ^ t42351;
    wire t42353 = t42352 ^ t42352;
    wire t42354 = t42353 ^ t42353;
    wire t42355 = t42354 ^ t42354;
    wire t42356 = t42355 ^ t42355;
    wire t42357 = t42356 ^ t42356;
    wire t42358 = t42357 ^ t42357;
    wire t42359 = t42358 ^ t42358;
    wire t42360 = t42359 ^ t42359;
    wire t42361 = t42360 ^ t42360;
    wire t42362 = t42361 ^ t42361;
    wire t42363 = t42362 ^ t42362;
    wire t42364 = t42363 ^ t42363;
    wire t42365 = t42364 ^ t42364;
    wire t42366 = t42365 ^ t42365;
    wire t42367 = t42366 ^ t42366;
    wire t42368 = t42367 ^ t42367;
    wire t42369 = t42368 ^ t42368;
    wire t42370 = t42369 ^ t42369;
    wire t42371 = t42370 ^ t42370;
    wire t42372 = t42371 ^ t42371;
    wire t42373 = t42372 ^ t42372;
    wire t42374 = t42373 ^ t42373;
    wire t42375 = t42374 ^ t42374;
    wire t42376 = t42375 ^ t42375;
    wire t42377 = t42376 ^ t42376;
    wire t42378 = t42377 ^ t42377;
    wire t42379 = t42378 ^ t42378;
    wire t42380 = t42379 ^ t42379;
    wire t42381 = t42380 ^ t42380;
    wire t42382 = t42381 ^ t42381;
    wire t42383 = t42382 ^ t42382;
    wire t42384 = t42383 ^ t42383;
    wire t42385 = t42384 ^ t42384;
    wire t42386 = t42385 ^ t42385;
    wire t42387 = t42386 ^ t42386;
    wire t42388 = t42387 ^ t42387;
    wire t42389 = t42388 ^ t42388;
    wire t42390 = t42389 ^ t42389;
    wire t42391 = t42390 ^ t42390;
    wire t42392 = t42391 ^ t42391;
    wire t42393 = t42392 ^ t42392;
    wire t42394 = t42393 ^ t42393;
    wire t42395 = t42394 ^ t42394;
    wire t42396 = t42395 ^ t42395;
    wire t42397 = t42396 ^ t42396;
    wire t42398 = t42397 ^ t42397;
    wire t42399 = t42398 ^ t42398;
    wire t42400 = t42399 ^ t42399;
    wire t42401 = t42400 ^ t42400;
    wire t42402 = t42401 ^ t42401;
    wire t42403 = t42402 ^ t42402;
    wire t42404 = t42403 ^ t42403;
    wire t42405 = t42404 ^ t42404;
    wire t42406 = t42405 ^ t42405;
    wire t42407 = t42406 ^ t42406;
    wire t42408 = t42407 ^ t42407;
    wire t42409 = t42408 ^ t42408;
    wire t42410 = t42409 ^ t42409;
    wire t42411 = t42410 ^ t42410;
    wire t42412 = t42411 ^ t42411;
    wire t42413 = t42412 ^ t42412;
    wire t42414 = t42413 ^ t42413;
    wire t42415 = t42414 ^ t42414;
    wire t42416 = t42415 ^ t42415;
    wire t42417 = t42416 ^ t42416;
    wire t42418 = t42417 ^ t42417;
    wire t42419 = t42418 ^ t42418;
    wire t42420 = t42419 ^ t42419;
    wire t42421 = t42420 ^ t42420;
    wire t42422 = t42421 ^ t42421;
    wire t42423 = t42422 ^ t42422;
    wire t42424 = t42423 ^ t42423;
    wire t42425 = t42424 ^ t42424;
    wire t42426 = t42425 ^ t42425;
    wire t42427 = t42426 ^ t42426;
    wire t42428 = t42427 ^ t42427;
    wire t42429 = t42428 ^ t42428;
    wire t42430 = t42429 ^ t42429;
    wire t42431 = t42430 ^ t42430;
    wire t42432 = t42431 ^ t42431;
    wire t42433 = t42432 ^ t42432;
    wire t42434 = t42433 ^ t42433;
    wire t42435 = t42434 ^ t42434;
    wire t42436 = t42435 ^ t42435;
    wire t42437 = t42436 ^ t42436;
    wire t42438 = t42437 ^ t42437;
    wire t42439 = t42438 ^ t42438;
    wire t42440 = t42439 ^ t42439;
    wire t42441 = t42440 ^ t42440;
    wire t42442 = t42441 ^ t42441;
    wire t42443 = t42442 ^ t42442;
    wire t42444 = t42443 ^ t42443;
    wire t42445 = t42444 ^ t42444;
    wire t42446 = t42445 ^ t42445;
    wire t42447 = t42446 ^ t42446;
    wire t42448 = t42447 ^ t42447;
    wire t42449 = t42448 ^ t42448;
    wire t42450 = t42449 ^ t42449;
    wire t42451 = t42450 ^ t42450;
    wire t42452 = t42451 ^ t42451;
    wire t42453 = t42452 ^ t42452;
    wire t42454 = t42453 ^ t42453;
    wire t42455 = t42454 ^ t42454;
    wire t42456 = t42455 ^ t42455;
    wire t42457 = t42456 ^ t42456;
    wire t42458 = t42457 ^ t42457;
    wire t42459 = t42458 ^ t42458;
    wire t42460 = t42459 ^ t42459;
    wire t42461 = t42460 ^ t42460;
    wire t42462 = t42461 ^ t42461;
    wire t42463 = t42462 ^ t42462;
    wire t42464 = t42463 ^ t42463;
    wire t42465 = t42464 ^ t42464;
    wire t42466 = t42465 ^ t42465;
    wire t42467 = t42466 ^ t42466;
    wire t42468 = t42467 ^ t42467;
    wire t42469 = t42468 ^ t42468;
    wire t42470 = t42469 ^ t42469;
    wire t42471 = t42470 ^ t42470;
    wire t42472 = t42471 ^ t42471;
    wire t42473 = t42472 ^ t42472;
    wire t42474 = t42473 ^ t42473;
    wire t42475 = t42474 ^ t42474;
    wire t42476 = t42475 ^ t42475;
    wire t42477 = t42476 ^ t42476;
    wire t42478 = t42477 ^ t42477;
    wire t42479 = t42478 ^ t42478;
    wire t42480 = t42479 ^ t42479;
    wire t42481 = t42480 ^ t42480;
    wire t42482 = t42481 ^ t42481;
    wire t42483 = t42482 ^ t42482;
    wire t42484 = t42483 ^ t42483;
    wire t42485 = t42484 ^ t42484;
    wire t42486 = t42485 ^ t42485;
    wire t42487 = t42486 ^ t42486;
    wire t42488 = t42487 ^ t42487;
    wire t42489 = t42488 ^ t42488;
    wire t42490 = t42489 ^ t42489;
    wire t42491 = t42490 ^ t42490;
    wire t42492 = t42491 ^ t42491;
    wire t42493 = t42492 ^ t42492;
    wire t42494 = t42493 ^ t42493;
    wire t42495 = t42494 ^ t42494;
    wire t42496 = t42495 ^ t42495;
    wire t42497 = t42496 ^ t42496;
    wire t42498 = t42497 ^ t42497;
    wire t42499 = t42498 ^ t42498;
    wire t42500 = t42499 ^ t42499;
    wire t42501 = t42500 ^ t42500;
    wire t42502 = t42501 ^ t42501;
    wire t42503 = t42502 ^ t42502;
    wire t42504 = t42503 ^ t42503;
    wire t42505 = t42504 ^ t42504;
    wire t42506 = t42505 ^ t42505;
    wire t42507 = t42506 ^ t42506;
    wire t42508 = t42507 ^ t42507;
    wire t42509 = t42508 ^ t42508;
    wire t42510 = t42509 ^ t42509;
    wire t42511 = t42510 ^ t42510;
    wire t42512 = t42511 ^ t42511;
    wire t42513 = t42512 ^ t42512;
    wire t42514 = t42513 ^ t42513;
    wire t42515 = t42514 ^ t42514;
    wire t42516 = t42515 ^ t42515;
    wire t42517 = t42516 ^ t42516;
    wire t42518 = t42517 ^ t42517;
    wire t42519 = t42518 ^ t42518;
    wire t42520 = t42519 ^ t42519;
    wire t42521 = t42520 ^ t42520;
    wire t42522 = t42521 ^ t42521;
    wire t42523 = t42522 ^ t42522;
    wire t42524 = t42523 ^ t42523;
    wire t42525 = t42524 ^ t42524;
    wire t42526 = t42525 ^ t42525;
    wire t42527 = t42526 ^ t42526;
    wire t42528 = t42527 ^ t42527;
    wire t42529 = t42528 ^ t42528;
    wire t42530 = t42529 ^ t42529;
    wire t42531 = t42530 ^ t42530;
    wire t42532 = t42531 ^ t42531;
    wire t42533 = t42532 ^ t42532;
    wire t42534 = t42533 ^ t42533;
    wire t42535 = t42534 ^ t42534;
    wire t42536 = t42535 ^ t42535;
    wire t42537 = t42536 ^ t42536;
    wire t42538 = t42537 ^ t42537;
    wire t42539 = t42538 ^ t42538;
    wire t42540 = t42539 ^ t42539;
    wire t42541 = t42540 ^ t42540;
    wire t42542 = t42541 ^ t42541;
    wire t42543 = t42542 ^ t42542;
    wire t42544 = t42543 ^ t42543;
    wire t42545 = t42544 ^ t42544;
    wire t42546 = t42545 ^ t42545;
    wire t42547 = t42546 ^ t42546;
    wire t42548 = t42547 ^ t42547;
    wire t42549 = t42548 ^ t42548;
    wire t42550 = t42549 ^ t42549;
    wire t42551 = t42550 ^ t42550;
    wire t42552 = t42551 ^ t42551;
    wire t42553 = t42552 ^ t42552;
    wire t42554 = t42553 ^ t42553;
    wire t42555 = t42554 ^ t42554;
    wire t42556 = t42555 ^ t42555;
    wire t42557 = t42556 ^ t42556;
    wire t42558 = t42557 ^ t42557;
    wire t42559 = t42558 ^ t42558;
    wire t42560 = t42559 ^ t42559;
    wire t42561 = t42560 ^ t42560;
    wire t42562 = t42561 ^ t42561;
    wire t42563 = t42562 ^ t42562;
    wire t42564 = t42563 ^ t42563;
    wire t42565 = t42564 ^ t42564;
    wire t42566 = t42565 ^ t42565;
    wire t42567 = t42566 ^ t42566;
    wire t42568 = t42567 ^ t42567;
    wire t42569 = t42568 ^ t42568;
    wire t42570 = t42569 ^ t42569;
    wire t42571 = t42570 ^ t42570;
    wire t42572 = t42571 ^ t42571;
    wire t42573 = t42572 ^ t42572;
    wire t42574 = t42573 ^ t42573;
    wire t42575 = t42574 ^ t42574;
    wire t42576 = t42575 ^ t42575;
    wire t42577 = t42576 ^ t42576;
    wire t42578 = t42577 ^ t42577;
    wire t42579 = t42578 ^ t42578;
    wire t42580 = t42579 ^ t42579;
    wire t42581 = t42580 ^ t42580;
    wire t42582 = t42581 ^ t42581;
    wire t42583 = t42582 ^ t42582;
    wire t42584 = t42583 ^ t42583;
    wire t42585 = t42584 ^ t42584;
    wire t42586 = t42585 ^ t42585;
    wire t42587 = t42586 ^ t42586;
    wire t42588 = t42587 ^ t42587;
    wire t42589 = t42588 ^ t42588;
    wire t42590 = t42589 ^ t42589;
    wire t42591 = t42590 ^ t42590;
    wire t42592 = t42591 ^ t42591;
    wire t42593 = t42592 ^ t42592;
    wire t42594 = t42593 ^ t42593;
    wire t42595 = t42594 ^ t42594;
    wire t42596 = t42595 ^ t42595;
    wire t42597 = t42596 ^ t42596;
    wire t42598 = t42597 ^ t42597;
    wire t42599 = t42598 ^ t42598;
    wire t42600 = t42599 ^ t42599;
    wire t42601 = t42600 ^ t42600;
    wire t42602 = t42601 ^ t42601;
    wire t42603 = t42602 ^ t42602;
    wire t42604 = t42603 ^ t42603;
    wire t42605 = t42604 ^ t42604;
    wire t42606 = t42605 ^ t42605;
    wire t42607 = t42606 ^ t42606;
    wire t42608 = t42607 ^ t42607;
    wire t42609 = t42608 ^ t42608;
    wire t42610 = t42609 ^ t42609;
    wire t42611 = t42610 ^ t42610;
    wire t42612 = t42611 ^ t42611;
    wire t42613 = t42612 ^ t42612;
    wire t42614 = t42613 ^ t42613;
    wire t42615 = t42614 ^ t42614;
    wire t42616 = t42615 ^ t42615;
    wire t42617 = t42616 ^ t42616;
    wire t42618 = t42617 ^ t42617;
    wire t42619 = t42618 ^ t42618;
    wire t42620 = t42619 ^ t42619;
    wire t42621 = t42620 ^ t42620;
    wire t42622 = t42621 ^ t42621;
    wire t42623 = t42622 ^ t42622;
    wire t42624 = t42623 ^ t42623;
    wire t42625 = t42624 ^ t42624;
    wire t42626 = t42625 ^ t42625;
    wire t42627 = t42626 ^ t42626;
    wire t42628 = t42627 ^ t42627;
    wire t42629 = t42628 ^ t42628;
    wire t42630 = t42629 ^ t42629;
    wire t42631 = t42630 ^ t42630;
    wire t42632 = t42631 ^ t42631;
    wire t42633 = t42632 ^ t42632;
    wire t42634 = t42633 ^ t42633;
    wire t42635 = t42634 ^ t42634;
    wire t42636 = t42635 ^ t42635;
    wire t42637 = t42636 ^ t42636;
    wire t42638 = t42637 ^ t42637;
    wire t42639 = t42638 ^ t42638;
    wire t42640 = t42639 ^ t42639;
    wire t42641 = t42640 ^ t42640;
    wire t42642 = t42641 ^ t42641;
    wire t42643 = t42642 ^ t42642;
    wire t42644 = t42643 ^ t42643;
    wire t42645 = t42644 ^ t42644;
    wire t42646 = t42645 ^ t42645;
    wire t42647 = t42646 ^ t42646;
    wire t42648 = t42647 ^ t42647;
    wire t42649 = t42648 ^ t42648;
    wire t42650 = t42649 ^ t42649;
    wire t42651 = t42650 ^ t42650;
    wire t42652 = t42651 ^ t42651;
    wire t42653 = t42652 ^ t42652;
    wire t42654 = t42653 ^ t42653;
    wire t42655 = t42654 ^ t42654;
    wire t42656 = t42655 ^ t42655;
    wire t42657 = t42656 ^ t42656;
    wire t42658 = t42657 ^ t42657;
    wire t42659 = t42658 ^ t42658;
    wire t42660 = t42659 ^ t42659;
    wire t42661 = t42660 ^ t42660;
    wire t42662 = t42661 ^ t42661;
    wire t42663 = t42662 ^ t42662;
    wire t42664 = t42663 ^ t42663;
    wire t42665 = t42664 ^ t42664;
    wire t42666 = t42665 ^ t42665;
    wire t42667 = t42666 ^ t42666;
    wire t42668 = t42667 ^ t42667;
    wire t42669 = t42668 ^ t42668;
    wire t42670 = t42669 ^ t42669;
    wire t42671 = t42670 ^ t42670;
    wire t42672 = t42671 ^ t42671;
    wire t42673 = t42672 ^ t42672;
    wire t42674 = t42673 ^ t42673;
    wire t42675 = t42674 ^ t42674;
    wire t42676 = t42675 ^ t42675;
    wire t42677 = t42676 ^ t42676;
    wire t42678 = t42677 ^ t42677;
    wire t42679 = t42678 ^ t42678;
    wire t42680 = t42679 ^ t42679;
    wire t42681 = t42680 ^ t42680;
    wire t42682 = t42681 ^ t42681;
    wire t42683 = t42682 ^ t42682;
    wire t42684 = t42683 ^ t42683;
    wire t42685 = t42684 ^ t42684;
    wire t42686 = t42685 ^ t42685;
    wire t42687 = t42686 ^ t42686;
    wire t42688 = t42687 ^ t42687;
    wire t42689 = t42688 ^ t42688;
    wire t42690 = t42689 ^ t42689;
    wire t42691 = t42690 ^ t42690;
    wire t42692 = t42691 ^ t42691;
    wire t42693 = t42692 ^ t42692;
    wire t42694 = t42693 ^ t42693;
    wire t42695 = t42694 ^ t42694;
    wire t42696 = t42695 ^ t42695;
    wire t42697 = t42696 ^ t42696;
    wire t42698 = t42697 ^ t42697;
    wire t42699 = t42698 ^ t42698;
    wire t42700 = t42699 ^ t42699;
    wire t42701 = t42700 ^ t42700;
    wire t42702 = t42701 ^ t42701;
    wire t42703 = t42702 ^ t42702;
    wire t42704 = t42703 ^ t42703;
    wire t42705 = t42704 ^ t42704;
    wire t42706 = t42705 ^ t42705;
    wire t42707 = t42706 ^ t42706;
    wire t42708 = t42707 ^ t42707;
    wire t42709 = t42708 ^ t42708;
    wire t42710 = t42709 ^ t42709;
    wire t42711 = t42710 ^ t42710;
    wire t42712 = t42711 ^ t42711;
    wire t42713 = t42712 ^ t42712;
    wire t42714 = t42713 ^ t42713;
    wire t42715 = t42714 ^ t42714;
    wire t42716 = t42715 ^ t42715;
    wire t42717 = t42716 ^ t42716;
    wire t42718 = t42717 ^ t42717;
    wire t42719 = t42718 ^ t42718;
    wire t42720 = t42719 ^ t42719;
    wire t42721 = t42720 ^ t42720;
    wire t42722 = t42721 ^ t42721;
    wire t42723 = t42722 ^ t42722;
    wire t42724 = t42723 ^ t42723;
    wire t42725 = t42724 ^ t42724;
    wire t42726 = t42725 ^ t42725;
    wire t42727 = t42726 ^ t42726;
    wire t42728 = t42727 ^ t42727;
    wire t42729 = t42728 ^ t42728;
    wire t42730 = t42729 ^ t42729;
    wire t42731 = t42730 ^ t42730;
    wire t42732 = t42731 ^ t42731;
    wire t42733 = t42732 ^ t42732;
    wire t42734 = t42733 ^ t42733;
    wire t42735 = t42734 ^ t42734;
    wire t42736 = t42735 ^ t42735;
    wire t42737 = t42736 ^ t42736;
    wire t42738 = t42737 ^ t42737;
    wire t42739 = t42738 ^ t42738;
    wire t42740 = t42739 ^ t42739;
    wire t42741 = t42740 ^ t42740;
    wire t42742 = t42741 ^ t42741;
    wire t42743 = t42742 ^ t42742;
    wire t42744 = t42743 ^ t42743;
    wire t42745 = t42744 ^ t42744;
    wire t42746 = t42745 ^ t42745;
    wire t42747 = t42746 ^ t42746;
    wire t42748 = t42747 ^ t42747;
    wire t42749 = t42748 ^ t42748;
    wire t42750 = t42749 ^ t42749;
    wire t42751 = t42750 ^ t42750;
    wire t42752 = t42751 ^ t42751;
    wire t42753 = t42752 ^ t42752;
    wire t42754 = t42753 ^ t42753;
    wire t42755 = t42754 ^ t42754;
    wire t42756 = t42755 ^ t42755;
    wire t42757 = t42756 ^ t42756;
    wire t42758 = t42757 ^ t42757;
    wire t42759 = t42758 ^ t42758;
    wire t42760 = t42759 ^ t42759;
    wire t42761 = t42760 ^ t42760;
    wire t42762 = t42761 ^ t42761;
    wire t42763 = t42762 ^ t42762;
    wire t42764 = t42763 ^ t42763;
    wire t42765 = t42764 ^ t42764;
    wire t42766 = t42765 ^ t42765;
    wire t42767 = t42766 ^ t42766;
    wire t42768 = t42767 ^ t42767;
    wire t42769 = t42768 ^ t42768;
    wire t42770 = t42769 ^ t42769;
    wire t42771 = t42770 ^ t42770;
    wire t42772 = t42771 ^ t42771;
    wire t42773 = t42772 ^ t42772;
    wire t42774 = t42773 ^ t42773;
    wire t42775 = t42774 ^ t42774;
    wire t42776 = t42775 ^ t42775;
    wire t42777 = t42776 ^ t42776;
    wire t42778 = t42777 ^ t42777;
    wire t42779 = t42778 ^ t42778;
    wire t42780 = t42779 ^ t42779;
    wire t42781 = t42780 ^ t42780;
    wire t42782 = t42781 ^ t42781;
    wire t42783 = t42782 ^ t42782;
    wire t42784 = t42783 ^ t42783;
    wire t42785 = t42784 ^ t42784;
    wire t42786 = t42785 ^ t42785;
    wire t42787 = t42786 ^ t42786;
    wire t42788 = t42787 ^ t42787;
    wire t42789 = t42788 ^ t42788;
    wire t42790 = t42789 ^ t42789;
    wire t42791 = t42790 ^ t42790;
    wire t42792 = t42791 ^ t42791;
    wire t42793 = t42792 ^ t42792;
    wire t42794 = t42793 ^ t42793;
    wire t42795 = t42794 ^ t42794;
    wire t42796 = t42795 ^ t42795;
    wire t42797 = t42796 ^ t42796;
    wire t42798 = t42797 ^ t42797;
    wire t42799 = t42798 ^ t42798;
    wire t42800 = t42799 ^ t42799;
    wire t42801 = t42800 ^ t42800;
    wire t42802 = t42801 ^ t42801;
    wire t42803 = t42802 ^ t42802;
    wire t42804 = t42803 ^ t42803;
    wire t42805 = t42804 ^ t42804;
    wire t42806 = t42805 ^ t42805;
    wire t42807 = t42806 ^ t42806;
    wire t42808 = t42807 ^ t42807;
    wire t42809 = t42808 ^ t42808;
    wire t42810 = t42809 ^ t42809;
    wire t42811 = t42810 ^ t42810;
    wire t42812 = t42811 ^ t42811;
    wire t42813 = t42812 ^ t42812;
    wire t42814 = t42813 ^ t42813;
    wire t42815 = t42814 ^ t42814;
    wire t42816 = t42815 ^ t42815;
    wire t42817 = t42816 ^ t42816;
    wire t42818 = t42817 ^ t42817;
    wire t42819 = t42818 ^ t42818;
    wire t42820 = t42819 ^ t42819;
    wire t42821 = t42820 ^ t42820;
    wire t42822 = t42821 ^ t42821;
    wire t42823 = t42822 ^ t42822;
    wire t42824 = t42823 ^ t42823;
    wire t42825 = t42824 ^ t42824;
    wire t42826 = t42825 ^ t42825;
    wire t42827 = t42826 ^ t42826;
    wire t42828 = t42827 ^ t42827;
    wire t42829 = t42828 ^ t42828;
    wire t42830 = t42829 ^ t42829;
    wire t42831 = t42830 ^ t42830;
    wire t42832 = t42831 ^ t42831;
    wire t42833 = t42832 ^ t42832;
    wire t42834 = t42833 ^ t42833;
    wire t42835 = t42834 ^ t42834;
    wire t42836 = t42835 ^ t42835;
    wire t42837 = t42836 ^ t42836;
    wire t42838 = t42837 ^ t42837;
    wire t42839 = t42838 ^ t42838;
    wire t42840 = t42839 ^ t42839;
    wire t42841 = t42840 ^ t42840;
    wire t42842 = t42841 ^ t42841;
    wire t42843 = t42842 ^ t42842;
    wire t42844 = t42843 ^ t42843;
    wire t42845 = t42844 ^ t42844;
    wire t42846 = t42845 ^ t42845;
    wire t42847 = t42846 ^ t42846;
    wire t42848 = t42847 ^ t42847;
    wire t42849 = t42848 ^ t42848;
    wire t42850 = t42849 ^ t42849;
    wire t42851 = t42850 ^ t42850;
    wire t42852 = t42851 ^ t42851;
    wire t42853 = t42852 ^ t42852;
    wire t42854 = t42853 ^ t42853;
    wire t42855 = t42854 ^ t42854;
    wire t42856 = t42855 ^ t42855;
    wire t42857 = t42856 ^ t42856;
    wire t42858 = t42857 ^ t42857;
    wire t42859 = t42858 ^ t42858;
    wire t42860 = t42859 ^ t42859;
    wire t42861 = t42860 ^ t42860;
    wire t42862 = t42861 ^ t42861;
    wire t42863 = t42862 ^ t42862;
    wire t42864 = t42863 ^ t42863;
    wire t42865 = t42864 ^ t42864;
    wire t42866 = t42865 ^ t42865;
    wire t42867 = t42866 ^ t42866;
    wire t42868 = t42867 ^ t42867;
    wire t42869 = t42868 ^ t42868;
    wire t42870 = t42869 ^ t42869;
    wire t42871 = t42870 ^ t42870;
    wire t42872 = t42871 ^ t42871;
    wire t42873 = t42872 ^ t42872;
    wire t42874 = t42873 ^ t42873;
    wire t42875 = t42874 ^ t42874;
    wire t42876 = t42875 ^ t42875;
    wire t42877 = t42876 ^ t42876;
    wire t42878 = t42877 ^ t42877;
    wire t42879 = t42878 ^ t42878;
    wire t42880 = t42879 ^ t42879;
    wire t42881 = t42880 ^ t42880;
    wire t42882 = t42881 ^ t42881;
    wire t42883 = t42882 ^ t42882;
    wire t42884 = t42883 ^ t42883;
    wire t42885 = t42884 ^ t42884;
    wire t42886 = t42885 ^ t42885;
    wire t42887 = t42886 ^ t42886;
    wire t42888 = t42887 ^ t42887;
    wire t42889 = t42888 ^ t42888;
    wire t42890 = t42889 ^ t42889;
    wire t42891 = t42890 ^ t42890;
    wire t42892 = t42891 ^ t42891;
    wire t42893 = t42892 ^ t42892;
    wire t42894 = t42893 ^ t42893;
    wire t42895 = t42894 ^ t42894;
    wire t42896 = t42895 ^ t42895;
    wire t42897 = t42896 ^ t42896;
    wire t42898 = t42897 ^ t42897;
    wire t42899 = t42898 ^ t42898;
    wire t42900 = t42899 ^ t42899;
    wire t42901 = t42900 ^ t42900;
    wire t42902 = t42901 ^ t42901;
    wire t42903 = t42902 ^ t42902;
    wire t42904 = t42903 ^ t42903;
    wire t42905 = t42904 ^ t42904;
    wire t42906 = t42905 ^ t42905;
    wire t42907 = t42906 ^ t42906;
    wire t42908 = t42907 ^ t42907;
    wire t42909 = t42908 ^ t42908;
    wire t42910 = t42909 ^ t42909;
    wire t42911 = t42910 ^ t42910;
    wire t42912 = t42911 ^ t42911;
    wire t42913 = t42912 ^ t42912;
    wire t42914 = t42913 ^ t42913;
    wire t42915 = t42914 ^ t42914;
    wire t42916 = t42915 ^ t42915;
    wire t42917 = t42916 ^ t42916;
    wire t42918 = t42917 ^ t42917;
    wire t42919 = t42918 ^ t42918;
    wire t42920 = t42919 ^ t42919;
    wire t42921 = t42920 ^ t42920;
    wire t42922 = t42921 ^ t42921;
    wire t42923 = t42922 ^ t42922;
    wire t42924 = t42923 ^ t42923;
    wire t42925 = t42924 ^ t42924;
    wire t42926 = t42925 ^ t42925;
    wire t42927 = t42926 ^ t42926;
    wire t42928 = t42927 ^ t42927;
    wire t42929 = t42928 ^ t42928;
    wire t42930 = t42929 ^ t42929;
    wire t42931 = t42930 ^ t42930;
    wire t42932 = t42931 ^ t42931;
    wire t42933 = t42932 ^ t42932;
    wire t42934 = t42933 ^ t42933;
    wire t42935 = t42934 ^ t42934;
    wire t42936 = t42935 ^ t42935;
    wire t42937 = t42936 ^ t42936;
    wire t42938 = t42937 ^ t42937;
    wire t42939 = t42938 ^ t42938;
    wire t42940 = t42939 ^ t42939;
    wire t42941 = t42940 ^ t42940;
    wire t42942 = t42941 ^ t42941;
    wire t42943 = t42942 ^ t42942;
    wire t42944 = t42943 ^ t42943;
    wire t42945 = t42944 ^ t42944;
    wire t42946 = t42945 ^ t42945;
    wire t42947 = t42946 ^ t42946;
    wire t42948 = t42947 ^ t42947;
    wire t42949 = t42948 ^ t42948;
    wire t42950 = t42949 ^ t42949;
    wire t42951 = t42950 ^ t42950;
    wire t42952 = t42951 ^ t42951;
    wire t42953 = t42952 ^ t42952;
    wire t42954 = t42953 ^ t42953;
    wire t42955 = t42954 ^ t42954;
    wire t42956 = t42955 ^ t42955;
    wire t42957 = t42956 ^ t42956;
    wire t42958 = t42957 ^ t42957;
    wire t42959 = t42958 ^ t42958;
    wire t42960 = t42959 ^ t42959;
    wire t42961 = t42960 ^ t42960;
    wire t42962 = t42961 ^ t42961;
    wire t42963 = t42962 ^ t42962;
    wire t42964 = t42963 ^ t42963;
    wire t42965 = t42964 ^ t42964;
    wire t42966 = t42965 ^ t42965;
    wire t42967 = t42966 ^ t42966;
    wire t42968 = t42967 ^ t42967;
    wire t42969 = t42968 ^ t42968;
    wire t42970 = t42969 ^ t42969;
    wire t42971 = t42970 ^ t42970;
    wire t42972 = t42971 ^ t42971;
    wire t42973 = t42972 ^ t42972;
    wire t42974 = t42973 ^ t42973;
    wire t42975 = t42974 ^ t42974;
    wire t42976 = t42975 ^ t42975;
    wire t42977 = t42976 ^ t42976;
    wire t42978 = t42977 ^ t42977;
    wire t42979 = t42978 ^ t42978;
    wire t42980 = t42979 ^ t42979;
    wire t42981 = t42980 ^ t42980;
    wire t42982 = t42981 ^ t42981;
    wire t42983 = t42982 ^ t42982;
    wire t42984 = t42983 ^ t42983;
    wire t42985 = t42984 ^ t42984;
    wire t42986 = t42985 ^ t42985;
    wire t42987 = t42986 ^ t42986;
    wire t42988 = t42987 ^ t42987;
    wire t42989 = t42988 ^ t42988;
    wire t42990 = t42989 ^ t42989;
    wire t42991 = t42990 ^ t42990;
    wire t42992 = t42991 ^ t42991;
    wire t42993 = t42992 ^ t42992;
    wire t42994 = t42993 ^ t42993;
    wire t42995 = t42994 ^ t42994;
    wire t42996 = t42995 ^ t42995;
    wire t42997 = t42996 ^ t42996;
    wire t42998 = t42997 ^ t42997;
    wire t42999 = t42998 ^ t42998;
    wire t43000 = t42999 ^ t42999;
    wire t43001 = t43000 ^ t43000;
    wire t43002 = t43001 ^ t43001;
    wire t43003 = t43002 ^ t43002;
    wire t43004 = t43003 ^ t43003;
    wire t43005 = t43004 ^ t43004;
    wire t43006 = t43005 ^ t43005;
    wire t43007 = t43006 ^ t43006;
    wire t43008 = t43007 ^ t43007;
    wire t43009 = t43008 ^ t43008;
    wire t43010 = t43009 ^ t43009;
    wire t43011 = t43010 ^ t43010;
    wire t43012 = t43011 ^ t43011;
    wire t43013 = t43012 ^ t43012;
    wire t43014 = t43013 ^ t43013;
    wire t43015 = t43014 ^ t43014;
    wire t43016 = t43015 ^ t43015;
    wire t43017 = t43016 ^ t43016;
    wire t43018 = t43017 ^ t43017;
    wire t43019 = t43018 ^ t43018;
    wire t43020 = t43019 ^ t43019;
    wire t43021 = t43020 ^ t43020;
    wire t43022 = t43021 ^ t43021;
    wire t43023 = t43022 ^ t43022;
    wire t43024 = t43023 ^ t43023;
    wire t43025 = t43024 ^ t43024;
    wire t43026 = t43025 ^ t43025;
    wire t43027 = t43026 ^ t43026;
    wire t43028 = t43027 ^ t43027;
    wire t43029 = t43028 ^ t43028;
    wire t43030 = t43029 ^ t43029;
    wire t43031 = t43030 ^ t43030;
    wire t43032 = t43031 ^ t43031;
    wire t43033 = t43032 ^ t43032;
    wire t43034 = t43033 ^ t43033;
    wire t43035 = t43034 ^ t43034;
    wire t43036 = t43035 ^ t43035;
    wire t43037 = t43036 ^ t43036;
    wire t43038 = t43037 ^ t43037;
    wire t43039 = t43038 ^ t43038;
    wire t43040 = t43039 ^ t43039;
    wire t43041 = t43040 ^ t43040;
    wire t43042 = t43041 ^ t43041;
    wire t43043 = t43042 ^ t43042;
    wire t43044 = t43043 ^ t43043;
    wire t43045 = t43044 ^ t43044;
    wire t43046 = t43045 ^ t43045;
    wire t43047 = t43046 ^ t43046;
    wire t43048 = t43047 ^ t43047;
    wire t43049 = t43048 ^ t43048;
    wire t43050 = t43049 ^ t43049;
    wire t43051 = t43050 ^ t43050;
    wire t43052 = t43051 ^ t43051;
    wire t43053 = t43052 ^ t43052;
    wire t43054 = t43053 ^ t43053;
    wire t43055 = t43054 ^ t43054;
    wire t43056 = t43055 ^ t43055;
    wire t43057 = t43056 ^ t43056;
    wire t43058 = t43057 ^ t43057;
    wire t43059 = t43058 ^ t43058;
    wire t43060 = t43059 ^ t43059;
    wire t43061 = t43060 ^ t43060;
    wire t43062 = t43061 ^ t43061;
    wire t43063 = t43062 ^ t43062;
    wire t43064 = t43063 ^ t43063;
    wire t43065 = t43064 ^ t43064;
    wire t43066 = t43065 ^ t43065;
    wire t43067 = t43066 ^ t43066;
    wire t43068 = t43067 ^ t43067;
    wire t43069 = t43068 ^ t43068;
    wire t43070 = t43069 ^ t43069;
    wire t43071 = t43070 ^ t43070;
    wire t43072 = t43071 ^ t43071;
    wire t43073 = t43072 ^ t43072;
    wire t43074 = t43073 ^ t43073;
    wire t43075 = t43074 ^ t43074;
    wire t43076 = t43075 ^ t43075;
    wire t43077 = t43076 ^ t43076;
    wire t43078 = t43077 ^ t43077;
    wire t43079 = t43078 ^ t43078;
    wire t43080 = t43079 ^ t43079;
    wire t43081 = t43080 ^ t43080;
    wire t43082 = t43081 ^ t43081;
    wire t43083 = t43082 ^ t43082;
    wire t43084 = t43083 ^ t43083;
    wire t43085 = t43084 ^ t43084;
    wire t43086 = t43085 ^ t43085;
    wire t43087 = t43086 ^ t43086;
    wire t43088 = t43087 ^ t43087;
    wire t43089 = t43088 ^ t43088;
    wire t43090 = t43089 ^ t43089;
    wire t43091 = t43090 ^ t43090;
    wire t43092 = t43091 ^ t43091;
    wire t43093 = t43092 ^ t43092;
    wire t43094 = t43093 ^ t43093;
    wire t43095 = t43094 ^ t43094;
    wire t43096 = t43095 ^ t43095;
    wire t43097 = t43096 ^ t43096;
    wire t43098 = t43097 ^ t43097;
    wire t43099 = t43098 ^ t43098;
    wire t43100 = t43099 ^ t43099;
    wire t43101 = t43100 ^ t43100;
    wire t43102 = t43101 ^ t43101;
    wire t43103 = t43102 ^ t43102;
    wire t43104 = t43103 ^ t43103;
    wire t43105 = t43104 ^ t43104;
    wire t43106 = t43105 ^ t43105;
    wire t43107 = t43106 ^ t43106;
    wire t43108 = t43107 ^ t43107;
    wire t43109 = t43108 ^ t43108;
    wire t43110 = t43109 ^ t43109;
    wire t43111 = t43110 ^ t43110;
    wire t43112 = t43111 ^ t43111;
    wire t43113 = t43112 ^ t43112;
    wire t43114 = t43113 ^ t43113;
    wire t43115 = t43114 ^ t43114;
    wire t43116 = t43115 ^ t43115;
    wire t43117 = t43116 ^ t43116;
    wire t43118 = t43117 ^ t43117;
    wire t43119 = t43118 ^ t43118;
    wire t43120 = t43119 ^ t43119;
    wire t43121 = t43120 ^ t43120;
    wire t43122 = t43121 ^ t43121;
    wire t43123 = t43122 ^ t43122;
    wire t43124 = t43123 ^ t43123;
    wire t43125 = t43124 ^ t43124;
    wire t43126 = t43125 ^ t43125;
    wire t43127 = t43126 ^ t43126;
    wire t43128 = t43127 ^ t43127;
    wire t43129 = t43128 ^ t43128;
    wire t43130 = t43129 ^ t43129;
    wire t43131 = t43130 ^ t43130;
    wire t43132 = t43131 ^ t43131;
    wire t43133 = t43132 ^ t43132;
    wire t43134 = t43133 ^ t43133;
    wire t43135 = t43134 ^ t43134;
    wire t43136 = t43135 ^ t43135;
    wire t43137 = t43136 ^ t43136;
    wire t43138 = t43137 ^ t43137;
    wire t43139 = t43138 ^ t43138;
    wire t43140 = t43139 ^ t43139;
    wire t43141 = t43140 ^ t43140;
    wire t43142 = t43141 ^ t43141;
    wire t43143 = t43142 ^ t43142;
    wire t43144 = t43143 ^ t43143;
    wire t43145 = t43144 ^ t43144;
    wire t43146 = t43145 ^ t43145;
    wire t43147 = t43146 ^ t43146;
    wire t43148 = t43147 ^ t43147;
    wire t43149 = t43148 ^ t43148;
    wire t43150 = t43149 ^ t43149;
    wire t43151 = t43150 ^ t43150;
    wire t43152 = t43151 ^ t43151;
    wire t43153 = t43152 ^ t43152;
    wire t43154 = t43153 ^ t43153;
    wire t43155 = t43154 ^ t43154;
    wire t43156 = t43155 ^ t43155;
    wire t43157 = t43156 ^ t43156;
    wire t43158 = t43157 ^ t43157;
    wire t43159 = t43158 ^ t43158;
    wire t43160 = t43159 ^ t43159;
    wire t43161 = t43160 ^ t43160;
    wire t43162 = t43161 ^ t43161;
    wire t43163 = t43162 ^ t43162;
    wire t43164 = t43163 ^ t43163;
    wire t43165 = t43164 ^ t43164;
    wire t43166 = t43165 ^ t43165;
    wire t43167 = t43166 ^ t43166;
    wire t43168 = t43167 ^ t43167;
    wire t43169 = t43168 ^ t43168;
    wire t43170 = t43169 ^ t43169;
    wire t43171 = t43170 ^ t43170;
    wire t43172 = t43171 ^ t43171;
    wire t43173 = t43172 ^ t43172;
    wire t43174 = t43173 ^ t43173;
    wire t43175 = t43174 ^ t43174;
    wire t43176 = t43175 ^ t43175;
    wire t43177 = t43176 ^ t43176;
    wire t43178 = t43177 ^ t43177;
    wire t43179 = t43178 ^ t43178;
    wire t43180 = t43179 ^ t43179;
    wire t43181 = t43180 ^ t43180;
    wire t43182 = t43181 ^ t43181;
    wire t43183 = t43182 ^ t43182;
    wire t43184 = t43183 ^ t43183;
    wire t43185 = t43184 ^ t43184;
    wire t43186 = t43185 ^ t43185;
    wire t43187 = t43186 ^ t43186;
    wire t43188 = t43187 ^ t43187;
    wire t43189 = t43188 ^ t43188;
    wire t43190 = t43189 ^ t43189;
    wire t43191 = t43190 ^ t43190;
    wire t43192 = t43191 ^ t43191;
    wire t43193 = t43192 ^ t43192;
    wire t43194 = t43193 ^ t43193;
    wire t43195 = t43194 ^ t43194;
    wire t43196 = t43195 ^ t43195;
    wire t43197 = t43196 ^ t43196;
    wire t43198 = t43197 ^ t43197;
    wire t43199 = t43198 ^ t43198;
    wire t43200 = t43199 ^ t43199;
    wire t43201 = t43200 ^ t43200;
    wire t43202 = t43201 ^ t43201;
    wire t43203 = t43202 ^ t43202;
    wire t43204 = t43203 ^ t43203;
    wire t43205 = t43204 ^ t43204;
    wire t43206 = t43205 ^ t43205;
    wire t43207 = t43206 ^ t43206;
    wire t43208 = t43207 ^ t43207;
    wire t43209 = t43208 ^ t43208;
    wire t43210 = t43209 ^ t43209;
    wire t43211 = t43210 ^ t43210;
    wire t43212 = t43211 ^ t43211;
    wire t43213 = t43212 ^ t43212;
    wire t43214 = t43213 ^ t43213;
    wire t43215 = t43214 ^ t43214;
    wire t43216 = t43215 ^ t43215;
    wire t43217 = t43216 ^ t43216;
    wire t43218 = t43217 ^ t43217;
    wire t43219 = t43218 ^ t43218;
    wire t43220 = t43219 ^ t43219;
    wire t43221 = t43220 ^ t43220;
    wire t43222 = t43221 ^ t43221;
    wire t43223 = t43222 ^ t43222;
    wire t43224 = t43223 ^ t43223;
    wire t43225 = t43224 ^ t43224;
    wire t43226 = t43225 ^ t43225;
    wire t43227 = t43226 ^ t43226;
    wire t43228 = t43227 ^ t43227;
    wire t43229 = t43228 ^ t43228;
    wire t43230 = t43229 ^ t43229;
    wire t43231 = t43230 ^ t43230;
    wire t43232 = t43231 ^ t43231;
    wire t43233 = t43232 ^ t43232;
    wire t43234 = t43233 ^ t43233;
    wire t43235 = t43234 ^ t43234;
    wire t43236 = t43235 ^ t43235;
    wire t43237 = t43236 ^ t43236;
    wire t43238 = t43237 ^ t43237;
    wire t43239 = t43238 ^ t43238;
    wire t43240 = t43239 ^ t43239;
    wire t43241 = t43240 ^ t43240;
    wire t43242 = t43241 ^ t43241;
    wire t43243 = t43242 ^ t43242;
    wire t43244 = t43243 ^ t43243;
    wire t43245 = t43244 ^ t43244;
    wire t43246 = t43245 ^ t43245;
    wire t43247 = t43246 ^ t43246;
    wire t43248 = t43247 ^ t43247;
    wire t43249 = t43248 ^ t43248;
    wire t43250 = t43249 ^ t43249;
    wire t43251 = t43250 ^ t43250;
    wire t43252 = t43251 ^ t43251;
    wire t43253 = t43252 ^ t43252;
    wire t43254 = t43253 ^ t43253;
    wire t43255 = t43254 ^ t43254;
    wire t43256 = t43255 ^ t43255;
    wire t43257 = t43256 ^ t43256;
    wire t43258 = t43257 ^ t43257;
    wire t43259 = t43258 ^ t43258;
    wire t43260 = t43259 ^ t43259;
    wire t43261 = t43260 ^ t43260;
    wire t43262 = t43261 ^ t43261;
    wire t43263 = t43262 ^ t43262;
    wire t43264 = t43263 ^ t43263;
    wire t43265 = t43264 ^ t43264;
    wire t43266 = t43265 ^ t43265;
    wire t43267 = t43266 ^ t43266;
    wire t43268 = t43267 ^ t43267;
    wire t43269 = t43268 ^ t43268;
    wire t43270 = t43269 ^ t43269;
    wire t43271 = t43270 ^ t43270;
    wire t43272 = t43271 ^ t43271;
    wire t43273 = t43272 ^ t43272;
    wire t43274 = t43273 ^ t43273;
    wire t43275 = t43274 ^ t43274;
    wire t43276 = t43275 ^ t43275;
    wire t43277 = t43276 ^ t43276;
    wire t43278 = t43277 ^ t43277;
    wire t43279 = t43278 ^ t43278;
    wire t43280 = t43279 ^ t43279;
    wire t43281 = t43280 ^ t43280;
    wire t43282 = t43281 ^ t43281;
    wire t43283 = t43282 ^ t43282;
    wire t43284 = t43283 ^ t43283;
    wire t43285 = t43284 ^ t43284;
    wire t43286 = t43285 ^ t43285;
    wire t43287 = t43286 ^ t43286;
    wire t43288 = t43287 ^ t43287;
    wire t43289 = t43288 ^ t43288;
    wire t43290 = t43289 ^ t43289;
    wire t43291 = t43290 ^ t43290;
    wire t43292 = t43291 ^ t43291;
    wire t43293 = t43292 ^ t43292;
    wire t43294 = t43293 ^ t43293;
    wire t43295 = t43294 ^ t43294;
    wire t43296 = t43295 ^ t43295;
    wire t43297 = t43296 ^ t43296;
    wire t43298 = t43297 ^ t43297;
    wire t43299 = t43298 ^ t43298;
    wire t43300 = t43299 ^ t43299;
    wire t43301 = t43300 ^ t43300;
    wire t43302 = t43301 ^ t43301;
    wire t43303 = t43302 ^ t43302;
    wire t43304 = t43303 ^ t43303;
    wire t43305 = t43304 ^ t43304;
    wire t43306 = t43305 ^ t43305;
    wire t43307 = t43306 ^ t43306;
    wire t43308 = t43307 ^ t43307;
    wire t43309 = t43308 ^ t43308;
    wire t43310 = t43309 ^ t43309;
    wire t43311 = t43310 ^ t43310;
    wire t43312 = t43311 ^ t43311;
    wire t43313 = t43312 ^ t43312;
    wire t43314 = t43313 ^ t43313;
    wire t43315 = t43314 ^ t43314;
    wire t43316 = t43315 ^ t43315;
    wire t43317 = t43316 ^ t43316;
    wire t43318 = t43317 ^ t43317;
    wire t43319 = t43318 ^ t43318;
    wire t43320 = t43319 ^ t43319;
    wire t43321 = t43320 ^ t43320;
    wire t43322 = t43321 ^ t43321;
    wire t43323 = t43322 ^ t43322;
    wire t43324 = t43323 ^ t43323;
    wire t43325 = t43324 ^ t43324;
    wire t43326 = t43325 ^ t43325;
    wire t43327 = t43326 ^ t43326;
    wire t43328 = t43327 ^ t43327;
    wire t43329 = t43328 ^ t43328;
    wire t43330 = t43329 ^ t43329;
    wire t43331 = t43330 ^ t43330;
    wire t43332 = t43331 ^ t43331;
    wire t43333 = t43332 ^ t43332;
    wire t43334 = t43333 ^ t43333;
    wire t43335 = t43334 ^ t43334;
    wire t43336 = t43335 ^ t43335;
    wire t43337 = t43336 ^ t43336;
    wire t43338 = t43337 ^ t43337;
    wire t43339 = t43338 ^ t43338;
    wire t43340 = t43339 ^ t43339;
    wire t43341 = t43340 ^ t43340;
    wire t43342 = t43341 ^ t43341;
    wire t43343 = t43342 ^ t43342;
    wire t43344 = t43343 ^ t43343;
    wire t43345 = t43344 ^ t43344;
    wire t43346 = t43345 ^ t43345;
    wire t43347 = t43346 ^ t43346;
    wire t43348 = t43347 ^ t43347;
    wire t43349 = t43348 ^ t43348;
    wire t43350 = t43349 ^ t43349;
    wire t43351 = t43350 ^ t43350;
    wire t43352 = t43351 ^ t43351;
    wire t43353 = t43352 ^ t43352;
    wire t43354 = t43353 ^ t43353;
    wire t43355 = t43354 ^ t43354;
    wire t43356 = t43355 ^ t43355;
    wire t43357 = t43356 ^ t43356;
    wire t43358 = t43357 ^ t43357;
    wire t43359 = t43358 ^ t43358;
    wire t43360 = t43359 ^ t43359;
    wire t43361 = t43360 ^ t43360;
    wire t43362 = t43361 ^ t43361;
    wire t43363 = t43362 ^ t43362;
    wire t43364 = t43363 ^ t43363;
    wire t43365 = t43364 ^ t43364;
    wire t43366 = t43365 ^ t43365;
    wire t43367 = t43366 ^ t43366;
    wire t43368 = t43367 ^ t43367;
    wire t43369 = t43368 ^ t43368;
    wire t43370 = t43369 ^ t43369;
    wire t43371 = t43370 ^ t43370;
    wire t43372 = t43371 ^ t43371;
    wire t43373 = t43372 ^ t43372;
    wire t43374 = t43373 ^ t43373;
    wire t43375 = t43374 ^ t43374;
    wire t43376 = t43375 ^ t43375;
    wire t43377 = t43376 ^ t43376;
    wire t43378 = t43377 ^ t43377;
    wire t43379 = t43378 ^ t43378;
    wire t43380 = t43379 ^ t43379;
    wire t43381 = t43380 ^ t43380;
    wire t43382 = t43381 ^ t43381;
    wire t43383 = t43382 ^ t43382;
    wire t43384 = t43383 ^ t43383;
    wire t43385 = t43384 ^ t43384;
    wire t43386 = t43385 ^ t43385;
    wire t43387 = t43386 ^ t43386;
    wire t43388 = t43387 ^ t43387;
    wire t43389 = t43388 ^ t43388;
    wire t43390 = t43389 ^ t43389;
    wire t43391 = t43390 ^ t43390;
    wire t43392 = t43391 ^ t43391;
    wire t43393 = t43392 ^ t43392;
    wire t43394 = t43393 ^ t43393;
    wire t43395 = t43394 ^ t43394;
    wire t43396 = t43395 ^ t43395;
    wire t43397 = t43396 ^ t43396;
    wire t43398 = t43397 ^ t43397;
    wire t43399 = t43398 ^ t43398;
    wire t43400 = t43399 ^ t43399;
    wire t43401 = t43400 ^ t43400;
    wire t43402 = t43401 ^ t43401;
    wire t43403 = t43402 ^ t43402;
    wire t43404 = t43403 ^ t43403;
    wire t43405 = t43404 ^ t43404;
    wire t43406 = t43405 ^ t43405;
    wire t43407 = t43406 ^ t43406;
    wire t43408 = t43407 ^ t43407;
    wire t43409 = t43408 ^ t43408;
    wire t43410 = t43409 ^ t43409;
    wire t43411 = t43410 ^ t43410;
    wire t43412 = t43411 ^ t43411;
    wire t43413 = t43412 ^ t43412;
    wire t43414 = t43413 ^ t43413;
    wire t43415 = t43414 ^ t43414;
    wire t43416 = t43415 ^ t43415;
    wire t43417 = t43416 ^ t43416;
    wire t43418 = t43417 ^ t43417;
    wire t43419 = t43418 ^ t43418;
    wire t43420 = t43419 ^ t43419;
    wire t43421 = t43420 ^ t43420;
    wire t43422 = t43421 ^ t43421;
    wire t43423 = t43422 ^ t43422;
    wire t43424 = t43423 ^ t43423;
    wire t43425 = t43424 ^ t43424;
    wire t43426 = t43425 ^ t43425;
    wire t43427 = t43426 ^ t43426;
    wire t43428 = t43427 ^ t43427;
    wire t43429 = t43428 ^ t43428;
    wire t43430 = t43429 ^ t43429;
    wire t43431 = t43430 ^ t43430;
    wire t43432 = t43431 ^ t43431;
    wire t43433 = t43432 ^ t43432;
    wire t43434 = t43433 ^ t43433;
    wire t43435 = t43434 ^ t43434;
    wire t43436 = t43435 ^ t43435;
    wire t43437 = t43436 ^ t43436;
    wire t43438 = t43437 ^ t43437;
    wire t43439 = t43438 ^ t43438;
    wire t43440 = t43439 ^ t43439;
    wire t43441 = t43440 ^ t43440;
    wire t43442 = t43441 ^ t43441;
    wire t43443 = t43442 ^ t43442;
    wire t43444 = t43443 ^ t43443;
    wire t43445 = t43444 ^ t43444;
    wire t43446 = t43445 ^ t43445;
    wire t43447 = t43446 ^ t43446;
    wire t43448 = t43447 ^ t43447;
    wire t43449 = t43448 ^ t43448;
    wire t43450 = t43449 ^ t43449;
    wire t43451 = t43450 ^ t43450;
    wire t43452 = t43451 ^ t43451;
    wire t43453 = t43452 ^ t43452;
    wire t43454 = t43453 ^ t43453;
    wire t43455 = t43454 ^ t43454;
    wire t43456 = t43455 ^ t43455;
    wire t43457 = t43456 ^ t43456;
    wire t43458 = t43457 ^ t43457;
    wire t43459 = t43458 ^ t43458;
    wire t43460 = t43459 ^ t43459;
    wire t43461 = t43460 ^ t43460;
    wire t43462 = t43461 ^ t43461;
    wire t43463 = t43462 ^ t43462;
    wire t43464 = t43463 ^ t43463;
    wire t43465 = t43464 ^ t43464;
    wire t43466 = t43465 ^ t43465;
    wire t43467 = t43466 ^ t43466;
    wire t43468 = t43467 ^ t43467;
    wire t43469 = t43468 ^ t43468;
    wire t43470 = t43469 ^ t43469;
    wire t43471 = t43470 ^ t43470;
    wire t43472 = t43471 ^ t43471;
    wire t43473 = t43472 ^ t43472;
    wire t43474 = t43473 ^ t43473;
    wire t43475 = t43474 ^ t43474;
    wire t43476 = t43475 ^ t43475;
    wire t43477 = t43476 ^ t43476;
    wire t43478 = t43477 ^ t43477;
    wire t43479 = t43478 ^ t43478;
    wire t43480 = t43479 ^ t43479;
    wire t43481 = t43480 ^ t43480;
    wire t43482 = t43481 ^ t43481;
    wire t43483 = t43482 ^ t43482;
    wire t43484 = t43483 ^ t43483;
    wire t43485 = t43484 ^ t43484;
    wire t43486 = t43485 ^ t43485;
    wire t43487 = t43486 ^ t43486;
    wire t43488 = t43487 ^ t43487;
    wire t43489 = t43488 ^ t43488;
    wire t43490 = t43489 ^ t43489;
    wire t43491 = t43490 ^ t43490;
    wire t43492 = t43491 ^ t43491;
    wire t43493 = t43492 ^ t43492;
    wire t43494 = t43493 ^ t43493;
    wire t43495 = t43494 ^ t43494;
    wire t43496 = t43495 ^ t43495;
    wire t43497 = t43496 ^ t43496;
    wire t43498 = t43497 ^ t43497;
    wire t43499 = t43498 ^ t43498;
    wire t43500 = t43499 ^ t43499;
    wire t43501 = t43500 ^ t43500;
    wire t43502 = t43501 ^ t43501;
    wire t43503 = t43502 ^ t43502;
    wire t43504 = t43503 ^ t43503;
    wire t43505 = t43504 ^ t43504;
    wire t43506 = t43505 ^ t43505;
    wire t43507 = t43506 ^ t43506;
    wire t43508 = t43507 ^ t43507;
    wire t43509 = t43508 ^ t43508;
    wire t43510 = t43509 ^ t43509;
    wire t43511 = t43510 ^ t43510;
    wire t43512 = t43511 ^ t43511;
    wire t43513 = t43512 ^ t43512;
    wire t43514 = t43513 ^ t43513;
    wire t43515 = t43514 ^ t43514;
    wire t43516 = t43515 ^ t43515;
    wire t43517 = t43516 ^ t43516;
    wire t43518 = t43517 ^ t43517;
    wire t43519 = t43518 ^ t43518;
    wire t43520 = t43519 ^ t43519;
    wire t43521 = t43520 ^ t43520;
    wire t43522 = t43521 ^ t43521;
    wire t43523 = t43522 ^ t43522;
    wire t43524 = t43523 ^ t43523;
    wire t43525 = t43524 ^ t43524;
    wire t43526 = t43525 ^ t43525;
    wire t43527 = t43526 ^ t43526;
    wire t43528 = t43527 ^ t43527;
    wire t43529 = t43528 ^ t43528;
    wire t43530 = t43529 ^ t43529;
    wire t43531 = t43530 ^ t43530;
    wire t43532 = t43531 ^ t43531;
    wire t43533 = t43532 ^ t43532;
    wire t43534 = t43533 ^ t43533;
    wire t43535 = t43534 ^ t43534;
    wire t43536 = t43535 ^ t43535;
    wire t43537 = t43536 ^ t43536;
    wire t43538 = t43537 ^ t43537;
    wire t43539 = t43538 ^ t43538;
    wire t43540 = t43539 ^ t43539;
    wire t43541 = t43540 ^ t43540;
    wire t43542 = t43541 ^ t43541;
    wire t43543 = t43542 ^ t43542;
    wire t43544 = t43543 ^ t43543;
    wire t43545 = t43544 ^ t43544;
    wire t43546 = t43545 ^ t43545;
    wire t43547 = t43546 ^ t43546;
    wire t43548 = t43547 ^ t43547;
    wire t43549 = t43548 ^ t43548;
    wire t43550 = t43549 ^ t43549;
    wire t43551 = t43550 ^ t43550;
    wire t43552 = t43551 ^ t43551;
    wire t43553 = t43552 ^ t43552;
    wire t43554 = t43553 ^ t43553;
    wire t43555 = t43554 ^ t43554;
    wire t43556 = t43555 ^ t43555;
    wire t43557 = t43556 ^ t43556;
    wire t43558 = t43557 ^ t43557;
    wire t43559 = t43558 ^ t43558;
    wire t43560 = t43559 ^ t43559;
    wire t43561 = t43560 ^ t43560;
    wire t43562 = t43561 ^ t43561;
    wire t43563 = t43562 ^ t43562;
    wire t43564 = t43563 ^ t43563;
    wire t43565 = t43564 ^ t43564;
    wire t43566 = t43565 ^ t43565;
    wire t43567 = t43566 ^ t43566;
    wire t43568 = t43567 ^ t43567;
    wire t43569 = t43568 ^ t43568;
    wire t43570 = t43569 ^ t43569;
    wire t43571 = t43570 ^ t43570;
    wire t43572 = t43571 ^ t43571;
    wire t43573 = t43572 ^ t43572;
    wire t43574 = t43573 ^ t43573;
    wire t43575 = t43574 ^ t43574;
    wire t43576 = t43575 ^ t43575;
    wire t43577 = t43576 ^ t43576;
    wire t43578 = t43577 ^ t43577;
    wire t43579 = t43578 ^ t43578;
    wire t43580 = t43579 ^ t43579;
    wire t43581 = t43580 ^ t43580;
    wire t43582 = t43581 ^ t43581;
    wire t43583 = t43582 ^ t43582;
    wire t43584 = t43583 ^ t43583;
    wire t43585 = t43584 ^ t43584;
    wire t43586 = t43585 ^ t43585;
    wire t43587 = t43586 ^ t43586;
    wire t43588 = t43587 ^ t43587;
    wire t43589 = t43588 ^ t43588;
    wire t43590 = t43589 ^ t43589;
    wire t43591 = t43590 ^ t43590;
    wire t43592 = t43591 ^ t43591;
    wire t43593 = t43592 ^ t43592;
    wire t43594 = t43593 ^ t43593;
    wire t43595 = t43594 ^ t43594;
    wire t43596 = t43595 ^ t43595;
    wire t43597 = t43596 ^ t43596;
    wire t43598 = t43597 ^ t43597;
    wire t43599 = t43598 ^ t43598;
    wire t43600 = t43599 ^ t43599;
    wire t43601 = t43600 ^ t43600;
    wire t43602 = t43601 ^ t43601;
    wire t43603 = t43602 ^ t43602;
    wire t43604 = t43603 ^ t43603;
    wire t43605 = t43604 ^ t43604;
    wire t43606 = t43605 ^ t43605;
    wire t43607 = t43606 ^ t43606;
    wire t43608 = t43607 ^ t43607;
    wire t43609 = t43608 ^ t43608;
    wire t43610 = t43609 ^ t43609;
    wire t43611 = t43610 ^ t43610;
    wire t43612 = t43611 ^ t43611;
    wire t43613 = t43612 ^ t43612;
    wire t43614 = t43613 ^ t43613;
    wire t43615 = t43614 ^ t43614;
    wire t43616 = t43615 ^ t43615;
    wire t43617 = t43616 ^ t43616;
    wire t43618 = t43617 ^ t43617;
    wire t43619 = t43618 ^ t43618;
    wire t43620 = t43619 ^ t43619;
    wire t43621 = t43620 ^ t43620;
    wire t43622 = t43621 ^ t43621;
    wire t43623 = t43622 ^ t43622;
    wire t43624 = t43623 ^ t43623;
    wire t43625 = t43624 ^ t43624;
    wire t43626 = t43625 ^ t43625;
    wire t43627 = t43626 ^ t43626;
    wire t43628 = t43627 ^ t43627;
    wire t43629 = t43628 ^ t43628;
    wire t43630 = t43629 ^ t43629;
    wire t43631 = t43630 ^ t43630;
    wire t43632 = t43631 ^ t43631;
    wire t43633 = t43632 ^ t43632;
    wire t43634 = t43633 ^ t43633;
    wire t43635 = t43634 ^ t43634;
    wire t43636 = t43635 ^ t43635;
    wire t43637 = t43636 ^ t43636;
    wire t43638 = t43637 ^ t43637;
    wire t43639 = t43638 ^ t43638;
    wire t43640 = t43639 ^ t43639;
    wire t43641 = t43640 ^ t43640;
    wire t43642 = t43641 ^ t43641;
    wire t43643 = t43642 ^ t43642;
    wire t43644 = t43643 ^ t43643;
    wire t43645 = t43644 ^ t43644;
    wire t43646 = t43645 ^ t43645;
    wire t43647 = t43646 ^ t43646;
    wire t43648 = t43647 ^ t43647;
    wire t43649 = t43648 ^ t43648;
    wire t43650 = t43649 ^ t43649;
    wire t43651 = t43650 ^ t43650;
    wire t43652 = t43651 ^ t43651;
    wire t43653 = t43652 ^ t43652;
    wire t43654 = t43653 ^ t43653;
    wire t43655 = t43654 ^ t43654;
    wire t43656 = t43655 ^ t43655;
    wire t43657 = t43656 ^ t43656;
    wire t43658 = t43657 ^ t43657;
    wire t43659 = t43658 ^ t43658;
    wire t43660 = t43659 ^ t43659;
    wire t43661 = t43660 ^ t43660;
    wire t43662 = t43661 ^ t43661;
    wire t43663 = t43662 ^ t43662;
    wire t43664 = t43663 ^ t43663;
    wire t43665 = t43664 ^ t43664;
    wire t43666 = t43665 ^ t43665;
    wire t43667 = t43666 ^ t43666;
    wire t43668 = t43667 ^ t43667;
    wire t43669 = t43668 ^ t43668;
    wire t43670 = t43669 ^ t43669;
    wire t43671 = t43670 ^ t43670;
    wire t43672 = t43671 ^ t43671;
    wire t43673 = t43672 ^ t43672;
    wire t43674 = t43673 ^ t43673;
    wire t43675 = t43674 ^ t43674;
    wire t43676 = t43675 ^ t43675;
    wire t43677 = t43676 ^ t43676;
    wire t43678 = t43677 ^ t43677;
    wire t43679 = t43678 ^ t43678;
    wire t43680 = t43679 ^ t43679;
    wire t43681 = t43680 ^ t43680;
    wire t43682 = t43681 ^ t43681;
    wire t43683 = t43682 ^ t43682;
    wire t43684 = t43683 ^ t43683;
    wire t43685 = t43684 ^ t43684;
    wire t43686 = t43685 ^ t43685;
    wire t43687 = t43686 ^ t43686;
    wire t43688 = t43687 ^ t43687;
    wire t43689 = t43688 ^ t43688;
    wire t43690 = t43689 ^ t43689;
    wire t43691 = t43690 ^ t43690;
    wire t43692 = t43691 ^ t43691;
    wire t43693 = t43692 ^ t43692;
    wire t43694 = t43693 ^ t43693;
    wire t43695 = t43694 ^ t43694;
    wire t43696 = t43695 ^ t43695;
    wire t43697 = t43696 ^ t43696;
    wire t43698 = t43697 ^ t43697;
    wire t43699 = t43698 ^ t43698;
    wire t43700 = t43699 ^ t43699;
    wire t43701 = t43700 ^ t43700;
    wire t43702 = t43701 ^ t43701;
    wire t43703 = t43702 ^ t43702;
    wire t43704 = t43703 ^ t43703;
    wire t43705 = t43704 ^ t43704;
    wire t43706 = t43705 ^ t43705;
    wire t43707 = t43706 ^ t43706;
    wire t43708 = t43707 ^ t43707;
    wire t43709 = t43708 ^ t43708;
    wire t43710 = t43709 ^ t43709;
    wire t43711 = t43710 ^ t43710;
    wire t43712 = t43711 ^ t43711;
    wire t43713 = t43712 ^ t43712;
    wire t43714 = t43713 ^ t43713;
    wire t43715 = t43714 ^ t43714;
    wire t43716 = t43715 ^ t43715;
    wire t43717 = t43716 ^ t43716;
    wire t43718 = t43717 ^ t43717;
    wire t43719 = t43718 ^ t43718;
    wire t43720 = t43719 ^ t43719;
    wire t43721 = t43720 ^ t43720;
    wire t43722 = t43721 ^ t43721;
    wire t43723 = t43722 ^ t43722;
    wire t43724 = t43723 ^ t43723;
    wire t43725 = t43724 ^ t43724;
    wire t43726 = t43725 ^ t43725;
    wire t43727 = t43726 ^ t43726;
    wire t43728 = t43727 ^ t43727;
    wire t43729 = t43728 ^ t43728;
    wire t43730 = t43729 ^ t43729;
    wire t43731 = t43730 ^ t43730;
    wire t43732 = t43731 ^ t43731;
    wire t43733 = t43732 ^ t43732;
    wire t43734 = t43733 ^ t43733;
    wire t43735 = t43734 ^ t43734;
    wire t43736 = t43735 ^ t43735;
    wire t43737 = t43736 ^ t43736;
    wire t43738 = t43737 ^ t43737;
    wire t43739 = t43738 ^ t43738;
    wire t43740 = t43739 ^ t43739;
    wire t43741 = t43740 ^ t43740;
    wire t43742 = t43741 ^ t43741;
    wire t43743 = t43742 ^ t43742;
    wire t43744 = t43743 ^ t43743;
    wire t43745 = t43744 ^ t43744;
    wire t43746 = t43745 ^ t43745;
    wire t43747 = t43746 ^ t43746;
    wire t43748 = t43747 ^ t43747;
    wire t43749 = t43748 ^ t43748;
    wire t43750 = t43749 ^ t43749;
    wire t43751 = t43750 ^ t43750;
    wire t43752 = t43751 ^ t43751;
    wire t43753 = t43752 ^ t43752;
    wire t43754 = t43753 ^ t43753;
    wire t43755 = t43754 ^ t43754;
    wire t43756 = t43755 ^ t43755;
    wire t43757 = t43756 ^ t43756;
    wire t43758 = t43757 ^ t43757;
    wire t43759 = t43758 ^ t43758;
    wire t43760 = t43759 ^ t43759;
    wire t43761 = t43760 ^ t43760;
    wire t43762 = t43761 ^ t43761;
    wire t43763 = t43762 ^ t43762;
    wire t43764 = t43763 ^ t43763;
    wire t43765 = t43764 ^ t43764;
    wire t43766 = t43765 ^ t43765;
    wire t43767 = t43766 ^ t43766;
    wire t43768 = t43767 ^ t43767;
    wire t43769 = t43768 ^ t43768;
    wire t43770 = t43769 ^ t43769;
    wire t43771 = t43770 ^ t43770;
    wire t43772 = t43771 ^ t43771;
    wire t43773 = t43772 ^ t43772;
    wire t43774 = t43773 ^ t43773;
    wire t43775 = t43774 ^ t43774;
    wire t43776 = t43775 ^ t43775;
    wire t43777 = t43776 ^ t43776;
    wire t43778 = t43777 ^ t43777;
    wire t43779 = t43778 ^ t43778;
    wire t43780 = t43779 ^ t43779;
    wire t43781 = t43780 ^ t43780;
    wire t43782 = t43781 ^ t43781;
    wire t43783 = t43782 ^ t43782;
    wire t43784 = t43783 ^ t43783;
    wire t43785 = t43784 ^ t43784;
    wire t43786 = t43785 ^ t43785;
    wire t43787 = t43786 ^ t43786;
    wire t43788 = t43787 ^ t43787;
    wire t43789 = t43788 ^ t43788;
    wire t43790 = t43789 ^ t43789;
    wire t43791 = t43790 ^ t43790;
    wire t43792 = t43791 ^ t43791;
    wire t43793 = t43792 ^ t43792;
    wire t43794 = t43793 ^ t43793;
    wire t43795 = t43794 ^ t43794;
    wire t43796 = t43795 ^ t43795;
    wire t43797 = t43796 ^ t43796;
    wire t43798 = t43797 ^ t43797;
    wire t43799 = t43798 ^ t43798;
    wire t43800 = t43799 ^ t43799;
    wire t43801 = t43800 ^ t43800;
    wire t43802 = t43801 ^ t43801;
    wire t43803 = t43802 ^ t43802;
    wire t43804 = t43803 ^ t43803;
    wire t43805 = t43804 ^ t43804;
    wire t43806 = t43805 ^ t43805;
    wire t43807 = t43806 ^ t43806;
    wire t43808 = t43807 ^ t43807;
    wire t43809 = t43808 ^ t43808;
    wire t43810 = t43809 ^ t43809;
    wire t43811 = t43810 ^ t43810;
    wire t43812 = t43811 ^ t43811;
    wire t43813 = t43812 ^ t43812;
    wire t43814 = t43813 ^ t43813;
    wire t43815 = t43814 ^ t43814;
    wire t43816 = t43815 ^ t43815;
    wire t43817 = t43816 ^ t43816;
    wire t43818 = t43817 ^ t43817;
    wire t43819 = t43818 ^ t43818;
    wire t43820 = t43819 ^ t43819;
    wire t43821 = t43820 ^ t43820;
    wire t43822 = t43821 ^ t43821;
    wire t43823 = t43822 ^ t43822;
    wire t43824 = t43823 ^ t43823;
    wire t43825 = t43824 ^ t43824;
    wire t43826 = t43825 ^ t43825;
    wire t43827 = t43826 ^ t43826;
    wire t43828 = t43827 ^ t43827;
    wire t43829 = t43828 ^ t43828;
    wire t43830 = t43829 ^ t43829;
    wire t43831 = t43830 ^ t43830;
    wire t43832 = t43831 ^ t43831;
    wire t43833 = t43832 ^ t43832;
    wire t43834 = t43833 ^ t43833;
    wire t43835 = t43834 ^ t43834;
    wire t43836 = t43835 ^ t43835;
    wire t43837 = t43836 ^ t43836;
    wire t43838 = t43837 ^ t43837;
    wire t43839 = t43838 ^ t43838;
    wire t43840 = t43839 ^ t43839;
    wire t43841 = t43840 ^ t43840;
    wire t43842 = t43841 ^ t43841;
    wire t43843 = t43842 ^ t43842;
    wire t43844 = t43843 ^ t43843;
    wire t43845 = t43844 ^ t43844;
    wire t43846 = t43845 ^ t43845;
    wire t43847 = t43846 ^ t43846;
    wire t43848 = t43847 ^ t43847;
    wire t43849 = t43848 ^ t43848;
    wire t43850 = t43849 ^ t43849;
    wire t43851 = t43850 ^ t43850;
    wire t43852 = t43851 ^ t43851;
    wire t43853 = t43852 ^ t43852;
    wire t43854 = t43853 ^ t43853;
    wire t43855 = t43854 ^ t43854;
    wire t43856 = t43855 ^ t43855;
    wire t43857 = t43856 ^ t43856;
    wire t43858 = t43857 ^ t43857;
    wire t43859 = t43858 ^ t43858;
    wire t43860 = t43859 ^ t43859;
    wire t43861 = t43860 ^ t43860;
    wire t43862 = t43861 ^ t43861;
    wire t43863 = t43862 ^ t43862;
    wire t43864 = t43863 ^ t43863;
    wire t43865 = t43864 ^ t43864;
    wire t43866 = t43865 ^ t43865;
    wire t43867 = t43866 ^ t43866;
    wire t43868 = t43867 ^ t43867;
    wire t43869 = t43868 ^ t43868;
    wire t43870 = t43869 ^ t43869;
    wire t43871 = t43870 ^ t43870;
    wire t43872 = t43871 ^ t43871;
    wire t43873 = t43872 ^ t43872;
    wire t43874 = t43873 ^ t43873;
    wire t43875 = t43874 ^ t43874;
    wire t43876 = t43875 ^ t43875;
    wire t43877 = t43876 ^ t43876;
    wire t43878 = t43877 ^ t43877;
    wire t43879 = t43878 ^ t43878;
    wire t43880 = t43879 ^ t43879;
    wire t43881 = t43880 ^ t43880;
    wire t43882 = t43881 ^ t43881;
    wire t43883 = t43882 ^ t43882;
    wire t43884 = t43883 ^ t43883;
    wire t43885 = t43884 ^ t43884;
    wire t43886 = t43885 ^ t43885;
    wire t43887 = t43886 ^ t43886;
    wire t43888 = t43887 ^ t43887;
    wire t43889 = t43888 ^ t43888;
    wire t43890 = t43889 ^ t43889;
    wire t43891 = t43890 ^ t43890;
    wire t43892 = t43891 ^ t43891;
    wire t43893 = t43892 ^ t43892;
    wire t43894 = t43893 ^ t43893;
    wire t43895 = t43894 ^ t43894;
    wire t43896 = t43895 ^ t43895;
    wire t43897 = t43896 ^ t43896;
    wire t43898 = t43897 ^ t43897;
    wire t43899 = t43898 ^ t43898;
    wire t43900 = t43899 ^ t43899;
    wire t43901 = t43900 ^ t43900;
    wire t43902 = t43901 ^ t43901;
    wire t43903 = t43902 ^ t43902;
    wire t43904 = t43903 ^ t43903;
    wire t43905 = t43904 ^ t43904;
    wire t43906 = t43905 ^ t43905;
    wire t43907 = t43906 ^ t43906;
    wire t43908 = t43907 ^ t43907;
    wire t43909 = t43908 ^ t43908;
    wire t43910 = t43909 ^ t43909;
    wire t43911 = t43910 ^ t43910;
    wire t43912 = t43911 ^ t43911;
    wire t43913 = t43912 ^ t43912;
    wire t43914 = t43913 ^ t43913;
    wire t43915 = t43914 ^ t43914;
    wire t43916 = t43915 ^ t43915;
    wire t43917 = t43916 ^ t43916;
    wire t43918 = t43917 ^ t43917;
    wire t43919 = t43918 ^ t43918;
    wire t43920 = t43919 ^ t43919;
    wire t43921 = t43920 ^ t43920;
    wire t43922 = t43921 ^ t43921;
    wire t43923 = t43922 ^ t43922;
    wire t43924 = t43923 ^ t43923;
    wire t43925 = t43924 ^ t43924;
    wire t43926 = t43925 ^ t43925;
    wire t43927 = t43926 ^ t43926;
    wire t43928 = t43927 ^ t43927;
    wire t43929 = t43928 ^ t43928;
    wire t43930 = t43929 ^ t43929;
    wire t43931 = t43930 ^ t43930;
    wire t43932 = t43931 ^ t43931;
    wire t43933 = t43932 ^ t43932;
    wire t43934 = t43933 ^ t43933;
    wire t43935 = t43934 ^ t43934;
    wire t43936 = t43935 ^ t43935;
    wire t43937 = t43936 ^ t43936;
    wire t43938 = t43937 ^ t43937;
    wire t43939 = t43938 ^ t43938;
    wire t43940 = t43939 ^ t43939;
    wire t43941 = t43940 ^ t43940;
    wire t43942 = t43941 ^ t43941;
    wire t43943 = t43942 ^ t43942;
    wire t43944 = t43943 ^ t43943;
    wire t43945 = t43944 ^ t43944;
    wire t43946 = t43945 ^ t43945;
    wire t43947 = t43946 ^ t43946;
    wire t43948 = t43947 ^ t43947;
    wire t43949 = t43948 ^ t43948;
    wire t43950 = t43949 ^ t43949;
    wire t43951 = t43950 ^ t43950;
    wire t43952 = t43951 ^ t43951;
    wire t43953 = t43952 ^ t43952;
    wire t43954 = t43953 ^ t43953;
    wire t43955 = t43954 ^ t43954;
    wire t43956 = t43955 ^ t43955;
    wire t43957 = t43956 ^ t43956;
    wire t43958 = t43957 ^ t43957;
    wire t43959 = t43958 ^ t43958;
    wire t43960 = t43959 ^ t43959;
    wire t43961 = t43960 ^ t43960;
    wire t43962 = t43961 ^ t43961;
    wire t43963 = t43962 ^ t43962;
    wire t43964 = t43963 ^ t43963;
    wire t43965 = t43964 ^ t43964;
    wire t43966 = t43965 ^ t43965;
    wire t43967 = t43966 ^ t43966;
    wire t43968 = t43967 ^ t43967;
    wire t43969 = t43968 ^ t43968;
    wire t43970 = t43969 ^ t43969;
    wire t43971 = t43970 ^ t43970;
    wire t43972 = t43971 ^ t43971;
    wire t43973 = t43972 ^ t43972;
    wire t43974 = t43973 ^ t43973;
    wire t43975 = t43974 ^ t43974;
    wire t43976 = t43975 ^ t43975;
    wire t43977 = t43976 ^ t43976;
    wire t43978 = t43977 ^ t43977;
    wire t43979 = t43978 ^ t43978;
    wire t43980 = t43979 ^ t43979;
    wire t43981 = t43980 ^ t43980;
    wire t43982 = t43981 ^ t43981;
    wire t43983 = t43982 ^ t43982;
    wire t43984 = t43983 ^ t43983;
    wire t43985 = t43984 ^ t43984;
    wire t43986 = t43985 ^ t43985;
    wire t43987 = t43986 ^ t43986;
    wire t43988 = t43987 ^ t43987;
    wire t43989 = t43988 ^ t43988;
    wire t43990 = t43989 ^ t43989;
    wire t43991 = t43990 ^ t43990;
    wire t43992 = t43991 ^ t43991;
    wire t43993 = t43992 ^ t43992;
    wire t43994 = t43993 ^ t43993;
    wire t43995 = t43994 ^ t43994;
    wire t43996 = t43995 ^ t43995;
    wire t43997 = t43996 ^ t43996;
    wire t43998 = t43997 ^ t43997;
    wire t43999 = t43998 ^ t43998;
    wire t44000 = t43999 ^ t43999;
    wire t44001 = t44000 ^ t44000;
    wire t44002 = t44001 ^ t44001;
    wire t44003 = t44002 ^ t44002;
    wire t44004 = t44003 ^ t44003;
    wire t44005 = t44004 ^ t44004;
    wire t44006 = t44005 ^ t44005;
    wire t44007 = t44006 ^ t44006;
    wire t44008 = t44007 ^ t44007;
    wire t44009 = t44008 ^ t44008;
    wire t44010 = t44009 ^ t44009;
    wire t44011 = t44010 ^ t44010;
    wire t44012 = t44011 ^ t44011;
    wire t44013 = t44012 ^ t44012;
    wire t44014 = t44013 ^ t44013;
    wire t44015 = t44014 ^ t44014;
    wire t44016 = t44015 ^ t44015;
    wire t44017 = t44016 ^ t44016;
    wire t44018 = t44017 ^ t44017;
    wire t44019 = t44018 ^ t44018;
    wire t44020 = t44019 ^ t44019;
    wire t44021 = t44020 ^ t44020;
    wire t44022 = t44021 ^ t44021;
    wire t44023 = t44022 ^ t44022;
    wire t44024 = t44023 ^ t44023;
    wire t44025 = t44024 ^ t44024;
    wire t44026 = t44025 ^ t44025;
    wire t44027 = t44026 ^ t44026;
    wire t44028 = t44027 ^ t44027;
    wire t44029 = t44028 ^ t44028;
    wire t44030 = t44029 ^ t44029;
    wire t44031 = t44030 ^ t44030;
    wire t44032 = t44031 ^ t44031;
    wire t44033 = t44032 ^ t44032;
    wire t44034 = t44033 ^ t44033;
    wire t44035 = t44034 ^ t44034;
    wire t44036 = t44035 ^ t44035;
    wire t44037 = t44036 ^ t44036;
    wire t44038 = t44037 ^ t44037;
    wire t44039 = t44038 ^ t44038;
    wire t44040 = t44039 ^ t44039;
    wire t44041 = t44040 ^ t44040;
    wire t44042 = t44041 ^ t44041;
    wire t44043 = t44042 ^ t44042;
    wire t44044 = t44043 ^ t44043;
    wire t44045 = t44044 ^ t44044;
    wire t44046 = t44045 ^ t44045;
    wire t44047 = t44046 ^ t44046;
    wire t44048 = t44047 ^ t44047;
    wire t44049 = t44048 ^ t44048;
    wire t44050 = t44049 ^ t44049;
    wire t44051 = t44050 ^ t44050;
    wire t44052 = t44051 ^ t44051;
    wire t44053 = t44052 ^ t44052;
    wire t44054 = t44053 ^ t44053;
    wire t44055 = t44054 ^ t44054;
    wire t44056 = t44055 ^ t44055;
    wire t44057 = t44056 ^ t44056;
    wire t44058 = t44057 ^ t44057;
    wire t44059 = t44058 ^ t44058;
    wire t44060 = t44059 ^ t44059;
    wire t44061 = t44060 ^ t44060;
    wire t44062 = t44061 ^ t44061;
    wire t44063 = t44062 ^ t44062;
    wire t44064 = t44063 ^ t44063;
    wire t44065 = t44064 ^ t44064;
    wire t44066 = t44065 ^ t44065;
    wire t44067 = t44066 ^ t44066;
    wire t44068 = t44067 ^ t44067;
    wire t44069 = t44068 ^ t44068;
    wire t44070 = t44069 ^ t44069;
    wire t44071 = t44070 ^ t44070;
    wire t44072 = t44071 ^ t44071;
    wire t44073 = t44072 ^ t44072;
    wire t44074 = t44073 ^ t44073;
    wire t44075 = t44074 ^ t44074;
    wire t44076 = t44075 ^ t44075;
    wire t44077 = t44076 ^ t44076;
    wire t44078 = t44077 ^ t44077;
    wire t44079 = t44078 ^ t44078;
    wire t44080 = t44079 ^ t44079;
    wire t44081 = t44080 ^ t44080;
    wire t44082 = t44081 ^ t44081;
    wire t44083 = t44082 ^ t44082;
    wire t44084 = t44083 ^ t44083;
    wire t44085 = t44084 ^ t44084;
    wire t44086 = t44085 ^ t44085;
    wire t44087 = t44086 ^ t44086;
    wire t44088 = t44087 ^ t44087;
    wire t44089 = t44088 ^ t44088;
    wire t44090 = t44089 ^ t44089;
    wire t44091 = t44090 ^ t44090;
    wire t44092 = t44091 ^ t44091;
    wire t44093 = t44092 ^ t44092;
    wire t44094 = t44093 ^ t44093;
    wire t44095 = t44094 ^ t44094;
    wire t44096 = t44095 ^ t44095;
    wire t44097 = t44096 ^ t44096;
    wire t44098 = t44097 ^ t44097;
    wire t44099 = t44098 ^ t44098;
    wire t44100 = t44099 ^ t44099;
    wire t44101 = t44100 ^ t44100;
    wire t44102 = t44101 ^ t44101;
    wire t44103 = t44102 ^ t44102;
    wire t44104 = t44103 ^ t44103;
    wire t44105 = t44104 ^ t44104;
    wire t44106 = t44105 ^ t44105;
    wire t44107 = t44106 ^ t44106;
    wire t44108 = t44107 ^ t44107;
    wire t44109 = t44108 ^ t44108;
    wire t44110 = t44109 ^ t44109;
    wire t44111 = t44110 ^ t44110;
    wire t44112 = t44111 ^ t44111;
    wire t44113 = t44112 ^ t44112;
    wire t44114 = t44113 ^ t44113;
    wire t44115 = t44114 ^ t44114;
    wire t44116 = t44115 ^ t44115;
    wire t44117 = t44116 ^ t44116;
    wire t44118 = t44117 ^ t44117;
    wire t44119 = t44118 ^ t44118;
    wire t44120 = t44119 ^ t44119;
    wire t44121 = t44120 ^ t44120;
    wire t44122 = t44121 ^ t44121;
    wire t44123 = t44122 ^ t44122;
    wire t44124 = t44123 ^ t44123;
    wire t44125 = t44124 ^ t44124;
    wire t44126 = t44125 ^ t44125;
    wire t44127 = t44126 ^ t44126;
    wire t44128 = t44127 ^ t44127;
    wire t44129 = t44128 ^ t44128;
    wire t44130 = t44129 ^ t44129;
    wire t44131 = t44130 ^ t44130;
    wire t44132 = t44131 ^ t44131;
    wire t44133 = t44132 ^ t44132;
    wire t44134 = t44133 ^ t44133;
    wire t44135 = t44134 ^ t44134;
    wire t44136 = t44135 ^ t44135;
    wire t44137 = t44136 ^ t44136;
    wire t44138 = t44137 ^ t44137;
    wire t44139 = t44138 ^ t44138;
    wire t44140 = t44139 ^ t44139;
    wire t44141 = t44140 ^ t44140;
    wire t44142 = t44141 ^ t44141;
    wire t44143 = t44142 ^ t44142;
    wire t44144 = t44143 ^ t44143;
    wire t44145 = t44144 ^ t44144;
    wire t44146 = t44145 ^ t44145;
    wire t44147 = t44146 ^ t44146;
    wire t44148 = t44147 ^ t44147;
    wire t44149 = t44148 ^ t44148;
    wire t44150 = t44149 ^ t44149;
    wire t44151 = t44150 ^ t44150;
    wire t44152 = t44151 ^ t44151;
    wire t44153 = t44152 ^ t44152;
    wire t44154 = t44153 ^ t44153;
    wire t44155 = t44154 ^ t44154;
    wire t44156 = t44155 ^ t44155;
    wire t44157 = t44156 ^ t44156;
    wire t44158 = t44157 ^ t44157;
    wire t44159 = t44158 ^ t44158;
    wire t44160 = t44159 ^ t44159;
    wire t44161 = t44160 ^ t44160;
    wire t44162 = t44161 ^ t44161;
    wire t44163 = t44162 ^ t44162;
    wire t44164 = t44163 ^ t44163;
    wire t44165 = t44164 ^ t44164;
    wire t44166 = t44165 ^ t44165;
    wire t44167 = t44166 ^ t44166;
    wire t44168 = t44167 ^ t44167;
    wire t44169 = t44168 ^ t44168;
    wire t44170 = t44169 ^ t44169;
    wire t44171 = t44170 ^ t44170;
    wire t44172 = t44171 ^ t44171;
    wire t44173 = t44172 ^ t44172;
    wire t44174 = t44173 ^ t44173;
    wire t44175 = t44174 ^ t44174;
    wire t44176 = t44175 ^ t44175;
    wire t44177 = t44176 ^ t44176;
    wire t44178 = t44177 ^ t44177;
    wire t44179 = t44178 ^ t44178;
    wire t44180 = t44179 ^ t44179;
    wire t44181 = t44180 ^ t44180;
    wire t44182 = t44181 ^ t44181;
    wire t44183 = t44182 ^ t44182;
    wire t44184 = t44183 ^ t44183;
    wire t44185 = t44184 ^ t44184;
    wire t44186 = t44185 ^ t44185;
    wire t44187 = t44186 ^ t44186;
    wire t44188 = t44187 ^ t44187;
    wire t44189 = t44188 ^ t44188;
    wire t44190 = t44189 ^ t44189;
    wire t44191 = t44190 ^ t44190;
    wire t44192 = t44191 ^ t44191;
    wire t44193 = t44192 ^ t44192;
    wire t44194 = t44193 ^ t44193;
    wire t44195 = t44194 ^ t44194;
    wire t44196 = t44195 ^ t44195;
    wire t44197 = t44196 ^ t44196;
    wire t44198 = t44197 ^ t44197;
    wire t44199 = t44198 ^ t44198;
    wire t44200 = t44199 ^ t44199;
    wire t44201 = t44200 ^ t44200;
    wire t44202 = t44201 ^ t44201;
    wire t44203 = t44202 ^ t44202;
    wire t44204 = t44203 ^ t44203;
    wire t44205 = t44204 ^ t44204;
    wire t44206 = t44205 ^ t44205;
    wire t44207 = t44206 ^ t44206;
    wire t44208 = t44207 ^ t44207;
    wire t44209 = t44208 ^ t44208;
    wire t44210 = t44209 ^ t44209;
    wire t44211 = t44210 ^ t44210;
    wire t44212 = t44211 ^ t44211;
    wire t44213 = t44212 ^ t44212;
    wire t44214 = t44213 ^ t44213;
    wire t44215 = t44214 ^ t44214;
    wire t44216 = t44215 ^ t44215;
    wire t44217 = t44216 ^ t44216;
    wire t44218 = t44217 ^ t44217;
    wire t44219 = t44218 ^ t44218;
    wire t44220 = t44219 ^ t44219;
    wire t44221 = t44220 ^ t44220;
    wire t44222 = t44221 ^ t44221;
    wire t44223 = t44222 ^ t44222;
    wire t44224 = t44223 ^ t44223;
    wire t44225 = t44224 ^ t44224;
    wire t44226 = t44225 ^ t44225;
    wire t44227 = t44226 ^ t44226;
    wire t44228 = t44227 ^ t44227;
    wire t44229 = t44228 ^ t44228;
    wire t44230 = t44229 ^ t44229;
    wire t44231 = t44230 ^ t44230;
    wire t44232 = t44231 ^ t44231;
    wire t44233 = t44232 ^ t44232;
    wire t44234 = t44233 ^ t44233;
    wire t44235 = t44234 ^ t44234;
    wire t44236 = t44235 ^ t44235;
    wire t44237 = t44236 ^ t44236;
    wire t44238 = t44237 ^ t44237;
    wire t44239 = t44238 ^ t44238;
    wire t44240 = t44239 ^ t44239;
    wire t44241 = t44240 ^ t44240;
    wire t44242 = t44241 ^ t44241;
    wire t44243 = t44242 ^ t44242;
    wire t44244 = t44243 ^ t44243;
    wire t44245 = t44244 ^ t44244;
    wire t44246 = t44245 ^ t44245;
    wire t44247 = t44246 ^ t44246;
    wire t44248 = t44247 ^ t44247;
    wire t44249 = t44248 ^ t44248;
    wire t44250 = t44249 ^ t44249;
    wire t44251 = t44250 ^ t44250;
    wire t44252 = t44251 ^ t44251;
    wire t44253 = t44252 ^ t44252;
    wire t44254 = t44253 ^ t44253;
    wire t44255 = t44254 ^ t44254;
    wire t44256 = t44255 ^ t44255;
    wire t44257 = t44256 ^ t44256;
    wire t44258 = t44257 ^ t44257;
    wire t44259 = t44258 ^ t44258;
    wire t44260 = t44259 ^ t44259;
    wire t44261 = t44260 ^ t44260;
    wire t44262 = t44261 ^ t44261;
    wire t44263 = t44262 ^ t44262;
    wire t44264 = t44263 ^ t44263;
    wire t44265 = t44264 ^ t44264;
    wire t44266 = t44265 ^ t44265;
    wire t44267 = t44266 ^ t44266;
    wire t44268 = t44267 ^ t44267;
    wire t44269 = t44268 ^ t44268;
    wire t44270 = t44269 ^ t44269;
    wire t44271 = t44270 ^ t44270;
    wire t44272 = t44271 ^ t44271;
    wire t44273 = t44272 ^ t44272;
    wire t44274 = t44273 ^ t44273;
    wire t44275 = t44274 ^ t44274;
    wire t44276 = t44275 ^ t44275;
    wire t44277 = t44276 ^ t44276;
    wire t44278 = t44277 ^ t44277;
    wire t44279 = t44278 ^ t44278;
    wire t44280 = t44279 ^ t44279;
    wire t44281 = t44280 ^ t44280;
    wire t44282 = t44281 ^ t44281;
    wire t44283 = t44282 ^ t44282;
    wire t44284 = t44283 ^ t44283;
    wire t44285 = t44284 ^ t44284;
    wire t44286 = t44285 ^ t44285;
    wire t44287 = t44286 ^ t44286;
    wire t44288 = t44287 ^ t44287;
    wire t44289 = t44288 ^ t44288;
    wire t44290 = t44289 ^ t44289;
    wire t44291 = t44290 ^ t44290;
    wire t44292 = t44291 ^ t44291;
    wire t44293 = t44292 ^ t44292;
    wire t44294 = t44293 ^ t44293;
    wire t44295 = t44294 ^ t44294;
    wire t44296 = t44295 ^ t44295;
    wire t44297 = t44296 ^ t44296;
    wire t44298 = t44297 ^ t44297;
    wire t44299 = t44298 ^ t44298;
    wire t44300 = t44299 ^ t44299;
    wire t44301 = t44300 ^ t44300;
    wire t44302 = t44301 ^ t44301;
    wire t44303 = t44302 ^ t44302;
    wire t44304 = t44303 ^ t44303;
    wire t44305 = t44304 ^ t44304;
    wire t44306 = t44305 ^ t44305;
    wire t44307 = t44306 ^ t44306;
    wire t44308 = t44307 ^ t44307;
    wire t44309 = t44308 ^ t44308;
    wire t44310 = t44309 ^ t44309;
    wire t44311 = t44310 ^ t44310;
    wire t44312 = t44311 ^ t44311;
    wire t44313 = t44312 ^ t44312;
    wire t44314 = t44313 ^ t44313;
    wire t44315 = t44314 ^ t44314;
    wire t44316 = t44315 ^ t44315;
    wire t44317 = t44316 ^ t44316;
    wire t44318 = t44317 ^ t44317;
    wire t44319 = t44318 ^ t44318;
    wire t44320 = t44319 ^ t44319;
    wire t44321 = t44320 ^ t44320;
    wire t44322 = t44321 ^ t44321;
    wire t44323 = t44322 ^ t44322;
    wire t44324 = t44323 ^ t44323;
    wire t44325 = t44324 ^ t44324;
    wire t44326 = t44325 ^ t44325;
    wire t44327 = t44326 ^ t44326;
    wire t44328 = t44327 ^ t44327;
    wire t44329 = t44328 ^ t44328;
    wire t44330 = t44329 ^ t44329;
    wire t44331 = t44330 ^ t44330;
    wire t44332 = t44331 ^ t44331;
    wire t44333 = t44332 ^ t44332;
    wire t44334 = t44333 ^ t44333;
    wire t44335 = t44334 ^ t44334;
    wire t44336 = t44335 ^ t44335;
    wire t44337 = t44336 ^ t44336;
    wire t44338 = t44337 ^ t44337;
    wire t44339 = t44338 ^ t44338;
    wire t44340 = t44339 ^ t44339;
    wire t44341 = t44340 ^ t44340;
    wire t44342 = t44341 ^ t44341;
    wire t44343 = t44342 ^ t44342;
    wire t44344 = t44343 ^ t44343;
    wire t44345 = t44344 ^ t44344;
    wire t44346 = t44345 ^ t44345;
    wire t44347 = t44346 ^ t44346;
    wire t44348 = t44347 ^ t44347;
    wire t44349 = t44348 ^ t44348;
    wire t44350 = t44349 ^ t44349;
    wire t44351 = t44350 ^ t44350;
    wire t44352 = t44351 ^ t44351;
    wire t44353 = t44352 ^ t44352;
    wire t44354 = t44353 ^ t44353;
    wire t44355 = t44354 ^ t44354;
    wire t44356 = t44355 ^ t44355;
    wire t44357 = t44356 ^ t44356;
    wire t44358 = t44357 ^ t44357;
    wire t44359 = t44358 ^ t44358;
    wire t44360 = t44359 ^ t44359;
    wire t44361 = t44360 ^ t44360;
    wire t44362 = t44361 ^ t44361;
    wire t44363 = t44362 ^ t44362;
    wire t44364 = t44363 ^ t44363;
    wire t44365 = t44364 ^ t44364;
    wire t44366 = t44365 ^ t44365;
    wire t44367 = t44366 ^ t44366;
    wire t44368 = t44367 ^ t44367;
    wire t44369 = t44368 ^ t44368;
    wire t44370 = t44369 ^ t44369;
    wire t44371 = t44370 ^ t44370;
    wire t44372 = t44371 ^ t44371;
    wire t44373 = t44372 ^ t44372;
    wire t44374 = t44373 ^ t44373;
    wire t44375 = t44374 ^ t44374;
    wire t44376 = t44375 ^ t44375;
    wire t44377 = t44376 ^ t44376;
    wire t44378 = t44377 ^ t44377;
    wire t44379 = t44378 ^ t44378;
    wire t44380 = t44379 ^ t44379;
    wire t44381 = t44380 ^ t44380;
    wire t44382 = t44381 ^ t44381;
    wire t44383 = t44382 ^ t44382;
    wire t44384 = t44383 ^ t44383;
    wire t44385 = t44384 ^ t44384;
    wire t44386 = t44385 ^ t44385;
    wire t44387 = t44386 ^ t44386;
    wire t44388 = t44387 ^ t44387;
    wire t44389 = t44388 ^ t44388;
    wire t44390 = t44389 ^ t44389;
    wire t44391 = t44390 ^ t44390;
    wire t44392 = t44391 ^ t44391;
    wire t44393 = t44392 ^ t44392;
    wire t44394 = t44393 ^ t44393;
    wire t44395 = t44394 ^ t44394;
    wire t44396 = t44395 ^ t44395;
    wire t44397 = t44396 ^ t44396;
    wire t44398 = t44397 ^ t44397;
    wire t44399 = t44398 ^ t44398;
    wire t44400 = t44399 ^ t44399;
    wire t44401 = t44400 ^ t44400;
    wire t44402 = t44401 ^ t44401;
    wire t44403 = t44402 ^ t44402;
    wire t44404 = t44403 ^ t44403;
    wire t44405 = t44404 ^ t44404;
    wire t44406 = t44405 ^ t44405;
    wire t44407 = t44406 ^ t44406;
    wire t44408 = t44407 ^ t44407;
    wire t44409 = t44408 ^ t44408;
    wire t44410 = t44409 ^ t44409;
    wire t44411 = t44410 ^ t44410;
    wire t44412 = t44411 ^ t44411;
    wire t44413 = t44412 ^ t44412;
    wire t44414 = t44413 ^ t44413;
    wire t44415 = t44414 ^ t44414;
    wire t44416 = t44415 ^ t44415;
    wire t44417 = t44416 ^ t44416;
    wire t44418 = t44417 ^ t44417;
    wire t44419 = t44418 ^ t44418;
    wire t44420 = t44419 ^ t44419;
    wire t44421 = t44420 ^ t44420;
    wire t44422 = t44421 ^ t44421;
    wire t44423 = t44422 ^ t44422;
    wire t44424 = t44423 ^ t44423;
    wire t44425 = t44424 ^ t44424;
    wire t44426 = t44425 ^ t44425;
    wire t44427 = t44426 ^ t44426;
    wire t44428 = t44427 ^ t44427;
    wire t44429 = t44428 ^ t44428;
    wire t44430 = t44429 ^ t44429;
    wire t44431 = t44430 ^ t44430;
    wire t44432 = t44431 ^ t44431;
    wire t44433 = t44432 ^ t44432;
    wire t44434 = t44433 ^ t44433;
    wire t44435 = t44434 ^ t44434;
    wire t44436 = t44435 ^ t44435;
    wire t44437 = t44436 ^ t44436;
    wire t44438 = t44437 ^ t44437;
    wire t44439 = t44438 ^ t44438;
    wire t44440 = t44439 ^ t44439;
    wire t44441 = t44440 ^ t44440;
    wire t44442 = t44441 ^ t44441;
    wire t44443 = t44442 ^ t44442;
    wire t44444 = t44443 ^ t44443;
    wire t44445 = t44444 ^ t44444;
    wire t44446 = t44445 ^ t44445;
    wire t44447 = t44446 ^ t44446;
    wire t44448 = t44447 ^ t44447;
    wire t44449 = t44448 ^ t44448;
    wire t44450 = t44449 ^ t44449;
    wire t44451 = t44450 ^ t44450;
    wire t44452 = t44451 ^ t44451;
    wire t44453 = t44452 ^ t44452;
    wire t44454 = t44453 ^ t44453;
    wire t44455 = t44454 ^ t44454;
    wire t44456 = t44455 ^ t44455;
    wire t44457 = t44456 ^ t44456;
    wire t44458 = t44457 ^ t44457;
    wire t44459 = t44458 ^ t44458;
    wire t44460 = t44459 ^ t44459;
    wire t44461 = t44460 ^ t44460;
    wire t44462 = t44461 ^ t44461;
    wire t44463 = t44462 ^ t44462;
    wire t44464 = t44463 ^ t44463;
    wire t44465 = t44464 ^ t44464;
    wire t44466 = t44465 ^ t44465;
    wire t44467 = t44466 ^ t44466;
    wire t44468 = t44467 ^ t44467;
    wire t44469 = t44468 ^ t44468;
    wire t44470 = t44469 ^ t44469;
    wire t44471 = t44470 ^ t44470;
    wire t44472 = t44471 ^ t44471;
    wire t44473 = t44472 ^ t44472;
    wire t44474 = t44473 ^ t44473;
    wire t44475 = t44474 ^ t44474;
    wire t44476 = t44475 ^ t44475;
    wire t44477 = t44476 ^ t44476;
    wire t44478 = t44477 ^ t44477;
    wire t44479 = t44478 ^ t44478;
    wire t44480 = t44479 ^ t44479;
    wire t44481 = t44480 ^ t44480;
    wire t44482 = t44481 ^ t44481;
    wire t44483 = t44482 ^ t44482;
    wire t44484 = t44483 ^ t44483;
    wire t44485 = t44484 ^ t44484;
    wire t44486 = t44485 ^ t44485;
    wire t44487 = t44486 ^ t44486;
    wire t44488 = t44487 ^ t44487;
    wire t44489 = t44488 ^ t44488;
    wire t44490 = t44489 ^ t44489;
    wire t44491 = t44490 ^ t44490;
    wire t44492 = t44491 ^ t44491;
    wire t44493 = t44492 ^ t44492;
    wire t44494 = t44493 ^ t44493;
    wire t44495 = t44494 ^ t44494;
    wire t44496 = t44495 ^ t44495;
    wire t44497 = t44496 ^ t44496;
    wire t44498 = t44497 ^ t44497;
    wire t44499 = t44498 ^ t44498;
    wire t44500 = t44499 ^ t44499;
    wire t44501 = t44500 ^ t44500;
    wire t44502 = t44501 ^ t44501;
    wire t44503 = t44502 ^ t44502;
    wire t44504 = t44503 ^ t44503;
    wire t44505 = t44504 ^ t44504;
    wire t44506 = t44505 ^ t44505;
    wire t44507 = t44506 ^ t44506;
    wire t44508 = t44507 ^ t44507;
    wire t44509 = t44508 ^ t44508;
    wire t44510 = t44509 ^ t44509;
    wire t44511 = t44510 ^ t44510;
    wire t44512 = t44511 ^ t44511;
    wire t44513 = t44512 ^ t44512;
    wire t44514 = t44513 ^ t44513;
    wire t44515 = t44514 ^ t44514;
    wire t44516 = t44515 ^ t44515;
    wire t44517 = t44516 ^ t44516;
    wire t44518 = t44517 ^ t44517;
    wire t44519 = t44518 ^ t44518;
    wire t44520 = t44519 ^ t44519;
    wire t44521 = t44520 ^ t44520;
    wire t44522 = t44521 ^ t44521;
    wire t44523 = t44522 ^ t44522;
    wire t44524 = t44523 ^ t44523;
    wire t44525 = t44524 ^ t44524;
    wire t44526 = t44525 ^ t44525;
    wire t44527 = t44526 ^ t44526;
    wire t44528 = t44527 ^ t44527;
    wire t44529 = t44528 ^ t44528;
    wire t44530 = t44529 ^ t44529;
    wire t44531 = t44530 ^ t44530;
    wire t44532 = t44531 ^ t44531;
    wire t44533 = t44532 ^ t44532;
    wire t44534 = t44533 ^ t44533;
    wire t44535 = t44534 ^ t44534;
    wire t44536 = t44535 ^ t44535;
    wire t44537 = t44536 ^ t44536;
    wire t44538 = t44537 ^ t44537;
    wire t44539 = t44538 ^ t44538;
    wire t44540 = t44539 ^ t44539;
    wire t44541 = t44540 ^ t44540;
    wire t44542 = t44541 ^ t44541;
    wire t44543 = t44542 ^ t44542;
    wire t44544 = t44543 ^ t44543;
    wire t44545 = t44544 ^ t44544;
    wire t44546 = t44545 ^ t44545;
    wire t44547 = t44546 ^ t44546;
    wire t44548 = t44547 ^ t44547;
    wire t44549 = t44548 ^ t44548;
    wire t44550 = t44549 ^ t44549;
    wire t44551 = t44550 ^ t44550;
    wire t44552 = t44551 ^ t44551;
    wire t44553 = t44552 ^ t44552;
    wire t44554 = t44553 ^ t44553;
    wire t44555 = t44554 ^ t44554;
    wire t44556 = t44555 ^ t44555;
    wire t44557 = t44556 ^ t44556;
    wire t44558 = t44557 ^ t44557;
    wire t44559 = t44558 ^ t44558;
    wire t44560 = t44559 ^ t44559;
    wire t44561 = t44560 ^ t44560;
    wire t44562 = t44561 ^ t44561;
    wire t44563 = t44562 ^ t44562;
    wire t44564 = t44563 ^ t44563;
    wire t44565 = t44564 ^ t44564;
    wire t44566 = t44565 ^ t44565;
    wire t44567 = t44566 ^ t44566;
    wire t44568 = t44567 ^ t44567;
    wire t44569 = t44568 ^ t44568;
    wire t44570 = t44569 ^ t44569;
    wire t44571 = t44570 ^ t44570;
    wire t44572 = t44571 ^ t44571;
    wire t44573 = t44572 ^ t44572;
    wire t44574 = t44573 ^ t44573;
    wire t44575 = t44574 ^ t44574;
    wire t44576 = t44575 ^ t44575;
    wire t44577 = t44576 ^ t44576;
    wire t44578 = t44577 ^ t44577;
    wire t44579 = t44578 ^ t44578;
    wire t44580 = t44579 ^ t44579;
    wire t44581 = t44580 ^ t44580;
    wire t44582 = t44581 ^ t44581;
    wire t44583 = t44582 ^ t44582;
    wire t44584 = t44583 ^ t44583;
    wire t44585 = t44584 ^ t44584;
    wire t44586 = t44585 ^ t44585;
    wire t44587 = t44586 ^ t44586;
    wire t44588 = t44587 ^ t44587;
    wire t44589 = t44588 ^ t44588;
    wire t44590 = t44589 ^ t44589;
    wire t44591 = t44590 ^ t44590;
    wire t44592 = t44591 ^ t44591;
    wire t44593 = t44592 ^ t44592;
    wire t44594 = t44593 ^ t44593;
    wire t44595 = t44594 ^ t44594;
    wire t44596 = t44595 ^ t44595;
    wire t44597 = t44596 ^ t44596;
    wire t44598 = t44597 ^ t44597;
    wire t44599 = t44598 ^ t44598;
    wire t44600 = t44599 ^ t44599;
    wire t44601 = t44600 ^ t44600;
    wire t44602 = t44601 ^ t44601;
    wire t44603 = t44602 ^ t44602;
    wire t44604 = t44603 ^ t44603;
    wire t44605 = t44604 ^ t44604;
    wire t44606 = t44605 ^ t44605;
    wire t44607 = t44606 ^ t44606;
    wire t44608 = t44607 ^ t44607;
    wire t44609 = t44608 ^ t44608;
    wire t44610 = t44609 ^ t44609;
    wire t44611 = t44610 ^ t44610;
    wire t44612 = t44611 ^ t44611;
    wire t44613 = t44612 ^ t44612;
    wire t44614 = t44613 ^ t44613;
    wire t44615 = t44614 ^ t44614;
    wire t44616 = t44615 ^ t44615;
    wire t44617 = t44616 ^ t44616;
    wire t44618 = t44617 ^ t44617;
    wire t44619 = t44618 ^ t44618;
    wire t44620 = t44619 ^ t44619;
    wire t44621 = t44620 ^ t44620;
    wire t44622 = t44621 ^ t44621;
    wire t44623 = t44622 ^ t44622;
    wire t44624 = t44623 ^ t44623;
    wire t44625 = t44624 ^ t44624;
    wire t44626 = t44625 ^ t44625;
    wire t44627 = t44626 ^ t44626;
    wire t44628 = t44627 ^ t44627;
    wire t44629 = t44628 ^ t44628;
    wire t44630 = t44629 ^ t44629;
    wire t44631 = t44630 ^ t44630;
    wire t44632 = t44631 ^ t44631;
    wire t44633 = t44632 ^ t44632;
    wire t44634 = t44633 ^ t44633;
    wire t44635 = t44634 ^ t44634;
    wire t44636 = t44635 ^ t44635;
    wire t44637 = t44636 ^ t44636;
    wire t44638 = t44637 ^ t44637;
    wire t44639 = t44638 ^ t44638;
    wire t44640 = t44639 ^ t44639;
    wire t44641 = t44640 ^ t44640;
    wire t44642 = t44641 ^ t44641;
    wire t44643 = t44642 ^ t44642;
    wire t44644 = t44643 ^ t44643;
    wire t44645 = t44644 ^ t44644;
    wire t44646 = t44645 ^ t44645;
    wire t44647 = t44646 ^ t44646;
    wire t44648 = t44647 ^ t44647;
    wire t44649 = t44648 ^ t44648;
    wire t44650 = t44649 ^ t44649;
    wire t44651 = t44650 ^ t44650;
    wire t44652 = t44651 ^ t44651;
    wire t44653 = t44652 ^ t44652;
    wire t44654 = t44653 ^ t44653;
    wire t44655 = t44654 ^ t44654;
    wire t44656 = t44655 ^ t44655;
    wire t44657 = t44656 ^ t44656;
    wire t44658 = t44657 ^ t44657;
    wire t44659 = t44658 ^ t44658;
    wire t44660 = t44659 ^ t44659;
    wire t44661 = t44660 ^ t44660;
    wire t44662 = t44661 ^ t44661;
    wire t44663 = t44662 ^ t44662;
    wire t44664 = t44663 ^ t44663;
    wire t44665 = t44664 ^ t44664;
    wire t44666 = t44665 ^ t44665;
    wire t44667 = t44666 ^ t44666;
    wire t44668 = t44667 ^ t44667;
    wire t44669 = t44668 ^ t44668;
    wire t44670 = t44669 ^ t44669;
    wire t44671 = t44670 ^ t44670;
    wire t44672 = t44671 ^ t44671;
    wire t44673 = t44672 ^ t44672;
    wire t44674 = t44673 ^ t44673;
    wire t44675 = t44674 ^ t44674;
    wire t44676 = t44675 ^ t44675;
    wire t44677 = t44676 ^ t44676;
    wire t44678 = t44677 ^ t44677;
    wire t44679 = t44678 ^ t44678;
    wire t44680 = t44679 ^ t44679;
    wire t44681 = t44680 ^ t44680;
    wire t44682 = t44681 ^ t44681;
    wire t44683 = t44682 ^ t44682;
    wire t44684 = t44683 ^ t44683;
    wire t44685 = t44684 ^ t44684;
    wire t44686 = t44685 ^ t44685;
    wire t44687 = t44686 ^ t44686;
    wire t44688 = t44687 ^ t44687;
    wire t44689 = t44688 ^ t44688;
    wire t44690 = t44689 ^ t44689;
    wire t44691 = t44690 ^ t44690;
    wire t44692 = t44691 ^ t44691;
    wire t44693 = t44692 ^ t44692;
    wire t44694 = t44693 ^ t44693;
    wire t44695 = t44694 ^ t44694;
    wire t44696 = t44695 ^ t44695;
    wire t44697 = t44696 ^ t44696;
    wire t44698 = t44697 ^ t44697;
    wire t44699 = t44698 ^ t44698;
    wire t44700 = t44699 ^ t44699;
    wire t44701 = t44700 ^ t44700;
    wire t44702 = t44701 ^ t44701;
    wire t44703 = t44702 ^ t44702;
    wire t44704 = t44703 ^ t44703;
    wire t44705 = t44704 ^ t44704;
    wire t44706 = t44705 ^ t44705;
    wire t44707 = t44706 ^ t44706;
    wire t44708 = t44707 ^ t44707;
    wire t44709 = t44708 ^ t44708;
    wire t44710 = t44709 ^ t44709;
    wire t44711 = t44710 ^ t44710;
    wire t44712 = t44711 ^ t44711;
    wire t44713 = t44712 ^ t44712;
    wire t44714 = t44713 ^ t44713;
    wire t44715 = t44714 ^ t44714;
    wire t44716 = t44715 ^ t44715;
    wire t44717 = t44716 ^ t44716;
    wire t44718 = t44717 ^ t44717;
    wire t44719 = t44718 ^ t44718;
    wire t44720 = t44719 ^ t44719;
    wire t44721 = t44720 ^ t44720;
    wire t44722 = t44721 ^ t44721;
    wire t44723 = t44722 ^ t44722;
    wire t44724 = t44723 ^ t44723;
    wire t44725 = t44724 ^ t44724;
    wire t44726 = t44725 ^ t44725;
    wire t44727 = t44726 ^ t44726;
    wire t44728 = t44727 ^ t44727;
    wire t44729 = t44728 ^ t44728;
    wire t44730 = t44729 ^ t44729;
    wire t44731 = t44730 ^ t44730;
    wire t44732 = t44731 ^ t44731;
    wire t44733 = t44732 ^ t44732;
    wire t44734 = t44733 ^ t44733;
    wire t44735 = t44734 ^ t44734;
    wire t44736 = t44735 ^ t44735;
    wire t44737 = t44736 ^ t44736;
    wire t44738 = t44737 ^ t44737;
    wire t44739 = t44738 ^ t44738;
    wire t44740 = t44739 ^ t44739;
    wire t44741 = t44740 ^ t44740;
    wire t44742 = t44741 ^ t44741;
    wire t44743 = t44742 ^ t44742;
    wire t44744 = t44743 ^ t44743;
    wire t44745 = t44744 ^ t44744;
    wire t44746 = t44745 ^ t44745;
    wire t44747 = t44746 ^ t44746;
    wire t44748 = t44747 ^ t44747;
    wire t44749 = t44748 ^ t44748;
    wire t44750 = t44749 ^ t44749;
    wire t44751 = t44750 ^ t44750;
    wire t44752 = t44751 ^ t44751;
    wire t44753 = t44752 ^ t44752;
    wire t44754 = t44753 ^ t44753;
    wire t44755 = t44754 ^ t44754;
    wire t44756 = t44755 ^ t44755;
    wire t44757 = t44756 ^ t44756;
    wire t44758 = t44757 ^ t44757;
    wire t44759 = t44758 ^ t44758;
    wire t44760 = t44759 ^ t44759;
    wire t44761 = t44760 ^ t44760;
    wire t44762 = t44761 ^ t44761;
    wire t44763 = t44762 ^ t44762;
    wire t44764 = t44763 ^ t44763;
    wire t44765 = t44764 ^ t44764;
    wire t44766 = t44765 ^ t44765;
    wire t44767 = t44766 ^ t44766;
    wire t44768 = t44767 ^ t44767;
    wire t44769 = t44768 ^ t44768;
    wire t44770 = t44769 ^ t44769;
    wire t44771 = t44770 ^ t44770;
    wire t44772 = t44771 ^ t44771;
    wire t44773 = t44772 ^ t44772;
    wire t44774 = t44773 ^ t44773;
    wire t44775 = t44774 ^ t44774;
    wire t44776 = t44775 ^ t44775;
    wire t44777 = t44776 ^ t44776;
    wire t44778 = t44777 ^ t44777;
    wire t44779 = t44778 ^ t44778;
    wire t44780 = t44779 ^ t44779;
    wire t44781 = t44780 ^ t44780;
    wire t44782 = t44781 ^ t44781;
    wire t44783 = t44782 ^ t44782;
    wire t44784 = t44783 ^ t44783;
    wire t44785 = t44784 ^ t44784;
    wire t44786 = t44785 ^ t44785;
    wire t44787 = t44786 ^ t44786;
    wire t44788 = t44787 ^ t44787;
    wire t44789 = t44788 ^ t44788;
    wire t44790 = t44789 ^ t44789;
    wire t44791 = t44790 ^ t44790;
    wire t44792 = t44791 ^ t44791;
    wire t44793 = t44792 ^ t44792;
    wire t44794 = t44793 ^ t44793;
    wire t44795 = t44794 ^ t44794;
    wire t44796 = t44795 ^ t44795;
    wire t44797 = t44796 ^ t44796;
    wire t44798 = t44797 ^ t44797;
    wire t44799 = t44798 ^ t44798;
    wire t44800 = t44799 ^ t44799;
    wire t44801 = t44800 ^ t44800;
    wire t44802 = t44801 ^ t44801;
    wire t44803 = t44802 ^ t44802;
    wire t44804 = t44803 ^ t44803;
    wire t44805 = t44804 ^ t44804;
    wire t44806 = t44805 ^ t44805;
    wire t44807 = t44806 ^ t44806;
    wire t44808 = t44807 ^ t44807;
    wire t44809 = t44808 ^ t44808;
    wire t44810 = t44809 ^ t44809;
    wire t44811 = t44810 ^ t44810;
    wire t44812 = t44811 ^ t44811;
    wire t44813 = t44812 ^ t44812;
    wire t44814 = t44813 ^ t44813;
    wire t44815 = t44814 ^ t44814;
    wire t44816 = t44815 ^ t44815;
    wire t44817 = t44816 ^ t44816;
    wire t44818 = t44817 ^ t44817;
    wire t44819 = t44818 ^ t44818;
    wire t44820 = t44819 ^ t44819;
    wire t44821 = t44820 ^ t44820;
    wire t44822 = t44821 ^ t44821;
    wire t44823 = t44822 ^ t44822;
    wire t44824 = t44823 ^ t44823;
    wire t44825 = t44824 ^ t44824;
    wire t44826 = t44825 ^ t44825;
    wire t44827 = t44826 ^ t44826;
    wire t44828 = t44827 ^ t44827;
    wire t44829 = t44828 ^ t44828;
    wire t44830 = t44829 ^ t44829;
    wire t44831 = t44830 ^ t44830;
    wire t44832 = t44831 ^ t44831;
    wire t44833 = t44832 ^ t44832;
    wire t44834 = t44833 ^ t44833;
    wire t44835 = t44834 ^ t44834;
    wire t44836 = t44835 ^ t44835;
    wire t44837 = t44836 ^ t44836;
    wire t44838 = t44837 ^ t44837;
    wire t44839 = t44838 ^ t44838;
    wire t44840 = t44839 ^ t44839;
    wire t44841 = t44840 ^ t44840;
    wire t44842 = t44841 ^ t44841;
    wire t44843 = t44842 ^ t44842;
    wire t44844 = t44843 ^ t44843;
    wire t44845 = t44844 ^ t44844;
    wire t44846 = t44845 ^ t44845;
    wire t44847 = t44846 ^ t44846;
    wire t44848 = t44847 ^ t44847;
    wire t44849 = t44848 ^ t44848;
    wire t44850 = t44849 ^ t44849;
    wire t44851 = t44850 ^ t44850;
    wire t44852 = t44851 ^ t44851;
    wire t44853 = t44852 ^ t44852;
    wire t44854 = t44853 ^ t44853;
    wire t44855 = t44854 ^ t44854;
    wire t44856 = t44855 ^ t44855;
    wire t44857 = t44856 ^ t44856;
    wire t44858 = t44857 ^ t44857;
    wire t44859 = t44858 ^ t44858;
    wire t44860 = t44859 ^ t44859;
    wire t44861 = t44860 ^ t44860;
    wire t44862 = t44861 ^ t44861;
    wire t44863 = t44862 ^ t44862;
    wire t44864 = t44863 ^ t44863;
    wire t44865 = t44864 ^ t44864;
    wire t44866 = t44865 ^ t44865;
    wire t44867 = t44866 ^ t44866;
    wire t44868 = t44867 ^ t44867;
    wire t44869 = t44868 ^ t44868;
    wire t44870 = t44869 ^ t44869;
    wire t44871 = t44870 ^ t44870;
    wire t44872 = t44871 ^ t44871;
    wire t44873 = t44872 ^ t44872;
    wire t44874 = t44873 ^ t44873;
    wire t44875 = t44874 ^ t44874;
    wire t44876 = t44875 ^ t44875;
    wire t44877 = t44876 ^ t44876;
    wire t44878 = t44877 ^ t44877;
    wire t44879 = t44878 ^ t44878;
    wire t44880 = t44879 ^ t44879;
    wire t44881 = t44880 ^ t44880;
    wire t44882 = t44881 ^ t44881;
    wire t44883 = t44882 ^ t44882;
    wire t44884 = t44883 ^ t44883;
    wire t44885 = t44884 ^ t44884;
    wire t44886 = t44885 ^ t44885;
    wire t44887 = t44886 ^ t44886;
    wire t44888 = t44887 ^ t44887;
    wire t44889 = t44888 ^ t44888;
    wire t44890 = t44889 ^ t44889;
    wire t44891 = t44890 ^ t44890;
    wire t44892 = t44891 ^ t44891;
    wire t44893 = t44892 ^ t44892;
    wire t44894 = t44893 ^ t44893;
    wire t44895 = t44894 ^ t44894;
    wire t44896 = t44895 ^ t44895;
    wire t44897 = t44896 ^ t44896;
    wire t44898 = t44897 ^ t44897;
    wire t44899 = t44898 ^ t44898;
    wire t44900 = t44899 ^ t44899;
    wire t44901 = t44900 ^ t44900;
    wire t44902 = t44901 ^ t44901;
    wire t44903 = t44902 ^ t44902;
    wire t44904 = t44903 ^ t44903;
    wire t44905 = t44904 ^ t44904;
    wire t44906 = t44905 ^ t44905;
    wire t44907 = t44906 ^ t44906;
    wire t44908 = t44907 ^ t44907;
    wire t44909 = t44908 ^ t44908;
    wire t44910 = t44909 ^ t44909;
    wire t44911 = t44910 ^ t44910;
    wire t44912 = t44911 ^ t44911;
    wire t44913 = t44912 ^ t44912;
    wire t44914 = t44913 ^ t44913;
    wire t44915 = t44914 ^ t44914;
    wire t44916 = t44915 ^ t44915;
    wire t44917 = t44916 ^ t44916;
    wire t44918 = t44917 ^ t44917;
    wire t44919 = t44918 ^ t44918;
    wire t44920 = t44919 ^ t44919;
    wire t44921 = t44920 ^ t44920;
    wire t44922 = t44921 ^ t44921;
    wire t44923 = t44922 ^ t44922;
    wire t44924 = t44923 ^ t44923;
    wire t44925 = t44924 ^ t44924;
    wire t44926 = t44925 ^ t44925;
    wire t44927 = t44926 ^ t44926;
    wire t44928 = t44927 ^ t44927;
    wire t44929 = t44928 ^ t44928;
    wire t44930 = t44929 ^ t44929;
    wire t44931 = t44930 ^ t44930;
    wire t44932 = t44931 ^ t44931;
    wire t44933 = t44932 ^ t44932;
    wire t44934 = t44933 ^ t44933;
    wire t44935 = t44934 ^ t44934;
    wire t44936 = t44935 ^ t44935;
    wire t44937 = t44936 ^ t44936;
    wire t44938 = t44937 ^ t44937;
    wire t44939 = t44938 ^ t44938;
    wire t44940 = t44939 ^ t44939;
    wire t44941 = t44940 ^ t44940;
    wire t44942 = t44941 ^ t44941;
    wire t44943 = t44942 ^ t44942;
    wire t44944 = t44943 ^ t44943;
    wire t44945 = t44944 ^ t44944;
    wire t44946 = t44945 ^ t44945;
    wire t44947 = t44946 ^ t44946;
    wire t44948 = t44947 ^ t44947;
    wire t44949 = t44948 ^ t44948;
    wire t44950 = t44949 ^ t44949;
    wire t44951 = t44950 ^ t44950;
    wire t44952 = t44951 ^ t44951;
    wire t44953 = t44952 ^ t44952;
    wire t44954 = t44953 ^ t44953;
    wire t44955 = t44954 ^ t44954;
    wire t44956 = t44955 ^ t44955;
    wire t44957 = t44956 ^ t44956;
    wire t44958 = t44957 ^ t44957;
    wire t44959 = t44958 ^ t44958;
    wire t44960 = t44959 ^ t44959;
    wire t44961 = t44960 ^ t44960;
    wire t44962 = t44961 ^ t44961;
    wire t44963 = t44962 ^ t44962;
    wire t44964 = t44963 ^ t44963;
    wire t44965 = t44964 ^ t44964;
    wire t44966 = t44965 ^ t44965;
    wire t44967 = t44966 ^ t44966;
    wire t44968 = t44967 ^ t44967;
    wire t44969 = t44968 ^ t44968;
    wire t44970 = t44969 ^ t44969;
    wire t44971 = t44970 ^ t44970;
    wire t44972 = t44971 ^ t44971;
    wire t44973 = t44972 ^ t44972;
    wire t44974 = t44973 ^ t44973;
    wire t44975 = t44974 ^ t44974;
    wire t44976 = t44975 ^ t44975;
    wire t44977 = t44976 ^ t44976;
    wire t44978 = t44977 ^ t44977;
    wire t44979 = t44978 ^ t44978;
    wire t44980 = t44979 ^ t44979;
    wire t44981 = t44980 ^ t44980;
    wire t44982 = t44981 ^ t44981;
    wire t44983 = t44982 ^ t44982;
    wire t44984 = t44983 ^ t44983;
    wire t44985 = t44984 ^ t44984;
    wire t44986 = t44985 ^ t44985;
    wire t44987 = t44986 ^ t44986;
    wire t44988 = t44987 ^ t44987;
    wire t44989 = t44988 ^ t44988;
    wire t44990 = t44989 ^ t44989;
    wire t44991 = t44990 ^ t44990;
    wire t44992 = t44991 ^ t44991;
    wire t44993 = t44992 ^ t44992;
    wire t44994 = t44993 ^ t44993;
    wire t44995 = t44994 ^ t44994;
    wire t44996 = t44995 ^ t44995;
    wire t44997 = t44996 ^ t44996;
    wire t44998 = t44997 ^ t44997;
    wire t44999 = t44998 ^ t44998;
    wire t45000 = t44999 ^ t44999;
    wire t45001 = t45000 ^ t45000;
    wire t45002 = t45001 ^ t45001;
    wire t45003 = t45002 ^ t45002;
    wire t45004 = t45003 ^ t45003;
    wire t45005 = t45004 ^ t45004;
    wire t45006 = t45005 ^ t45005;
    wire t45007 = t45006 ^ t45006;
    wire t45008 = t45007 ^ t45007;
    wire t45009 = t45008 ^ t45008;
    wire t45010 = t45009 ^ t45009;
    wire t45011 = t45010 ^ t45010;
    wire t45012 = t45011 ^ t45011;
    wire t45013 = t45012 ^ t45012;
    wire t45014 = t45013 ^ t45013;
    wire t45015 = t45014 ^ t45014;
    wire t45016 = t45015 ^ t45015;
    wire t45017 = t45016 ^ t45016;
    wire t45018 = t45017 ^ t45017;
    wire t45019 = t45018 ^ t45018;
    wire t45020 = t45019 ^ t45019;
    wire t45021 = t45020 ^ t45020;
    wire t45022 = t45021 ^ t45021;
    wire t45023 = t45022 ^ t45022;
    wire t45024 = t45023 ^ t45023;
    wire t45025 = t45024 ^ t45024;
    wire t45026 = t45025 ^ t45025;
    wire t45027 = t45026 ^ t45026;
    wire t45028 = t45027 ^ t45027;
    wire t45029 = t45028 ^ t45028;
    wire t45030 = t45029 ^ t45029;
    wire t45031 = t45030 ^ t45030;
    wire t45032 = t45031 ^ t45031;
    wire t45033 = t45032 ^ t45032;
    wire t45034 = t45033 ^ t45033;
    wire t45035 = t45034 ^ t45034;
    wire t45036 = t45035 ^ t45035;
    wire t45037 = t45036 ^ t45036;
    wire t45038 = t45037 ^ t45037;
    wire t45039 = t45038 ^ t45038;
    wire t45040 = t45039 ^ t45039;
    wire t45041 = t45040 ^ t45040;
    wire t45042 = t45041 ^ t45041;
    wire t45043 = t45042 ^ t45042;
    wire t45044 = t45043 ^ t45043;
    wire t45045 = t45044 ^ t45044;
    wire t45046 = t45045 ^ t45045;
    wire t45047 = t45046 ^ t45046;
    wire t45048 = t45047 ^ t45047;
    wire t45049 = t45048 ^ t45048;
    wire t45050 = t45049 ^ t45049;
    wire t45051 = t45050 ^ t45050;
    wire t45052 = t45051 ^ t45051;
    wire t45053 = t45052 ^ t45052;
    wire t45054 = t45053 ^ t45053;
    wire t45055 = t45054 ^ t45054;
    wire t45056 = t45055 ^ t45055;
    wire t45057 = t45056 ^ t45056;
    wire t45058 = t45057 ^ t45057;
    wire t45059 = t45058 ^ t45058;
    wire t45060 = t45059 ^ t45059;
    wire t45061 = t45060 ^ t45060;
    wire t45062 = t45061 ^ t45061;
    wire t45063 = t45062 ^ t45062;
    wire t45064 = t45063 ^ t45063;
    wire t45065 = t45064 ^ t45064;
    wire t45066 = t45065 ^ t45065;
    wire t45067 = t45066 ^ t45066;
    wire t45068 = t45067 ^ t45067;
    wire t45069 = t45068 ^ t45068;
    wire t45070 = t45069 ^ t45069;
    wire t45071 = t45070 ^ t45070;
    wire t45072 = t45071 ^ t45071;
    wire t45073 = t45072 ^ t45072;
    wire t45074 = t45073 ^ t45073;
    wire t45075 = t45074 ^ t45074;
    wire t45076 = t45075 ^ t45075;
    wire t45077 = t45076 ^ t45076;
    wire t45078 = t45077 ^ t45077;
    wire t45079 = t45078 ^ t45078;
    wire t45080 = t45079 ^ t45079;
    wire t45081 = t45080 ^ t45080;
    wire t45082 = t45081 ^ t45081;
    wire t45083 = t45082 ^ t45082;
    wire t45084 = t45083 ^ t45083;
    wire t45085 = t45084 ^ t45084;
    wire t45086 = t45085 ^ t45085;
    wire t45087 = t45086 ^ t45086;
    wire t45088 = t45087 ^ t45087;
    wire t45089 = t45088 ^ t45088;
    wire t45090 = t45089 ^ t45089;
    wire t45091 = t45090 ^ t45090;
    wire t45092 = t45091 ^ t45091;
    wire t45093 = t45092 ^ t45092;
    wire t45094 = t45093 ^ t45093;
    wire t45095 = t45094 ^ t45094;
    wire t45096 = t45095 ^ t45095;
    wire t45097 = t45096 ^ t45096;
    wire t45098 = t45097 ^ t45097;
    wire t45099 = t45098 ^ t45098;
    wire t45100 = t45099 ^ t45099;
    wire t45101 = t45100 ^ t45100;
    wire t45102 = t45101 ^ t45101;
    wire t45103 = t45102 ^ t45102;
    wire t45104 = t45103 ^ t45103;
    wire t45105 = t45104 ^ t45104;
    wire t45106 = t45105 ^ t45105;
    wire t45107 = t45106 ^ t45106;
    wire t45108 = t45107 ^ t45107;
    wire t45109 = t45108 ^ t45108;
    wire t45110 = t45109 ^ t45109;
    wire t45111 = t45110 ^ t45110;
    wire t45112 = t45111 ^ t45111;
    wire t45113 = t45112 ^ t45112;
    wire t45114 = t45113 ^ t45113;
    wire t45115 = t45114 ^ t45114;
    wire t45116 = t45115 ^ t45115;
    wire t45117 = t45116 ^ t45116;
    wire t45118 = t45117 ^ t45117;
    wire t45119 = t45118 ^ t45118;
    wire t45120 = t45119 ^ t45119;
    wire t45121 = t45120 ^ t45120;
    wire t45122 = t45121 ^ t45121;
    wire t45123 = t45122 ^ t45122;
    wire t45124 = t45123 ^ t45123;
    wire t45125 = t45124 ^ t45124;
    wire t45126 = t45125 ^ t45125;
    wire t45127 = t45126 ^ t45126;
    wire t45128 = t45127 ^ t45127;
    wire t45129 = t45128 ^ t45128;
    wire t45130 = t45129 ^ t45129;
    wire t45131 = t45130 ^ t45130;
    wire t45132 = t45131 ^ t45131;
    wire t45133 = t45132 ^ t45132;
    wire t45134 = t45133 ^ t45133;
    wire t45135 = t45134 ^ t45134;
    wire t45136 = t45135 ^ t45135;
    wire t45137 = t45136 ^ t45136;
    wire t45138 = t45137 ^ t45137;
    wire t45139 = t45138 ^ t45138;
    wire t45140 = t45139 ^ t45139;
    wire t45141 = t45140 ^ t45140;
    wire t45142 = t45141 ^ t45141;
    wire t45143 = t45142 ^ t45142;
    wire t45144 = t45143 ^ t45143;
    wire t45145 = t45144 ^ t45144;
    wire t45146 = t45145 ^ t45145;
    wire t45147 = t45146 ^ t45146;
    wire t45148 = t45147 ^ t45147;
    wire t45149 = t45148 ^ t45148;
    wire t45150 = t45149 ^ t45149;
    wire t45151 = t45150 ^ t45150;
    wire t45152 = t45151 ^ t45151;
    wire t45153 = t45152 ^ t45152;
    wire t45154 = t45153 ^ t45153;
    wire t45155 = t45154 ^ t45154;
    wire t45156 = t45155 ^ t45155;
    wire t45157 = t45156 ^ t45156;
    wire t45158 = t45157 ^ t45157;
    wire t45159 = t45158 ^ t45158;
    wire t45160 = t45159 ^ t45159;
    wire t45161 = t45160 ^ t45160;
    wire t45162 = t45161 ^ t45161;
    wire t45163 = t45162 ^ t45162;
    wire t45164 = t45163 ^ t45163;
    wire t45165 = t45164 ^ t45164;
    wire t45166 = t45165 ^ t45165;
    wire t45167 = t45166 ^ t45166;
    wire t45168 = t45167 ^ t45167;
    wire t45169 = t45168 ^ t45168;
    wire t45170 = t45169 ^ t45169;
    wire t45171 = t45170 ^ t45170;
    wire t45172 = t45171 ^ t45171;
    wire t45173 = t45172 ^ t45172;
    wire t45174 = t45173 ^ t45173;
    wire t45175 = t45174 ^ t45174;
    wire t45176 = t45175 ^ t45175;
    wire t45177 = t45176 ^ t45176;
    wire t45178 = t45177 ^ t45177;
    wire t45179 = t45178 ^ t45178;
    wire t45180 = t45179 ^ t45179;
    wire t45181 = t45180 ^ t45180;
    wire t45182 = t45181 ^ t45181;
    wire t45183 = t45182 ^ t45182;
    wire t45184 = t45183 ^ t45183;
    wire t45185 = t45184 ^ t45184;
    wire t45186 = t45185 ^ t45185;
    wire t45187 = t45186 ^ t45186;
    wire t45188 = t45187 ^ t45187;
    wire t45189 = t45188 ^ t45188;
    wire t45190 = t45189 ^ t45189;
    wire t45191 = t45190 ^ t45190;
    wire t45192 = t45191 ^ t45191;
    wire t45193 = t45192 ^ t45192;
    wire t45194 = t45193 ^ t45193;
    wire t45195 = t45194 ^ t45194;
    wire t45196 = t45195 ^ t45195;
    wire t45197 = t45196 ^ t45196;
    wire t45198 = t45197 ^ t45197;
    wire t45199 = t45198 ^ t45198;
    wire t45200 = t45199 ^ t45199;
    wire t45201 = t45200 ^ t45200;
    wire t45202 = t45201 ^ t45201;
    wire t45203 = t45202 ^ t45202;
    wire t45204 = t45203 ^ t45203;
    wire t45205 = t45204 ^ t45204;
    wire t45206 = t45205 ^ t45205;
    wire t45207 = t45206 ^ t45206;
    wire t45208 = t45207 ^ t45207;
    wire t45209 = t45208 ^ t45208;
    wire t45210 = t45209 ^ t45209;
    wire t45211 = t45210 ^ t45210;
    wire t45212 = t45211 ^ t45211;
    wire t45213 = t45212 ^ t45212;
    wire t45214 = t45213 ^ t45213;
    wire t45215 = t45214 ^ t45214;
    wire t45216 = t45215 ^ t45215;
    wire t45217 = t45216 ^ t45216;
    wire t45218 = t45217 ^ t45217;
    wire t45219 = t45218 ^ t45218;
    wire t45220 = t45219 ^ t45219;
    wire t45221 = t45220 ^ t45220;
    wire t45222 = t45221 ^ t45221;
    wire t45223 = t45222 ^ t45222;
    wire t45224 = t45223 ^ t45223;
    wire t45225 = t45224 ^ t45224;
    wire t45226 = t45225 ^ t45225;
    wire t45227 = t45226 ^ t45226;
    wire t45228 = t45227 ^ t45227;
    wire t45229 = t45228 ^ t45228;
    wire t45230 = t45229 ^ t45229;
    wire t45231 = t45230 ^ t45230;
    wire t45232 = t45231 ^ t45231;
    wire t45233 = t45232 ^ t45232;
    wire t45234 = t45233 ^ t45233;
    wire t45235 = t45234 ^ t45234;
    wire t45236 = t45235 ^ t45235;
    wire t45237 = t45236 ^ t45236;
    wire t45238 = t45237 ^ t45237;
    wire t45239 = t45238 ^ t45238;
    wire t45240 = t45239 ^ t45239;
    wire t45241 = t45240 ^ t45240;
    wire t45242 = t45241 ^ t45241;
    wire t45243 = t45242 ^ t45242;
    wire t45244 = t45243 ^ t45243;
    wire t45245 = t45244 ^ t45244;
    wire t45246 = t45245 ^ t45245;
    wire t45247 = t45246 ^ t45246;
    wire t45248 = t45247 ^ t45247;
    wire t45249 = t45248 ^ t45248;
    wire t45250 = t45249 ^ t45249;
    wire t45251 = t45250 ^ t45250;
    wire t45252 = t45251 ^ t45251;
    wire t45253 = t45252 ^ t45252;
    wire t45254 = t45253 ^ t45253;
    wire t45255 = t45254 ^ t45254;
    wire t45256 = t45255 ^ t45255;
    wire t45257 = t45256 ^ t45256;
    wire t45258 = t45257 ^ t45257;
    wire t45259 = t45258 ^ t45258;
    wire t45260 = t45259 ^ t45259;
    wire t45261 = t45260 ^ t45260;
    wire t45262 = t45261 ^ t45261;
    wire t45263 = t45262 ^ t45262;
    wire t45264 = t45263 ^ t45263;
    wire t45265 = t45264 ^ t45264;
    wire t45266 = t45265 ^ t45265;
    wire t45267 = t45266 ^ t45266;
    wire t45268 = t45267 ^ t45267;
    wire t45269 = t45268 ^ t45268;
    wire t45270 = t45269 ^ t45269;
    wire t45271 = t45270 ^ t45270;
    wire t45272 = t45271 ^ t45271;
    wire t45273 = t45272 ^ t45272;
    wire t45274 = t45273 ^ t45273;
    wire t45275 = t45274 ^ t45274;
    wire t45276 = t45275 ^ t45275;
    wire t45277 = t45276 ^ t45276;
    wire t45278 = t45277 ^ t45277;
    wire t45279 = t45278 ^ t45278;
    wire t45280 = t45279 ^ t45279;
    wire t45281 = t45280 ^ t45280;
    wire t45282 = t45281 ^ t45281;
    wire t45283 = t45282 ^ t45282;
    wire t45284 = t45283 ^ t45283;
    wire t45285 = t45284 ^ t45284;
    wire t45286 = t45285 ^ t45285;
    wire t45287 = t45286 ^ t45286;
    wire t45288 = t45287 ^ t45287;
    wire t45289 = t45288 ^ t45288;
    wire t45290 = t45289 ^ t45289;
    wire t45291 = t45290 ^ t45290;
    wire t45292 = t45291 ^ t45291;
    wire t45293 = t45292 ^ t45292;
    wire t45294 = t45293 ^ t45293;
    wire t45295 = t45294 ^ t45294;
    wire t45296 = t45295 ^ t45295;
    wire t45297 = t45296 ^ t45296;
    wire t45298 = t45297 ^ t45297;
    wire t45299 = t45298 ^ t45298;
    wire t45300 = t45299 ^ t45299;
    wire t45301 = t45300 ^ t45300;
    wire t45302 = t45301 ^ t45301;
    wire t45303 = t45302 ^ t45302;
    wire t45304 = t45303 ^ t45303;
    wire t45305 = t45304 ^ t45304;
    wire t45306 = t45305 ^ t45305;
    wire t45307 = t45306 ^ t45306;
    wire t45308 = t45307 ^ t45307;
    wire t45309 = t45308 ^ t45308;
    wire t45310 = t45309 ^ t45309;
    wire t45311 = t45310 ^ t45310;
    wire t45312 = t45311 ^ t45311;
    wire t45313 = t45312 ^ t45312;
    wire t45314 = t45313 ^ t45313;
    wire t45315 = t45314 ^ t45314;
    wire t45316 = t45315 ^ t45315;
    wire t45317 = t45316 ^ t45316;
    wire t45318 = t45317 ^ t45317;
    wire t45319 = t45318 ^ t45318;
    wire t45320 = t45319 ^ t45319;
    wire t45321 = t45320 ^ t45320;
    wire t45322 = t45321 ^ t45321;
    wire t45323 = t45322 ^ t45322;
    wire t45324 = t45323 ^ t45323;
    wire t45325 = t45324 ^ t45324;
    wire t45326 = t45325 ^ t45325;
    wire t45327 = t45326 ^ t45326;
    wire t45328 = t45327 ^ t45327;
    wire t45329 = t45328 ^ t45328;
    wire t45330 = t45329 ^ t45329;
    wire t45331 = t45330 ^ t45330;
    wire t45332 = t45331 ^ t45331;
    wire t45333 = t45332 ^ t45332;
    wire t45334 = t45333 ^ t45333;
    wire t45335 = t45334 ^ t45334;
    wire t45336 = t45335 ^ t45335;
    wire t45337 = t45336 ^ t45336;
    wire t45338 = t45337 ^ t45337;
    wire t45339 = t45338 ^ t45338;
    wire t45340 = t45339 ^ t45339;
    wire t45341 = t45340 ^ t45340;
    wire t45342 = t45341 ^ t45341;
    wire t45343 = t45342 ^ t45342;
    wire t45344 = t45343 ^ t45343;
    wire t45345 = t45344 ^ t45344;
    wire t45346 = t45345 ^ t45345;
    wire t45347 = t45346 ^ t45346;
    wire t45348 = t45347 ^ t45347;
    wire t45349 = t45348 ^ t45348;
    wire t45350 = t45349 ^ t45349;
    wire t45351 = t45350 ^ t45350;
    wire t45352 = t45351 ^ t45351;
    wire t45353 = t45352 ^ t45352;
    wire t45354 = t45353 ^ t45353;
    wire t45355 = t45354 ^ t45354;
    wire t45356 = t45355 ^ t45355;
    wire t45357 = t45356 ^ t45356;
    wire t45358 = t45357 ^ t45357;
    wire t45359 = t45358 ^ t45358;
    wire t45360 = t45359 ^ t45359;
    wire t45361 = t45360 ^ t45360;
    wire t45362 = t45361 ^ t45361;
    wire t45363 = t45362 ^ t45362;
    wire t45364 = t45363 ^ t45363;
    wire t45365 = t45364 ^ t45364;
    wire t45366 = t45365 ^ t45365;
    wire t45367 = t45366 ^ t45366;
    wire t45368 = t45367 ^ t45367;
    wire t45369 = t45368 ^ t45368;
    wire t45370 = t45369 ^ t45369;
    wire t45371 = t45370 ^ t45370;
    wire t45372 = t45371 ^ t45371;
    wire t45373 = t45372 ^ t45372;
    wire t45374 = t45373 ^ t45373;
    wire t45375 = t45374 ^ t45374;
    wire t45376 = t45375 ^ t45375;
    wire t45377 = t45376 ^ t45376;
    wire t45378 = t45377 ^ t45377;
    wire t45379 = t45378 ^ t45378;
    wire t45380 = t45379 ^ t45379;
    wire t45381 = t45380 ^ t45380;
    wire t45382 = t45381 ^ t45381;
    wire t45383 = t45382 ^ t45382;
    wire t45384 = t45383 ^ t45383;
    wire t45385 = t45384 ^ t45384;
    wire t45386 = t45385 ^ t45385;
    wire t45387 = t45386 ^ t45386;
    wire t45388 = t45387 ^ t45387;
    wire t45389 = t45388 ^ t45388;
    wire t45390 = t45389 ^ t45389;
    wire t45391 = t45390 ^ t45390;
    wire t45392 = t45391 ^ t45391;
    wire t45393 = t45392 ^ t45392;
    wire t45394 = t45393 ^ t45393;
    wire t45395 = t45394 ^ t45394;
    wire t45396 = t45395 ^ t45395;
    wire t45397 = t45396 ^ t45396;
    wire t45398 = t45397 ^ t45397;
    wire t45399 = t45398 ^ t45398;
    wire t45400 = t45399 ^ t45399;
    wire t45401 = t45400 ^ t45400;
    wire t45402 = t45401 ^ t45401;
    wire t45403 = t45402 ^ t45402;
    wire t45404 = t45403 ^ t45403;
    wire t45405 = t45404 ^ t45404;
    wire t45406 = t45405 ^ t45405;
    wire t45407 = t45406 ^ t45406;
    wire t45408 = t45407 ^ t45407;
    wire t45409 = t45408 ^ t45408;
    wire t45410 = t45409 ^ t45409;
    wire t45411 = t45410 ^ t45410;
    wire t45412 = t45411 ^ t45411;
    wire t45413 = t45412 ^ t45412;
    wire t45414 = t45413 ^ t45413;
    wire t45415 = t45414 ^ t45414;
    wire t45416 = t45415 ^ t45415;
    wire t45417 = t45416 ^ t45416;
    wire t45418 = t45417 ^ t45417;
    wire t45419 = t45418 ^ t45418;
    wire t45420 = t45419 ^ t45419;
    wire t45421 = t45420 ^ t45420;
    wire t45422 = t45421 ^ t45421;
    wire t45423 = t45422 ^ t45422;
    wire t45424 = t45423 ^ t45423;
    wire t45425 = t45424 ^ t45424;
    wire t45426 = t45425 ^ t45425;
    wire t45427 = t45426 ^ t45426;
    wire t45428 = t45427 ^ t45427;
    wire t45429 = t45428 ^ t45428;
    wire t45430 = t45429 ^ t45429;
    wire t45431 = t45430 ^ t45430;
    wire t45432 = t45431 ^ t45431;
    wire t45433 = t45432 ^ t45432;
    wire t45434 = t45433 ^ t45433;
    wire t45435 = t45434 ^ t45434;
    wire t45436 = t45435 ^ t45435;
    wire t45437 = t45436 ^ t45436;
    wire t45438 = t45437 ^ t45437;
    wire t45439 = t45438 ^ t45438;
    wire t45440 = t45439 ^ t45439;
    wire t45441 = t45440 ^ t45440;
    wire t45442 = t45441 ^ t45441;
    wire t45443 = t45442 ^ t45442;
    wire t45444 = t45443 ^ t45443;
    wire t45445 = t45444 ^ t45444;
    wire t45446 = t45445 ^ t45445;
    wire t45447 = t45446 ^ t45446;
    wire t45448 = t45447 ^ t45447;
    wire t45449 = t45448 ^ t45448;
    wire t45450 = t45449 ^ t45449;
    wire t45451 = t45450 ^ t45450;
    wire t45452 = t45451 ^ t45451;
    wire t45453 = t45452 ^ t45452;
    wire t45454 = t45453 ^ t45453;
    wire t45455 = t45454 ^ t45454;
    wire t45456 = t45455 ^ t45455;
    wire t45457 = t45456 ^ t45456;
    wire t45458 = t45457 ^ t45457;
    wire t45459 = t45458 ^ t45458;
    wire t45460 = t45459 ^ t45459;
    wire t45461 = t45460 ^ t45460;
    wire t45462 = t45461 ^ t45461;
    wire t45463 = t45462 ^ t45462;
    wire t45464 = t45463 ^ t45463;
    wire t45465 = t45464 ^ t45464;
    wire t45466 = t45465 ^ t45465;
    wire t45467 = t45466 ^ t45466;
    wire t45468 = t45467 ^ t45467;
    wire t45469 = t45468 ^ t45468;
    wire t45470 = t45469 ^ t45469;
    wire t45471 = t45470 ^ t45470;
    wire t45472 = t45471 ^ t45471;
    wire t45473 = t45472 ^ t45472;
    wire t45474 = t45473 ^ t45473;
    wire t45475 = t45474 ^ t45474;
    wire t45476 = t45475 ^ t45475;
    wire t45477 = t45476 ^ t45476;
    wire t45478 = t45477 ^ t45477;
    wire t45479 = t45478 ^ t45478;
    wire t45480 = t45479 ^ t45479;
    wire t45481 = t45480 ^ t45480;
    wire t45482 = t45481 ^ t45481;
    wire t45483 = t45482 ^ t45482;
    wire t45484 = t45483 ^ t45483;
    wire t45485 = t45484 ^ t45484;
    wire t45486 = t45485 ^ t45485;
    wire t45487 = t45486 ^ t45486;
    wire t45488 = t45487 ^ t45487;
    wire t45489 = t45488 ^ t45488;
    wire t45490 = t45489 ^ t45489;
    wire t45491 = t45490 ^ t45490;
    wire t45492 = t45491 ^ t45491;
    wire t45493 = t45492 ^ t45492;
    wire t45494 = t45493 ^ t45493;
    wire t45495 = t45494 ^ t45494;
    wire t45496 = t45495 ^ t45495;
    wire t45497 = t45496 ^ t45496;
    wire t45498 = t45497 ^ t45497;
    wire t45499 = t45498 ^ t45498;
    wire t45500 = t45499 ^ t45499;
    wire t45501 = t45500 ^ t45500;
    wire t45502 = t45501 ^ t45501;
    wire t45503 = t45502 ^ t45502;
    wire t45504 = t45503 ^ t45503;
    wire t45505 = t45504 ^ t45504;
    wire t45506 = t45505 ^ t45505;
    wire t45507 = t45506 ^ t45506;
    wire t45508 = t45507 ^ t45507;
    wire t45509 = t45508 ^ t45508;
    wire t45510 = t45509 ^ t45509;
    wire t45511 = t45510 ^ t45510;
    wire t45512 = t45511 ^ t45511;
    wire t45513 = t45512 ^ t45512;
    wire t45514 = t45513 ^ t45513;
    wire t45515 = t45514 ^ t45514;
    wire t45516 = t45515 ^ t45515;
    wire t45517 = t45516 ^ t45516;
    wire t45518 = t45517 ^ t45517;
    wire t45519 = t45518 ^ t45518;
    wire t45520 = t45519 ^ t45519;
    wire t45521 = t45520 ^ t45520;
    wire t45522 = t45521 ^ t45521;
    wire t45523 = t45522 ^ t45522;
    wire t45524 = t45523 ^ t45523;
    wire t45525 = t45524 ^ t45524;
    wire t45526 = t45525 ^ t45525;
    wire t45527 = t45526 ^ t45526;
    wire t45528 = t45527 ^ t45527;
    wire t45529 = t45528 ^ t45528;
    wire t45530 = t45529 ^ t45529;
    wire t45531 = t45530 ^ t45530;
    wire t45532 = t45531 ^ t45531;
    wire t45533 = t45532 ^ t45532;
    wire t45534 = t45533 ^ t45533;
    wire t45535 = t45534 ^ t45534;
    wire t45536 = t45535 ^ t45535;
    wire t45537 = t45536 ^ t45536;
    wire t45538 = t45537 ^ t45537;
    wire t45539 = t45538 ^ t45538;
    wire t45540 = t45539 ^ t45539;
    wire t45541 = t45540 ^ t45540;
    wire t45542 = t45541 ^ t45541;
    wire t45543 = t45542 ^ t45542;
    wire t45544 = t45543 ^ t45543;
    wire t45545 = t45544 ^ t45544;
    wire t45546 = t45545 ^ t45545;
    wire t45547 = t45546 ^ t45546;
    wire t45548 = t45547 ^ t45547;
    wire t45549 = t45548 ^ t45548;
    wire t45550 = t45549 ^ t45549;
    wire t45551 = t45550 ^ t45550;
    wire t45552 = t45551 ^ t45551;
    wire t45553 = t45552 ^ t45552;
    wire t45554 = t45553 ^ t45553;
    wire t45555 = t45554 ^ t45554;
    wire t45556 = t45555 ^ t45555;
    wire t45557 = t45556 ^ t45556;
    wire t45558 = t45557 ^ t45557;
    wire t45559 = t45558 ^ t45558;
    wire t45560 = t45559 ^ t45559;
    wire t45561 = t45560 ^ t45560;
    wire t45562 = t45561 ^ t45561;
    wire t45563 = t45562 ^ t45562;
    wire t45564 = t45563 ^ t45563;
    wire t45565 = t45564 ^ t45564;
    wire t45566 = t45565 ^ t45565;
    wire t45567 = t45566 ^ t45566;
    wire t45568 = t45567 ^ t45567;
    wire t45569 = t45568 ^ t45568;
    wire t45570 = t45569 ^ t45569;
    wire t45571 = t45570 ^ t45570;
    wire t45572 = t45571 ^ t45571;
    wire t45573 = t45572 ^ t45572;
    wire t45574 = t45573 ^ t45573;
    wire t45575 = t45574 ^ t45574;
    wire t45576 = t45575 ^ t45575;
    wire t45577 = t45576 ^ t45576;
    wire t45578 = t45577 ^ t45577;
    wire t45579 = t45578 ^ t45578;
    wire t45580 = t45579 ^ t45579;
    wire t45581 = t45580 ^ t45580;
    wire t45582 = t45581 ^ t45581;
    wire t45583 = t45582 ^ t45582;
    wire t45584 = t45583 ^ t45583;
    wire t45585 = t45584 ^ t45584;
    wire t45586 = t45585 ^ t45585;
    wire t45587 = t45586 ^ t45586;
    wire t45588 = t45587 ^ t45587;
    wire t45589 = t45588 ^ t45588;
    wire t45590 = t45589 ^ t45589;
    wire t45591 = t45590 ^ t45590;
    wire t45592 = t45591 ^ t45591;
    wire t45593 = t45592 ^ t45592;
    wire t45594 = t45593 ^ t45593;
    wire t45595 = t45594 ^ t45594;
    wire t45596 = t45595 ^ t45595;
    wire t45597 = t45596 ^ t45596;
    wire t45598 = t45597 ^ t45597;
    wire t45599 = t45598 ^ t45598;
    wire t45600 = t45599 ^ t45599;
    wire t45601 = t45600 ^ t45600;
    wire t45602 = t45601 ^ t45601;
    wire t45603 = t45602 ^ t45602;
    wire t45604 = t45603 ^ t45603;
    wire t45605 = t45604 ^ t45604;
    wire t45606 = t45605 ^ t45605;
    wire t45607 = t45606 ^ t45606;
    wire t45608 = t45607 ^ t45607;
    wire t45609 = t45608 ^ t45608;
    wire t45610 = t45609 ^ t45609;
    wire t45611 = t45610 ^ t45610;
    wire t45612 = t45611 ^ t45611;
    wire t45613 = t45612 ^ t45612;
    wire t45614 = t45613 ^ t45613;
    wire t45615 = t45614 ^ t45614;
    wire t45616 = t45615 ^ t45615;
    wire t45617 = t45616 ^ t45616;
    wire t45618 = t45617 ^ t45617;
    wire t45619 = t45618 ^ t45618;
    wire t45620 = t45619 ^ t45619;
    wire t45621 = t45620 ^ t45620;
    wire t45622 = t45621 ^ t45621;
    wire t45623 = t45622 ^ t45622;
    wire t45624 = t45623 ^ t45623;
    wire t45625 = t45624 ^ t45624;
    wire t45626 = t45625 ^ t45625;
    wire t45627 = t45626 ^ t45626;
    wire t45628 = t45627 ^ t45627;
    wire t45629 = t45628 ^ t45628;
    wire t45630 = t45629 ^ t45629;
    wire t45631 = t45630 ^ t45630;
    wire t45632 = t45631 ^ t45631;
    wire t45633 = t45632 ^ t45632;
    wire t45634 = t45633 ^ t45633;
    wire t45635 = t45634 ^ t45634;
    wire t45636 = t45635 ^ t45635;
    wire t45637 = t45636 ^ t45636;
    wire t45638 = t45637 ^ t45637;
    wire t45639 = t45638 ^ t45638;
    wire t45640 = t45639 ^ t45639;
    wire t45641 = t45640 ^ t45640;
    wire t45642 = t45641 ^ t45641;
    wire t45643 = t45642 ^ t45642;
    wire t45644 = t45643 ^ t45643;
    wire t45645 = t45644 ^ t45644;
    wire t45646 = t45645 ^ t45645;
    wire t45647 = t45646 ^ t45646;
    wire t45648 = t45647 ^ t45647;
    wire t45649 = t45648 ^ t45648;
    wire t45650 = t45649 ^ t45649;
    wire t45651 = t45650 ^ t45650;
    wire t45652 = t45651 ^ t45651;
    wire t45653 = t45652 ^ t45652;
    wire t45654 = t45653 ^ t45653;
    wire t45655 = t45654 ^ t45654;
    wire t45656 = t45655 ^ t45655;
    wire t45657 = t45656 ^ t45656;
    wire t45658 = t45657 ^ t45657;
    wire t45659 = t45658 ^ t45658;
    wire t45660 = t45659 ^ t45659;
    wire t45661 = t45660 ^ t45660;
    wire t45662 = t45661 ^ t45661;
    wire t45663 = t45662 ^ t45662;
    wire t45664 = t45663 ^ t45663;
    wire t45665 = t45664 ^ t45664;
    wire t45666 = t45665 ^ t45665;
    wire t45667 = t45666 ^ t45666;
    wire t45668 = t45667 ^ t45667;
    wire t45669 = t45668 ^ t45668;
    wire t45670 = t45669 ^ t45669;
    wire t45671 = t45670 ^ t45670;
    wire t45672 = t45671 ^ t45671;
    wire t45673 = t45672 ^ t45672;
    wire t45674 = t45673 ^ t45673;
    wire t45675 = t45674 ^ t45674;
    wire t45676 = t45675 ^ t45675;
    wire t45677 = t45676 ^ t45676;
    wire t45678 = t45677 ^ t45677;
    wire t45679 = t45678 ^ t45678;
    wire t45680 = t45679 ^ t45679;
    wire t45681 = t45680 ^ t45680;
    wire t45682 = t45681 ^ t45681;
    wire t45683 = t45682 ^ t45682;
    wire t45684 = t45683 ^ t45683;
    wire t45685 = t45684 ^ t45684;
    wire t45686 = t45685 ^ t45685;
    wire t45687 = t45686 ^ t45686;
    wire t45688 = t45687 ^ t45687;
    wire t45689 = t45688 ^ t45688;
    wire t45690 = t45689 ^ t45689;
    wire t45691 = t45690 ^ t45690;
    wire t45692 = t45691 ^ t45691;
    wire t45693 = t45692 ^ t45692;
    wire t45694 = t45693 ^ t45693;
    wire t45695 = t45694 ^ t45694;
    wire t45696 = t45695 ^ t45695;
    wire t45697 = t45696 ^ t45696;
    wire t45698 = t45697 ^ t45697;
    wire t45699 = t45698 ^ t45698;
    wire t45700 = t45699 ^ t45699;
    wire t45701 = t45700 ^ t45700;
    wire t45702 = t45701 ^ t45701;
    wire t45703 = t45702 ^ t45702;
    wire t45704 = t45703 ^ t45703;
    wire t45705 = t45704 ^ t45704;
    wire t45706 = t45705 ^ t45705;
    wire t45707 = t45706 ^ t45706;
    wire t45708 = t45707 ^ t45707;
    wire t45709 = t45708 ^ t45708;
    wire t45710 = t45709 ^ t45709;
    wire t45711 = t45710 ^ t45710;
    wire t45712 = t45711 ^ t45711;
    wire t45713 = t45712 ^ t45712;
    wire t45714 = t45713 ^ t45713;
    wire t45715 = t45714 ^ t45714;
    wire t45716 = t45715 ^ t45715;
    wire t45717 = t45716 ^ t45716;
    wire t45718 = t45717 ^ t45717;
    wire t45719 = t45718 ^ t45718;
    wire t45720 = t45719 ^ t45719;
    wire t45721 = t45720 ^ t45720;
    wire t45722 = t45721 ^ t45721;
    wire t45723 = t45722 ^ t45722;
    wire t45724 = t45723 ^ t45723;
    wire t45725 = t45724 ^ t45724;
    wire t45726 = t45725 ^ t45725;
    wire t45727 = t45726 ^ t45726;
    wire t45728 = t45727 ^ t45727;
    wire t45729 = t45728 ^ t45728;
    wire t45730 = t45729 ^ t45729;
    wire t45731 = t45730 ^ t45730;
    wire t45732 = t45731 ^ t45731;
    wire t45733 = t45732 ^ t45732;
    wire t45734 = t45733 ^ t45733;
    wire t45735 = t45734 ^ t45734;
    wire t45736 = t45735 ^ t45735;
    wire t45737 = t45736 ^ t45736;
    wire t45738 = t45737 ^ t45737;
    wire t45739 = t45738 ^ t45738;
    wire t45740 = t45739 ^ t45739;
    wire t45741 = t45740 ^ t45740;
    wire t45742 = t45741 ^ t45741;
    wire t45743 = t45742 ^ t45742;
    wire t45744 = t45743 ^ t45743;
    wire t45745 = t45744 ^ t45744;
    wire t45746 = t45745 ^ t45745;
    wire t45747 = t45746 ^ t45746;
    wire t45748 = t45747 ^ t45747;
    wire t45749 = t45748 ^ t45748;
    wire t45750 = t45749 ^ t45749;
    wire t45751 = t45750 ^ t45750;
    wire t45752 = t45751 ^ t45751;
    wire t45753 = t45752 ^ t45752;
    wire t45754 = t45753 ^ t45753;
    wire t45755 = t45754 ^ t45754;
    wire t45756 = t45755 ^ t45755;
    wire t45757 = t45756 ^ t45756;
    wire t45758 = t45757 ^ t45757;
    wire t45759 = t45758 ^ t45758;
    wire t45760 = t45759 ^ t45759;
    wire t45761 = t45760 ^ t45760;
    wire t45762 = t45761 ^ t45761;
    wire t45763 = t45762 ^ t45762;
    wire t45764 = t45763 ^ t45763;
    wire t45765 = t45764 ^ t45764;
    wire t45766 = t45765 ^ t45765;
    wire t45767 = t45766 ^ t45766;
    wire t45768 = t45767 ^ t45767;
    wire t45769 = t45768 ^ t45768;
    wire t45770 = t45769 ^ t45769;
    wire t45771 = t45770 ^ t45770;
    wire t45772 = t45771 ^ t45771;
    wire t45773 = t45772 ^ t45772;
    wire t45774 = t45773 ^ t45773;
    wire t45775 = t45774 ^ t45774;
    wire t45776 = t45775 ^ t45775;
    wire t45777 = t45776 ^ t45776;
    wire t45778 = t45777 ^ t45777;
    wire t45779 = t45778 ^ t45778;
    wire t45780 = t45779 ^ t45779;
    wire t45781 = t45780 ^ t45780;
    wire t45782 = t45781 ^ t45781;
    wire t45783 = t45782 ^ t45782;
    wire t45784 = t45783 ^ t45783;
    wire t45785 = t45784 ^ t45784;
    wire t45786 = t45785 ^ t45785;
    wire t45787 = t45786 ^ t45786;
    wire t45788 = t45787 ^ t45787;
    wire t45789 = t45788 ^ t45788;
    wire t45790 = t45789 ^ t45789;
    wire t45791 = t45790 ^ t45790;
    wire t45792 = t45791 ^ t45791;
    wire t45793 = t45792 ^ t45792;
    wire t45794 = t45793 ^ t45793;
    wire t45795 = t45794 ^ t45794;
    wire t45796 = t45795 ^ t45795;
    wire t45797 = t45796 ^ t45796;
    wire t45798 = t45797 ^ t45797;
    wire t45799 = t45798 ^ t45798;
    wire t45800 = t45799 ^ t45799;
    wire t45801 = t45800 ^ t45800;
    wire t45802 = t45801 ^ t45801;
    wire t45803 = t45802 ^ t45802;
    wire t45804 = t45803 ^ t45803;
    wire t45805 = t45804 ^ t45804;
    wire t45806 = t45805 ^ t45805;
    wire t45807 = t45806 ^ t45806;
    wire t45808 = t45807 ^ t45807;
    wire t45809 = t45808 ^ t45808;
    wire t45810 = t45809 ^ t45809;
    wire t45811 = t45810 ^ t45810;
    wire t45812 = t45811 ^ t45811;
    wire t45813 = t45812 ^ t45812;
    wire t45814 = t45813 ^ t45813;
    wire t45815 = t45814 ^ t45814;
    wire t45816 = t45815 ^ t45815;
    wire t45817 = t45816 ^ t45816;
    wire t45818 = t45817 ^ t45817;
    wire t45819 = t45818 ^ t45818;
    wire t45820 = t45819 ^ t45819;
    wire t45821 = t45820 ^ t45820;
    wire t45822 = t45821 ^ t45821;
    wire t45823 = t45822 ^ t45822;
    wire t45824 = t45823 ^ t45823;
    wire t45825 = t45824 ^ t45824;
    wire t45826 = t45825 ^ t45825;
    wire t45827 = t45826 ^ t45826;
    wire t45828 = t45827 ^ t45827;
    wire t45829 = t45828 ^ t45828;
    wire t45830 = t45829 ^ t45829;
    wire t45831 = t45830 ^ t45830;
    wire t45832 = t45831 ^ t45831;
    wire t45833 = t45832 ^ t45832;
    wire t45834 = t45833 ^ t45833;
    wire t45835 = t45834 ^ t45834;
    wire t45836 = t45835 ^ t45835;
    wire t45837 = t45836 ^ t45836;
    wire t45838 = t45837 ^ t45837;
    wire t45839 = t45838 ^ t45838;
    wire t45840 = t45839 ^ t45839;
    wire t45841 = t45840 ^ t45840;
    wire t45842 = t45841 ^ t45841;
    wire t45843 = t45842 ^ t45842;
    wire t45844 = t45843 ^ t45843;
    wire t45845 = t45844 ^ t45844;
    wire t45846 = t45845 ^ t45845;
    wire t45847 = t45846 ^ t45846;
    wire t45848 = t45847 ^ t45847;
    wire t45849 = t45848 ^ t45848;
    wire t45850 = t45849 ^ t45849;
    wire t45851 = t45850 ^ t45850;
    wire t45852 = t45851 ^ t45851;
    wire t45853 = t45852 ^ t45852;
    wire t45854 = t45853 ^ t45853;
    wire t45855 = t45854 ^ t45854;
    wire t45856 = t45855 ^ t45855;
    wire t45857 = t45856 ^ t45856;
    wire t45858 = t45857 ^ t45857;
    wire t45859 = t45858 ^ t45858;
    wire t45860 = t45859 ^ t45859;
    wire t45861 = t45860 ^ t45860;
    wire t45862 = t45861 ^ t45861;
    wire t45863 = t45862 ^ t45862;
    wire t45864 = t45863 ^ t45863;
    wire t45865 = t45864 ^ t45864;
    wire t45866 = t45865 ^ t45865;
    wire t45867 = t45866 ^ t45866;
    wire t45868 = t45867 ^ t45867;
    wire t45869 = t45868 ^ t45868;
    wire t45870 = t45869 ^ t45869;
    wire t45871 = t45870 ^ t45870;
    wire t45872 = t45871 ^ t45871;
    wire t45873 = t45872 ^ t45872;
    wire t45874 = t45873 ^ t45873;
    wire t45875 = t45874 ^ t45874;
    wire t45876 = t45875 ^ t45875;
    wire t45877 = t45876 ^ t45876;
    wire t45878 = t45877 ^ t45877;
    wire t45879 = t45878 ^ t45878;
    wire t45880 = t45879 ^ t45879;
    wire t45881 = t45880 ^ t45880;
    wire t45882 = t45881 ^ t45881;
    wire t45883 = t45882 ^ t45882;
    wire t45884 = t45883 ^ t45883;
    wire t45885 = t45884 ^ t45884;
    wire t45886 = t45885 ^ t45885;
    wire t45887 = t45886 ^ t45886;
    wire t45888 = t45887 ^ t45887;
    wire t45889 = t45888 ^ t45888;
    wire t45890 = t45889 ^ t45889;
    wire t45891 = t45890 ^ t45890;
    wire t45892 = t45891 ^ t45891;
    wire t45893 = t45892 ^ t45892;
    wire t45894 = t45893 ^ t45893;
    wire t45895 = t45894 ^ t45894;
    wire t45896 = t45895 ^ t45895;
    wire t45897 = t45896 ^ t45896;
    wire t45898 = t45897 ^ t45897;
    wire t45899 = t45898 ^ t45898;
    wire t45900 = t45899 ^ t45899;
    wire t45901 = t45900 ^ t45900;
    wire t45902 = t45901 ^ t45901;
    wire t45903 = t45902 ^ t45902;
    wire t45904 = t45903 ^ t45903;
    wire t45905 = t45904 ^ t45904;
    wire t45906 = t45905 ^ t45905;
    wire t45907 = t45906 ^ t45906;
    wire t45908 = t45907 ^ t45907;
    wire t45909 = t45908 ^ t45908;
    wire t45910 = t45909 ^ t45909;
    wire t45911 = t45910 ^ t45910;
    wire t45912 = t45911 ^ t45911;
    wire t45913 = t45912 ^ t45912;
    wire t45914 = t45913 ^ t45913;
    wire t45915 = t45914 ^ t45914;
    wire t45916 = t45915 ^ t45915;
    wire t45917 = t45916 ^ t45916;
    wire t45918 = t45917 ^ t45917;
    wire t45919 = t45918 ^ t45918;
    wire t45920 = t45919 ^ t45919;
    wire t45921 = t45920 ^ t45920;
    wire t45922 = t45921 ^ t45921;
    wire t45923 = t45922 ^ t45922;
    wire t45924 = t45923 ^ t45923;
    wire t45925 = t45924 ^ t45924;
    wire t45926 = t45925 ^ t45925;
    wire t45927 = t45926 ^ t45926;
    wire t45928 = t45927 ^ t45927;
    wire t45929 = t45928 ^ t45928;
    wire t45930 = t45929 ^ t45929;
    wire t45931 = t45930 ^ t45930;
    wire t45932 = t45931 ^ t45931;
    wire t45933 = t45932 ^ t45932;
    wire t45934 = t45933 ^ t45933;
    wire t45935 = t45934 ^ t45934;
    wire t45936 = t45935 ^ t45935;
    wire t45937 = t45936 ^ t45936;
    wire t45938 = t45937 ^ t45937;
    wire t45939 = t45938 ^ t45938;
    wire t45940 = t45939 ^ t45939;
    wire t45941 = t45940 ^ t45940;
    wire t45942 = t45941 ^ t45941;
    wire t45943 = t45942 ^ t45942;
    wire t45944 = t45943 ^ t45943;
    wire t45945 = t45944 ^ t45944;
    wire t45946 = t45945 ^ t45945;
    wire t45947 = t45946 ^ t45946;
    wire t45948 = t45947 ^ t45947;
    wire t45949 = t45948 ^ t45948;
    wire t45950 = t45949 ^ t45949;
    wire t45951 = t45950 ^ t45950;
    wire t45952 = t45951 ^ t45951;
    wire t45953 = t45952 ^ t45952;
    wire t45954 = t45953 ^ t45953;
    wire t45955 = t45954 ^ t45954;
    wire t45956 = t45955 ^ t45955;
    wire t45957 = t45956 ^ t45956;
    wire t45958 = t45957 ^ t45957;
    wire t45959 = t45958 ^ t45958;
    wire t45960 = t45959 ^ t45959;
    wire t45961 = t45960 ^ t45960;
    wire t45962 = t45961 ^ t45961;
    wire t45963 = t45962 ^ t45962;
    wire t45964 = t45963 ^ t45963;
    wire t45965 = t45964 ^ t45964;
    wire t45966 = t45965 ^ t45965;
    wire t45967 = t45966 ^ t45966;
    wire t45968 = t45967 ^ t45967;
    wire t45969 = t45968 ^ t45968;
    wire t45970 = t45969 ^ t45969;
    wire t45971 = t45970 ^ t45970;
    wire t45972 = t45971 ^ t45971;
    wire t45973 = t45972 ^ t45972;
    wire t45974 = t45973 ^ t45973;
    wire t45975 = t45974 ^ t45974;
    wire t45976 = t45975 ^ t45975;
    wire t45977 = t45976 ^ t45976;
    wire t45978 = t45977 ^ t45977;
    wire t45979 = t45978 ^ t45978;
    wire t45980 = t45979 ^ t45979;
    wire t45981 = t45980 ^ t45980;
    wire t45982 = t45981 ^ t45981;
    wire t45983 = t45982 ^ t45982;
    wire t45984 = t45983 ^ t45983;
    wire t45985 = t45984 ^ t45984;
    wire t45986 = t45985 ^ t45985;
    wire t45987 = t45986 ^ t45986;
    wire t45988 = t45987 ^ t45987;
    wire t45989 = t45988 ^ t45988;
    wire t45990 = t45989 ^ t45989;
    wire t45991 = t45990 ^ t45990;
    wire t45992 = t45991 ^ t45991;
    wire t45993 = t45992 ^ t45992;
    wire t45994 = t45993 ^ t45993;
    wire t45995 = t45994 ^ t45994;
    wire t45996 = t45995 ^ t45995;
    wire t45997 = t45996 ^ t45996;
    wire t45998 = t45997 ^ t45997;
    wire t45999 = t45998 ^ t45998;
    wire t46000 = t45999 ^ t45999;
    wire t46001 = t46000 ^ t46000;
    wire t46002 = t46001 ^ t46001;
    wire t46003 = t46002 ^ t46002;
    wire t46004 = t46003 ^ t46003;
    wire t46005 = t46004 ^ t46004;
    wire t46006 = t46005 ^ t46005;
    wire t46007 = t46006 ^ t46006;
    wire t46008 = t46007 ^ t46007;
    wire t46009 = t46008 ^ t46008;
    wire t46010 = t46009 ^ t46009;
    wire t46011 = t46010 ^ t46010;
    wire t46012 = t46011 ^ t46011;
    wire t46013 = t46012 ^ t46012;
    wire t46014 = t46013 ^ t46013;
    wire t46015 = t46014 ^ t46014;
    wire t46016 = t46015 ^ t46015;
    wire t46017 = t46016 ^ t46016;
    wire t46018 = t46017 ^ t46017;
    wire t46019 = t46018 ^ t46018;
    wire t46020 = t46019 ^ t46019;
    wire t46021 = t46020 ^ t46020;
    wire t46022 = t46021 ^ t46021;
    wire t46023 = t46022 ^ t46022;
    wire t46024 = t46023 ^ t46023;
    wire t46025 = t46024 ^ t46024;
    wire t46026 = t46025 ^ t46025;
    wire t46027 = t46026 ^ t46026;
    wire t46028 = t46027 ^ t46027;
    wire t46029 = t46028 ^ t46028;
    wire t46030 = t46029 ^ t46029;
    wire t46031 = t46030 ^ t46030;
    wire t46032 = t46031 ^ t46031;
    wire t46033 = t46032 ^ t46032;
    wire t46034 = t46033 ^ t46033;
    wire t46035 = t46034 ^ t46034;
    wire t46036 = t46035 ^ t46035;
    wire t46037 = t46036 ^ t46036;
    wire t46038 = t46037 ^ t46037;
    wire t46039 = t46038 ^ t46038;
    wire t46040 = t46039 ^ t46039;
    wire t46041 = t46040 ^ t46040;
    wire t46042 = t46041 ^ t46041;
    wire t46043 = t46042 ^ t46042;
    wire t46044 = t46043 ^ t46043;
    wire t46045 = t46044 ^ t46044;
    wire t46046 = t46045 ^ t46045;
    wire t46047 = t46046 ^ t46046;
    wire t46048 = t46047 ^ t46047;
    wire t46049 = t46048 ^ t46048;
    wire t46050 = t46049 ^ t46049;
    wire t46051 = t46050 ^ t46050;
    wire t46052 = t46051 ^ t46051;
    wire t46053 = t46052 ^ t46052;
    wire t46054 = t46053 ^ t46053;
    wire t46055 = t46054 ^ t46054;
    wire t46056 = t46055 ^ t46055;
    wire t46057 = t46056 ^ t46056;
    wire t46058 = t46057 ^ t46057;
    wire t46059 = t46058 ^ t46058;
    wire t46060 = t46059 ^ t46059;
    wire t46061 = t46060 ^ t46060;
    wire t46062 = t46061 ^ t46061;
    wire t46063 = t46062 ^ t46062;
    wire t46064 = t46063 ^ t46063;
    wire t46065 = t46064 ^ t46064;
    wire t46066 = t46065 ^ t46065;
    wire t46067 = t46066 ^ t46066;
    wire t46068 = t46067 ^ t46067;
    wire t46069 = t46068 ^ t46068;
    wire t46070 = t46069 ^ t46069;
    wire t46071 = t46070 ^ t46070;
    wire t46072 = t46071 ^ t46071;
    wire t46073 = t46072 ^ t46072;
    wire t46074 = t46073 ^ t46073;
    wire t46075 = t46074 ^ t46074;
    wire t46076 = t46075 ^ t46075;
    wire t46077 = t46076 ^ t46076;
    wire t46078 = t46077 ^ t46077;
    wire t46079 = t46078 ^ t46078;
    wire t46080 = t46079 ^ t46079;
    wire t46081 = t46080 ^ t46080;
    wire t46082 = t46081 ^ t46081;
    wire t46083 = t46082 ^ t46082;
    wire t46084 = t46083 ^ t46083;
    wire t46085 = t46084 ^ t46084;
    wire t46086 = t46085 ^ t46085;
    wire t46087 = t46086 ^ t46086;
    wire t46088 = t46087 ^ t46087;
    wire t46089 = t46088 ^ t46088;
    wire t46090 = t46089 ^ t46089;
    wire t46091 = t46090 ^ t46090;
    wire t46092 = t46091 ^ t46091;
    wire t46093 = t46092 ^ t46092;
    wire t46094 = t46093 ^ t46093;
    wire t46095 = t46094 ^ t46094;
    wire t46096 = t46095 ^ t46095;
    wire t46097 = t46096 ^ t46096;
    wire t46098 = t46097 ^ t46097;
    wire t46099 = t46098 ^ t46098;
    wire t46100 = t46099 ^ t46099;
    wire t46101 = t46100 ^ t46100;
    wire t46102 = t46101 ^ t46101;
    wire t46103 = t46102 ^ t46102;
    wire t46104 = t46103 ^ t46103;
    wire t46105 = t46104 ^ t46104;
    wire t46106 = t46105 ^ t46105;
    wire t46107 = t46106 ^ t46106;
    wire t46108 = t46107 ^ t46107;
    wire t46109 = t46108 ^ t46108;
    wire t46110 = t46109 ^ t46109;
    wire t46111 = t46110 ^ t46110;
    wire t46112 = t46111 ^ t46111;
    wire t46113 = t46112 ^ t46112;
    wire t46114 = t46113 ^ t46113;
    wire t46115 = t46114 ^ t46114;
    wire t46116 = t46115 ^ t46115;
    wire t46117 = t46116 ^ t46116;
    wire t46118 = t46117 ^ t46117;
    wire t46119 = t46118 ^ t46118;
    wire t46120 = t46119 ^ t46119;
    wire t46121 = t46120 ^ t46120;
    wire t46122 = t46121 ^ t46121;
    wire t46123 = t46122 ^ t46122;
    wire t46124 = t46123 ^ t46123;
    wire t46125 = t46124 ^ t46124;
    wire t46126 = t46125 ^ t46125;
    wire t46127 = t46126 ^ t46126;
    wire t46128 = t46127 ^ t46127;
    wire t46129 = t46128 ^ t46128;
    wire t46130 = t46129 ^ t46129;
    wire t46131 = t46130 ^ t46130;
    wire t46132 = t46131 ^ t46131;
    wire t46133 = t46132 ^ t46132;
    wire t46134 = t46133 ^ t46133;
    wire t46135 = t46134 ^ t46134;
    wire t46136 = t46135 ^ t46135;
    wire t46137 = t46136 ^ t46136;
    wire t46138 = t46137 ^ t46137;
    wire t46139 = t46138 ^ t46138;
    wire t46140 = t46139 ^ t46139;
    wire t46141 = t46140 ^ t46140;
    wire t46142 = t46141 ^ t46141;
    wire t46143 = t46142 ^ t46142;
    wire t46144 = t46143 ^ t46143;
    wire t46145 = t46144 ^ t46144;
    wire t46146 = t46145 ^ t46145;
    wire t46147 = t46146 ^ t46146;
    wire t46148 = t46147 ^ t46147;
    wire t46149 = t46148 ^ t46148;
    wire t46150 = t46149 ^ t46149;
    wire t46151 = t46150 ^ t46150;
    wire t46152 = t46151 ^ t46151;
    wire t46153 = t46152 ^ t46152;
    wire t46154 = t46153 ^ t46153;
    wire t46155 = t46154 ^ t46154;
    wire t46156 = t46155 ^ t46155;
    wire t46157 = t46156 ^ t46156;
    wire t46158 = t46157 ^ t46157;
    wire t46159 = t46158 ^ t46158;
    wire t46160 = t46159 ^ t46159;
    wire t46161 = t46160 ^ t46160;
    wire t46162 = t46161 ^ t46161;
    wire t46163 = t46162 ^ t46162;
    wire t46164 = t46163 ^ t46163;
    wire t46165 = t46164 ^ t46164;
    wire t46166 = t46165 ^ t46165;
    wire t46167 = t46166 ^ t46166;
    wire t46168 = t46167 ^ t46167;
    wire t46169 = t46168 ^ t46168;
    wire t46170 = t46169 ^ t46169;
    wire t46171 = t46170 ^ t46170;
    wire t46172 = t46171 ^ t46171;
    wire t46173 = t46172 ^ t46172;
    wire t46174 = t46173 ^ t46173;
    wire t46175 = t46174 ^ t46174;
    wire t46176 = t46175 ^ t46175;
    wire t46177 = t46176 ^ t46176;
    wire t46178 = t46177 ^ t46177;
    wire t46179 = t46178 ^ t46178;
    wire t46180 = t46179 ^ t46179;
    wire t46181 = t46180 ^ t46180;
    wire t46182 = t46181 ^ t46181;
    wire t46183 = t46182 ^ t46182;
    wire t46184 = t46183 ^ t46183;
    wire t46185 = t46184 ^ t46184;
    wire t46186 = t46185 ^ t46185;
    wire t46187 = t46186 ^ t46186;
    wire t46188 = t46187 ^ t46187;
    wire t46189 = t46188 ^ t46188;
    wire t46190 = t46189 ^ t46189;
    wire t46191 = t46190 ^ t46190;
    wire t46192 = t46191 ^ t46191;
    wire t46193 = t46192 ^ t46192;
    wire t46194 = t46193 ^ t46193;
    wire t46195 = t46194 ^ t46194;
    wire t46196 = t46195 ^ t46195;
    wire t46197 = t46196 ^ t46196;
    wire t46198 = t46197 ^ t46197;
    wire t46199 = t46198 ^ t46198;
    wire t46200 = t46199 ^ t46199;
    wire t46201 = t46200 ^ t46200;
    wire t46202 = t46201 ^ t46201;
    wire t46203 = t46202 ^ t46202;
    wire t46204 = t46203 ^ t46203;
    wire t46205 = t46204 ^ t46204;
    wire t46206 = t46205 ^ t46205;
    wire t46207 = t46206 ^ t46206;
    wire t46208 = t46207 ^ t46207;
    wire t46209 = t46208 ^ t46208;
    wire t46210 = t46209 ^ t46209;
    wire t46211 = t46210 ^ t46210;
    wire t46212 = t46211 ^ t46211;
    wire t46213 = t46212 ^ t46212;
    wire t46214 = t46213 ^ t46213;
    wire t46215 = t46214 ^ t46214;
    wire t46216 = t46215 ^ t46215;
    wire t46217 = t46216 ^ t46216;
    wire t46218 = t46217 ^ t46217;
    wire t46219 = t46218 ^ t46218;
    wire t46220 = t46219 ^ t46219;
    wire t46221 = t46220 ^ t46220;
    wire t46222 = t46221 ^ t46221;
    wire t46223 = t46222 ^ t46222;
    wire t46224 = t46223 ^ t46223;
    wire t46225 = t46224 ^ t46224;
    wire t46226 = t46225 ^ t46225;
    wire t46227 = t46226 ^ t46226;
    wire t46228 = t46227 ^ t46227;
    wire t46229 = t46228 ^ t46228;
    wire t46230 = t46229 ^ t46229;
    wire t46231 = t46230 ^ t46230;
    wire t46232 = t46231 ^ t46231;
    wire t46233 = t46232 ^ t46232;
    wire t46234 = t46233 ^ t46233;
    wire t46235 = t46234 ^ t46234;
    wire t46236 = t46235 ^ t46235;
    wire t46237 = t46236 ^ t46236;
    wire t46238 = t46237 ^ t46237;
    wire t46239 = t46238 ^ t46238;
    wire t46240 = t46239 ^ t46239;
    wire t46241 = t46240 ^ t46240;
    wire t46242 = t46241 ^ t46241;
    wire t46243 = t46242 ^ t46242;
    wire t46244 = t46243 ^ t46243;
    wire t46245 = t46244 ^ t46244;
    wire t46246 = t46245 ^ t46245;
    wire t46247 = t46246 ^ t46246;
    wire t46248 = t46247 ^ t46247;
    wire t46249 = t46248 ^ t46248;
    wire t46250 = t46249 ^ t46249;
    wire t46251 = t46250 ^ t46250;
    wire t46252 = t46251 ^ t46251;
    wire t46253 = t46252 ^ t46252;
    wire t46254 = t46253 ^ t46253;
    wire t46255 = t46254 ^ t46254;
    wire t46256 = t46255 ^ t46255;
    wire t46257 = t46256 ^ t46256;
    wire t46258 = t46257 ^ t46257;
    wire t46259 = t46258 ^ t46258;
    wire t46260 = t46259 ^ t46259;
    wire t46261 = t46260 ^ t46260;
    wire t46262 = t46261 ^ t46261;
    wire t46263 = t46262 ^ t46262;
    wire t46264 = t46263 ^ t46263;
    wire t46265 = t46264 ^ t46264;
    wire t46266 = t46265 ^ t46265;
    wire t46267 = t46266 ^ t46266;
    wire t46268 = t46267 ^ t46267;
    wire t46269 = t46268 ^ t46268;
    wire t46270 = t46269 ^ t46269;
    wire t46271 = t46270 ^ t46270;
    wire t46272 = t46271 ^ t46271;
    wire t46273 = t46272 ^ t46272;
    wire t46274 = t46273 ^ t46273;
    wire t46275 = t46274 ^ t46274;
    wire t46276 = t46275 ^ t46275;
    wire t46277 = t46276 ^ t46276;
    wire t46278 = t46277 ^ t46277;
    wire t46279 = t46278 ^ t46278;
    wire t46280 = t46279 ^ t46279;
    wire t46281 = t46280 ^ t46280;
    wire t46282 = t46281 ^ t46281;
    wire t46283 = t46282 ^ t46282;
    wire t46284 = t46283 ^ t46283;
    wire t46285 = t46284 ^ t46284;
    wire t46286 = t46285 ^ t46285;
    wire t46287 = t46286 ^ t46286;
    wire t46288 = t46287 ^ t46287;
    wire t46289 = t46288 ^ t46288;
    wire t46290 = t46289 ^ t46289;
    wire t46291 = t46290 ^ t46290;
    wire t46292 = t46291 ^ t46291;
    wire t46293 = t46292 ^ t46292;
    wire t46294 = t46293 ^ t46293;
    wire t46295 = t46294 ^ t46294;
    wire t46296 = t46295 ^ t46295;
    wire t46297 = t46296 ^ t46296;
    wire t46298 = t46297 ^ t46297;
    wire t46299 = t46298 ^ t46298;
    wire t46300 = t46299 ^ t46299;
    wire t46301 = t46300 ^ t46300;
    wire t46302 = t46301 ^ t46301;
    wire t46303 = t46302 ^ t46302;
    wire t46304 = t46303 ^ t46303;
    wire t46305 = t46304 ^ t46304;
    wire t46306 = t46305 ^ t46305;
    wire t46307 = t46306 ^ t46306;
    wire t46308 = t46307 ^ t46307;
    wire t46309 = t46308 ^ t46308;
    wire t46310 = t46309 ^ t46309;
    wire t46311 = t46310 ^ t46310;
    wire t46312 = t46311 ^ t46311;
    wire t46313 = t46312 ^ t46312;
    wire t46314 = t46313 ^ t46313;
    wire t46315 = t46314 ^ t46314;
    wire t46316 = t46315 ^ t46315;
    wire t46317 = t46316 ^ t46316;
    wire t46318 = t46317 ^ t46317;
    wire t46319 = t46318 ^ t46318;
    wire t46320 = t46319 ^ t46319;
    wire t46321 = t46320 ^ t46320;
    wire t46322 = t46321 ^ t46321;
    wire t46323 = t46322 ^ t46322;
    wire t46324 = t46323 ^ t46323;
    wire t46325 = t46324 ^ t46324;
    wire t46326 = t46325 ^ t46325;
    wire t46327 = t46326 ^ t46326;
    wire t46328 = t46327 ^ t46327;
    wire t46329 = t46328 ^ t46328;
    wire t46330 = t46329 ^ t46329;
    wire t46331 = t46330 ^ t46330;
    wire t46332 = t46331 ^ t46331;
    wire t46333 = t46332 ^ t46332;
    wire t46334 = t46333 ^ t46333;
    wire t46335 = t46334 ^ t46334;
    wire t46336 = t46335 ^ t46335;
    wire t46337 = t46336 ^ t46336;
    wire t46338 = t46337 ^ t46337;
    wire t46339 = t46338 ^ t46338;
    wire t46340 = t46339 ^ t46339;
    wire t46341 = t46340 ^ t46340;
    wire t46342 = t46341 ^ t46341;
    wire t46343 = t46342 ^ t46342;
    wire t46344 = t46343 ^ t46343;
    wire t46345 = t46344 ^ t46344;
    wire t46346 = t46345 ^ t46345;
    wire t46347 = t46346 ^ t46346;
    wire t46348 = t46347 ^ t46347;
    wire t46349 = t46348 ^ t46348;
    wire t46350 = t46349 ^ t46349;
    wire t46351 = t46350 ^ t46350;
    wire t46352 = t46351 ^ t46351;
    wire t46353 = t46352 ^ t46352;
    wire t46354 = t46353 ^ t46353;
    wire t46355 = t46354 ^ t46354;
    wire t46356 = t46355 ^ t46355;
    wire t46357 = t46356 ^ t46356;
    wire t46358 = t46357 ^ t46357;
    wire t46359 = t46358 ^ t46358;
    wire t46360 = t46359 ^ t46359;
    wire t46361 = t46360 ^ t46360;
    wire t46362 = t46361 ^ t46361;
    wire t46363 = t46362 ^ t46362;
    wire t46364 = t46363 ^ t46363;
    wire t46365 = t46364 ^ t46364;
    wire t46366 = t46365 ^ t46365;
    wire t46367 = t46366 ^ t46366;
    wire t46368 = t46367 ^ t46367;
    wire t46369 = t46368 ^ t46368;
    wire t46370 = t46369 ^ t46369;
    wire t46371 = t46370 ^ t46370;
    wire t46372 = t46371 ^ t46371;
    wire t46373 = t46372 ^ t46372;
    wire t46374 = t46373 ^ t46373;
    wire t46375 = t46374 ^ t46374;
    wire t46376 = t46375 ^ t46375;
    wire t46377 = t46376 ^ t46376;
    wire t46378 = t46377 ^ t46377;
    wire t46379 = t46378 ^ t46378;
    wire t46380 = t46379 ^ t46379;
    wire t46381 = t46380 ^ t46380;
    wire t46382 = t46381 ^ t46381;
    wire t46383 = t46382 ^ t46382;
    wire t46384 = t46383 ^ t46383;
    wire t46385 = t46384 ^ t46384;
    wire t46386 = t46385 ^ t46385;
    wire t46387 = t46386 ^ t46386;
    wire t46388 = t46387 ^ t46387;
    wire t46389 = t46388 ^ t46388;
    wire t46390 = t46389 ^ t46389;
    wire t46391 = t46390 ^ t46390;
    wire t46392 = t46391 ^ t46391;
    wire t46393 = t46392 ^ t46392;
    wire t46394 = t46393 ^ t46393;
    wire t46395 = t46394 ^ t46394;
    wire t46396 = t46395 ^ t46395;
    wire t46397 = t46396 ^ t46396;
    wire t46398 = t46397 ^ t46397;
    wire t46399 = t46398 ^ t46398;
    wire t46400 = t46399 ^ t46399;
    wire t46401 = t46400 ^ t46400;
    wire t46402 = t46401 ^ t46401;
    wire t46403 = t46402 ^ t46402;
    wire t46404 = t46403 ^ t46403;
    wire t46405 = t46404 ^ t46404;
    wire t46406 = t46405 ^ t46405;
    wire t46407 = t46406 ^ t46406;
    wire t46408 = t46407 ^ t46407;
    wire t46409 = t46408 ^ t46408;
    wire t46410 = t46409 ^ t46409;
    wire t46411 = t46410 ^ t46410;
    wire t46412 = t46411 ^ t46411;
    wire t46413 = t46412 ^ t46412;
    wire t46414 = t46413 ^ t46413;
    wire t46415 = t46414 ^ t46414;
    wire t46416 = t46415 ^ t46415;
    wire t46417 = t46416 ^ t46416;
    wire t46418 = t46417 ^ t46417;
    wire t46419 = t46418 ^ t46418;
    wire t46420 = t46419 ^ t46419;
    wire t46421 = t46420 ^ t46420;
    wire t46422 = t46421 ^ t46421;
    wire t46423 = t46422 ^ t46422;
    wire t46424 = t46423 ^ t46423;
    wire t46425 = t46424 ^ t46424;
    wire t46426 = t46425 ^ t46425;
    wire t46427 = t46426 ^ t46426;
    wire t46428 = t46427 ^ t46427;
    wire t46429 = t46428 ^ t46428;
    wire t46430 = t46429 ^ t46429;
    wire t46431 = t46430 ^ t46430;
    wire t46432 = t46431 ^ t46431;
    wire t46433 = t46432 ^ t46432;
    wire t46434 = t46433 ^ t46433;
    wire t46435 = t46434 ^ t46434;
    wire t46436 = t46435 ^ t46435;
    wire t46437 = t46436 ^ t46436;
    wire t46438 = t46437 ^ t46437;
    wire t46439 = t46438 ^ t46438;
    wire t46440 = t46439 ^ t46439;
    wire t46441 = t46440 ^ t46440;
    wire t46442 = t46441 ^ t46441;
    wire t46443 = t46442 ^ t46442;
    wire t46444 = t46443 ^ t46443;
    wire t46445 = t46444 ^ t46444;
    wire t46446 = t46445 ^ t46445;
    wire t46447 = t46446 ^ t46446;
    wire t46448 = t46447 ^ t46447;
    wire t46449 = t46448 ^ t46448;
    wire t46450 = t46449 ^ t46449;
    wire t46451 = t46450 ^ t46450;
    wire t46452 = t46451 ^ t46451;
    wire t46453 = t46452 ^ t46452;
    wire t46454 = t46453 ^ t46453;
    wire t46455 = t46454 ^ t46454;
    wire t46456 = t46455 ^ t46455;
    wire t46457 = t46456 ^ t46456;
    wire t46458 = t46457 ^ t46457;
    wire t46459 = t46458 ^ t46458;
    wire t46460 = t46459 ^ t46459;
    wire t46461 = t46460 ^ t46460;
    wire t46462 = t46461 ^ t46461;
    wire t46463 = t46462 ^ t46462;
    wire t46464 = t46463 ^ t46463;
    wire t46465 = t46464 ^ t46464;
    wire t46466 = t46465 ^ t46465;
    wire t46467 = t46466 ^ t46466;
    wire t46468 = t46467 ^ t46467;
    wire t46469 = t46468 ^ t46468;
    wire t46470 = t46469 ^ t46469;
    wire t46471 = t46470 ^ t46470;
    wire t46472 = t46471 ^ t46471;
    wire t46473 = t46472 ^ t46472;
    wire t46474 = t46473 ^ t46473;
    wire t46475 = t46474 ^ t46474;
    wire t46476 = t46475 ^ t46475;
    wire t46477 = t46476 ^ t46476;
    wire t46478 = t46477 ^ t46477;
    wire t46479 = t46478 ^ t46478;
    wire t46480 = t46479 ^ t46479;
    wire t46481 = t46480 ^ t46480;
    wire t46482 = t46481 ^ t46481;
    wire t46483 = t46482 ^ t46482;
    wire t46484 = t46483 ^ t46483;
    wire t46485 = t46484 ^ t46484;
    wire t46486 = t46485 ^ t46485;
    wire t46487 = t46486 ^ t46486;
    wire t46488 = t46487 ^ t46487;
    wire t46489 = t46488 ^ t46488;
    wire t46490 = t46489 ^ t46489;
    wire t46491 = t46490 ^ t46490;
    wire t46492 = t46491 ^ t46491;
    wire t46493 = t46492 ^ t46492;
    wire t46494 = t46493 ^ t46493;
    wire t46495 = t46494 ^ t46494;
    wire t46496 = t46495 ^ t46495;
    wire t46497 = t46496 ^ t46496;
    wire t46498 = t46497 ^ t46497;
    wire t46499 = t46498 ^ t46498;
    wire t46500 = t46499 ^ t46499;
    wire t46501 = t46500 ^ t46500;
    wire t46502 = t46501 ^ t46501;
    wire t46503 = t46502 ^ t46502;
    wire t46504 = t46503 ^ t46503;
    wire t46505 = t46504 ^ t46504;
    wire t46506 = t46505 ^ t46505;
    wire t46507 = t46506 ^ t46506;
    wire t46508 = t46507 ^ t46507;
    wire t46509 = t46508 ^ t46508;
    wire t46510 = t46509 ^ t46509;
    wire t46511 = t46510 ^ t46510;
    wire t46512 = t46511 ^ t46511;
    wire t46513 = t46512 ^ t46512;
    wire t46514 = t46513 ^ t46513;
    wire t46515 = t46514 ^ t46514;
    wire t46516 = t46515 ^ t46515;
    wire t46517 = t46516 ^ t46516;
    wire t46518 = t46517 ^ t46517;
    wire t46519 = t46518 ^ t46518;
    wire t46520 = t46519 ^ t46519;
    wire t46521 = t46520 ^ t46520;
    wire t46522 = t46521 ^ t46521;
    wire t46523 = t46522 ^ t46522;
    wire t46524 = t46523 ^ t46523;
    wire t46525 = t46524 ^ t46524;
    wire t46526 = t46525 ^ t46525;
    wire t46527 = t46526 ^ t46526;
    wire t46528 = t46527 ^ t46527;
    wire t46529 = t46528 ^ t46528;
    wire t46530 = t46529 ^ t46529;
    wire t46531 = t46530 ^ t46530;
    wire t46532 = t46531 ^ t46531;
    wire t46533 = t46532 ^ t46532;
    wire t46534 = t46533 ^ t46533;
    wire t46535 = t46534 ^ t46534;
    wire t46536 = t46535 ^ t46535;
    wire t46537 = t46536 ^ t46536;
    wire t46538 = t46537 ^ t46537;
    wire t46539 = t46538 ^ t46538;
    wire t46540 = t46539 ^ t46539;
    wire t46541 = t46540 ^ t46540;
    wire t46542 = t46541 ^ t46541;
    wire t46543 = t46542 ^ t46542;
    wire t46544 = t46543 ^ t46543;
    wire t46545 = t46544 ^ t46544;
    wire t46546 = t46545 ^ t46545;
    wire t46547 = t46546 ^ t46546;
    wire t46548 = t46547 ^ t46547;
    wire t46549 = t46548 ^ t46548;
    wire t46550 = t46549 ^ t46549;
    wire t46551 = t46550 ^ t46550;
    wire t46552 = t46551 ^ t46551;
    wire t46553 = t46552 ^ t46552;
    wire t46554 = t46553 ^ t46553;
    wire t46555 = t46554 ^ t46554;
    wire t46556 = t46555 ^ t46555;
    wire t46557 = t46556 ^ t46556;
    wire t46558 = t46557 ^ t46557;
    wire t46559 = t46558 ^ t46558;
    wire t46560 = t46559 ^ t46559;
    wire t46561 = t46560 ^ t46560;
    wire t46562 = t46561 ^ t46561;
    wire t46563 = t46562 ^ t46562;
    wire t46564 = t46563 ^ t46563;
    wire t46565 = t46564 ^ t46564;
    wire t46566 = t46565 ^ t46565;
    wire t46567 = t46566 ^ t46566;
    wire t46568 = t46567 ^ t46567;
    wire t46569 = t46568 ^ t46568;
    wire t46570 = t46569 ^ t46569;
    wire t46571 = t46570 ^ t46570;
    wire t46572 = t46571 ^ t46571;
    wire t46573 = t46572 ^ t46572;
    wire t46574 = t46573 ^ t46573;
    wire t46575 = t46574 ^ t46574;
    wire t46576 = t46575 ^ t46575;
    wire t46577 = t46576 ^ t46576;
    wire t46578 = t46577 ^ t46577;
    wire t46579 = t46578 ^ t46578;
    wire t46580 = t46579 ^ t46579;
    wire t46581 = t46580 ^ t46580;
    wire t46582 = t46581 ^ t46581;
    wire t46583 = t46582 ^ t46582;
    wire t46584 = t46583 ^ t46583;
    wire t46585 = t46584 ^ t46584;
    wire t46586 = t46585 ^ t46585;
    wire t46587 = t46586 ^ t46586;
    wire t46588 = t46587 ^ t46587;
    wire t46589 = t46588 ^ t46588;
    wire t46590 = t46589 ^ t46589;
    wire t46591 = t46590 ^ t46590;
    wire t46592 = t46591 ^ t46591;
    wire t46593 = t46592 ^ t46592;
    wire t46594 = t46593 ^ t46593;
    wire t46595 = t46594 ^ t46594;
    wire t46596 = t46595 ^ t46595;
    wire t46597 = t46596 ^ t46596;
    wire t46598 = t46597 ^ t46597;
    wire t46599 = t46598 ^ t46598;
    wire t46600 = t46599 ^ t46599;
    wire t46601 = t46600 ^ t46600;
    wire t46602 = t46601 ^ t46601;
    wire t46603 = t46602 ^ t46602;
    wire t46604 = t46603 ^ t46603;
    wire t46605 = t46604 ^ t46604;
    wire t46606 = t46605 ^ t46605;
    wire t46607 = t46606 ^ t46606;
    wire t46608 = t46607 ^ t46607;
    wire t46609 = t46608 ^ t46608;
    wire t46610 = t46609 ^ t46609;
    wire t46611 = t46610 ^ t46610;
    wire t46612 = t46611 ^ t46611;
    wire t46613 = t46612 ^ t46612;
    wire t46614 = t46613 ^ t46613;
    wire t46615 = t46614 ^ t46614;
    wire t46616 = t46615 ^ t46615;
    wire t46617 = t46616 ^ t46616;
    wire t46618 = t46617 ^ t46617;
    wire t46619 = t46618 ^ t46618;
    wire t46620 = t46619 ^ t46619;
    wire t46621 = t46620 ^ t46620;
    wire t46622 = t46621 ^ t46621;
    wire t46623 = t46622 ^ t46622;
    wire t46624 = t46623 ^ t46623;
    wire t46625 = t46624 ^ t46624;
    wire t46626 = t46625 ^ t46625;
    wire t46627 = t46626 ^ t46626;
    wire t46628 = t46627 ^ t46627;
    wire t46629 = t46628 ^ t46628;
    wire t46630 = t46629 ^ t46629;
    wire t46631 = t46630 ^ t46630;
    wire t46632 = t46631 ^ t46631;
    wire t46633 = t46632 ^ t46632;
    wire t46634 = t46633 ^ t46633;
    wire t46635 = t46634 ^ t46634;
    wire t46636 = t46635 ^ t46635;
    wire t46637 = t46636 ^ t46636;
    wire t46638 = t46637 ^ t46637;
    wire t46639 = t46638 ^ t46638;
    wire t46640 = t46639 ^ t46639;
    wire t46641 = t46640 ^ t46640;
    wire t46642 = t46641 ^ t46641;
    wire t46643 = t46642 ^ t46642;
    wire t46644 = t46643 ^ t46643;
    wire t46645 = t46644 ^ t46644;
    wire t46646 = t46645 ^ t46645;
    wire t46647 = t46646 ^ t46646;
    wire t46648 = t46647 ^ t46647;
    wire t46649 = t46648 ^ t46648;
    wire t46650 = t46649 ^ t46649;
    wire t46651 = t46650 ^ t46650;
    wire t46652 = t46651 ^ t46651;
    wire t46653 = t46652 ^ t46652;
    wire t46654 = t46653 ^ t46653;
    wire t46655 = t46654 ^ t46654;
    wire t46656 = t46655 ^ t46655;
    wire t46657 = t46656 ^ t46656;
    wire t46658 = t46657 ^ t46657;
    wire t46659 = t46658 ^ t46658;
    wire t46660 = t46659 ^ t46659;
    wire t46661 = t46660 ^ t46660;
    wire t46662 = t46661 ^ t46661;
    wire t46663 = t46662 ^ t46662;
    wire t46664 = t46663 ^ t46663;
    wire t46665 = t46664 ^ t46664;
    wire t46666 = t46665 ^ t46665;
    wire t46667 = t46666 ^ t46666;
    wire t46668 = t46667 ^ t46667;
    wire t46669 = t46668 ^ t46668;
    wire t46670 = t46669 ^ t46669;
    wire t46671 = t46670 ^ t46670;
    wire t46672 = t46671 ^ t46671;
    wire t46673 = t46672 ^ t46672;
    wire t46674 = t46673 ^ t46673;
    wire t46675 = t46674 ^ t46674;
    wire t46676 = t46675 ^ t46675;
    wire t46677 = t46676 ^ t46676;
    wire t46678 = t46677 ^ t46677;
    wire t46679 = t46678 ^ t46678;
    wire t46680 = t46679 ^ t46679;
    wire t46681 = t46680 ^ t46680;
    wire t46682 = t46681 ^ t46681;
    wire t46683 = t46682 ^ t46682;
    wire t46684 = t46683 ^ t46683;
    wire t46685 = t46684 ^ t46684;
    wire t46686 = t46685 ^ t46685;
    wire t46687 = t46686 ^ t46686;
    wire t46688 = t46687 ^ t46687;
    wire t46689 = t46688 ^ t46688;
    wire t46690 = t46689 ^ t46689;
    wire t46691 = t46690 ^ t46690;
    wire t46692 = t46691 ^ t46691;
    wire t46693 = t46692 ^ t46692;
    wire t46694 = t46693 ^ t46693;
    wire t46695 = t46694 ^ t46694;
    wire t46696 = t46695 ^ t46695;
    wire t46697 = t46696 ^ t46696;
    wire t46698 = t46697 ^ t46697;
    wire t46699 = t46698 ^ t46698;
    wire t46700 = t46699 ^ t46699;
    wire t46701 = t46700 ^ t46700;
    wire t46702 = t46701 ^ t46701;
    wire t46703 = t46702 ^ t46702;
    wire t46704 = t46703 ^ t46703;
    wire t46705 = t46704 ^ t46704;
    wire t46706 = t46705 ^ t46705;
    wire t46707 = t46706 ^ t46706;
    wire t46708 = t46707 ^ t46707;
    wire t46709 = t46708 ^ t46708;
    wire t46710 = t46709 ^ t46709;
    wire t46711 = t46710 ^ t46710;
    wire t46712 = t46711 ^ t46711;
    wire t46713 = t46712 ^ t46712;
    wire t46714 = t46713 ^ t46713;
    wire t46715 = t46714 ^ t46714;
    wire t46716 = t46715 ^ t46715;
    wire t46717 = t46716 ^ t46716;
    wire t46718 = t46717 ^ t46717;
    wire t46719 = t46718 ^ t46718;
    wire t46720 = t46719 ^ t46719;
    wire t46721 = t46720 ^ t46720;
    wire t46722 = t46721 ^ t46721;
    wire t46723 = t46722 ^ t46722;
    wire t46724 = t46723 ^ t46723;
    wire t46725 = t46724 ^ t46724;
    wire t46726 = t46725 ^ t46725;
    wire t46727 = t46726 ^ t46726;
    wire t46728 = t46727 ^ t46727;
    wire t46729 = t46728 ^ t46728;
    wire t46730 = t46729 ^ t46729;
    wire t46731 = t46730 ^ t46730;
    wire t46732 = t46731 ^ t46731;
    wire t46733 = t46732 ^ t46732;
    wire t46734 = t46733 ^ t46733;
    wire t46735 = t46734 ^ t46734;
    wire t46736 = t46735 ^ t46735;
    wire t46737 = t46736 ^ t46736;
    wire t46738 = t46737 ^ t46737;
    wire t46739 = t46738 ^ t46738;
    wire t46740 = t46739 ^ t46739;
    wire t46741 = t46740 ^ t46740;
    wire t46742 = t46741 ^ t46741;
    wire t46743 = t46742 ^ t46742;
    wire t46744 = t46743 ^ t46743;
    wire t46745 = t46744 ^ t46744;
    wire t46746 = t46745 ^ t46745;
    wire t46747 = t46746 ^ t46746;
    wire t46748 = t46747 ^ t46747;
    wire t46749 = t46748 ^ t46748;
    wire t46750 = t46749 ^ t46749;
    wire t46751 = t46750 ^ t46750;
    wire t46752 = t46751 ^ t46751;
    wire t46753 = t46752 ^ t46752;
    wire t46754 = t46753 ^ t46753;
    wire t46755 = t46754 ^ t46754;
    wire t46756 = t46755 ^ t46755;
    wire t46757 = t46756 ^ t46756;
    wire t46758 = t46757 ^ t46757;
    wire t46759 = t46758 ^ t46758;
    wire t46760 = t46759 ^ t46759;
    wire t46761 = t46760 ^ t46760;
    wire t46762 = t46761 ^ t46761;
    wire t46763 = t46762 ^ t46762;
    wire t46764 = t46763 ^ t46763;
    wire t46765 = t46764 ^ t46764;
    wire t46766 = t46765 ^ t46765;
    wire t46767 = t46766 ^ t46766;
    wire t46768 = t46767 ^ t46767;
    wire t46769 = t46768 ^ t46768;
    wire t46770 = t46769 ^ t46769;
    wire t46771 = t46770 ^ t46770;
    wire t46772 = t46771 ^ t46771;
    wire t46773 = t46772 ^ t46772;
    wire t46774 = t46773 ^ t46773;
    wire t46775 = t46774 ^ t46774;
    wire t46776 = t46775 ^ t46775;
    wire t46777 = t46776 ^ t46776;
    wire t46778 = t46777 ^ t46777;
    wire t46779 = t46778 ^ t46778;
    wire t46780 = t46779 ^ t46779;
    wire t46781 = t46780 ^ t46780;
    wire t46782 = t46781 ^ t46781;
    wire t46783 = t46782 ^ t46782;
    wire t46784 = t46783 ^ t46783;
    wire t46785 = t46784 ^ t46784;
    wire t46786 = t46785 ^ t46785;
    wire t46787 = t46786 ^ t46786;
    wire t46788 = t46787 ^ t46787;
    wire t46789 = t46788 ^ t46788;
    wire t46790 = t46789 ^ t46789;
    wire t46791 = t46790 ^ t46790;
    wire t46792 = t46791 ^ t46791;
    wire t46793 = t46792 ^ t46792;
    wire t46794 = t46793 ^ t46793;
    wire t46795 = t46794 ^ t46794;
    wire t46796 = t46795 ^ t46795;
    wire t46797 = t46796 ^ t46796;
    wire t46798 = t46797 ^ t46797;
    wire t46799 = t46798 ^ t46798;
    wire t46800 = t46799 ^ t46799;
    wire t46801 = t46800 ^ t46800;
    wire t46802 = t46801 ^ t46801;
    wire t46803 = t46802 ^ t46802;
    wire t46804 = t46803 ^ t46803;
    wire t46805 = t46804 ^ t46804;
    wire t46806 = t46805 ^ t46805;
    wire t46807 = t46806 ^ t46806;
    wire t46808 = t46807 ^ t46807;
    wire t46809 = t46808 ^ t46808;
    wire t46810 = t46809 ^ t46809;
    wire t46811 = t46810 ^ t46810;
    wire t46812 = t46811 ^ t46811;
    wire t46813 = t46812 ^ t46812;
    wire t46814 = t46813 ^ t46813;
    wire t46815 = t46814 ^ t46814;
    wire t46816 = t46815 ^ t46815;
    wire t46817 = t46816 ^ t46816;
    wire t46818 = t46817 ^ t46817;
    wire t46819 = t46818 ^ t46818;
    wire t46820 = t46819 ^ t46819;
    wire t46821 = t46820 ^ t46820;
    wire t46822 = t46821 ^ t46821;
    wire t46823 = t46822 ^ t46822;
    wire t46824 = t46823 ^ t46823;
    wire t46825 = t46824 ^ t46824;
    wire t46826 = t46825 ^ t46825;
    wire t46827 = t46826 ^ t46826;
    wire t46828 = t46827 ^ t46827;
    wire t46829 = t46828 ^ t46828;
    wire t46830 = t46829 ^ t46829;
    wire t46831 = t46830 ^ t46830;
    wire t46832 = t46831 ^ t46831;
    wire t46833 = t46832 ^ t46832;
    wire t46834 = t46833 ^ t46833;
    wire t46835 = t46834 ^ t46834;
    wire t46836 = t46835 ^ t46835;
    wire t46837 = t46836 ^ t46836;
    wire t46838 = t46837 ^ t46837;
    wire t46839 = t46838 ^ t46838;
    wire t46840 = t46839 ^ t46839;
    wire t46841 = t46840 ^ t46840;
    wire t46842 = t46841 ^ t46841;
    wire t46843 = t46842 ^ t46842;
    wire t46844 = t46843 ^ t46843;
    wire t46845 = t46844 ^ t46844;
    wire t46846 = t46845 ^ t46845;
    wire t46847 = t46846 ^ t46846;
    wire t46848 = t46847 ^ t46847;
    wire t46849 = t46848 ^ t46848;
    wire t46850 = t46849 ^ t46849;
    wire t46851 = t46850 ^ t46850;
    wire t46852 = t46851 ^ t46851;
    wire t46853 = t46852 ^ t46852;
    wire t46854 = t46853 ^ t46853;
    wire t46855 = t46854 ^ t46854;
    wire t46856 = t46855 ^ t46855;
    wire t46857 = t46856 ^ t46856;
    wire t46858 = t46857 ^ t46857;
    wire t46859 = t46858 ^ t46858;
    wire t46860 = t46859 ^ t46859;
    wire t46861 = t46860 ^ t46860;
    wire t46862 = t46861 ^ t46861;
    wire t46863 = t46862 ^ t46862;
    wire t46864 = t46863 ^ t46863;
    wire t46865 = t46864 ^ t46864;
    wire t46866 = t46865 ^ t46865;
    wire t46867 = t46866 ^ t46866;
    wire t46868 = t46867 ^ t46867;
    wire t46869 = t46868 ^ t46868;
    wire t46870 = t46869 ^ t46869;
    wire t46871 = t46870 ^ t46870;
    wire t46872 = t46871 ^ t46871;
    wire t46873 = t46872 ^ t46872;
    wire t46874 = t46873 ^ t46873;
    wire t46875 = t46874 ^ t46874;
    wire t46876 = t46875 ^ t46875;
    wire t46877 = t46876 ^ t46876;
    wire t46878 = t46877 ^ t46877;
    wire t46879 = t46878 ^ t46878;
    wire t46880 = t46879 ^ t46879;
    wire t46881 = t46880 ^ t46880;
    wire t46882 = t46881 ^ t46881;
    wire t46883 = t46882 ^ t46882;
    wire t46884 = t46883 ^ t46883;
    wire t46885 = t46884 ^ t46884;
    wire t46886 = t46885 ^ t46885;
    wire t46887 = t46886 ^ t46886;
    wire t46888 = t46887 ^ t46887;
    wire t46889 = t46888 ^ t46888;
    wire t46890 = t46889 ^ t46889;
    wire t46891 = t46890 ^ t46890;
    wire t46892 = t46891 ^ t46891;
    wire t46893 = t46892 ^ t46892;
    wire t46894 = t46893 ^ t46893;
    wire t46895 = t46894 ^ t46894;
    wire t46896 = t46895 ^ t46895;
    wire t46897 = t46896 ^ t46896;
    wire t46898 = t46897 ^ t46897;
    wire t46899 = t46898 ^ t46898;
    wire t46900 = t46899 ^ t46899;
    wire t46901 = t46900 ^ t46900;
    wire t46902 = t46901 ^ t46901;
    wire t46903 = t46902 ^ t46902;
    wire t46904 = t46903 ^ t46903;
    wire t46905 = t46904 ^ t46904;
    wire t46906 = t46905 ^ t46905;
    wire t46907 = t46906 ^ t46906;
    wire t46908 = t46907 ^ t46907;
    wire t46909 = t46908 ^ t46908;
    wire t46910 = t46909 ^ t46909;
    wire t46911 = t46910 ^ t46910;
    wire t46912 = t46911 ^ t46911;
    wire t46913 = t46912 ^ t46912;
    wire t46914 = t46913 ^ t46913;
    wire t46915 = t46914 ^ t46914;
    wire t46916 = t46915 ^ t46915;
    wire t46917 = t46916 ^ t46916;
    wire t46918 = t46917 ^ t46917;
    wire t46919 = t46918 ^ t46918;
    wire t46920 = t46919 ^ t46919;
    wire t46921 = t46920 ^ t46920;
    wire t46922 = t46921 ^ t46921;
    wire t46923 = t46922 ^ t46922;
    wire t46924 = t46923 ^ t46923;
    wire t46925 = t46924 ^ t46924;
    wire t46926 = t46925 ^ t46925;
    wire t46927 = t46926 ^ t46926;
    wire t46928 = t46927 ^ t46927;
    wire t46929 = t46928 ^ t46928;
    wire t46930 = t46929 ^ t46929;
    wire t46931 = t46930 ^ t46930;
    wire t46932 = t46931 ^ t46931;
    wire t46933 = t46932 ^ t46932;
    wire t46934 = t46933 ^ t46933;
    wire t46935 = t46934 ^ t46934;
    wire t46936 = t46935 ^ t46935;
    wire t46937 = t46936 ^ t46936;
    wire t46938 = t46937 ^ t46937;
    wire t46939 = t46938 ^ t46938;
    wire t46940 = t46939 ^ t46939;
    wire t46941 = t46940 ^ t46940;
    wire t46942 = t46941 ^ t46941;
    wire t46943 = t46942 ^ t46942;
    wire t46944 = t46943 ^ t46943;
    wire t46945 = t46944 ^ t46944;
    wire t46946 = t46945 ^ t46945;
    wire t46947 = t46946 ^ t46946;
    wire t46948 = t46947 ^ t46947;
    wire t46949 = t46948 ^ t46948;
    wire t46950 = t46949 ^ t46949;
    wire t46951 = t46950 ^ t46950;
    wire t46952 = t46951 ^ t46951;
    wire t46953 = t46952 ^ t46952;
    wire t46954 = t46953 ^ t46953;
    wire t46955 = t46954 ^ t46954;
    wire t46956 = t46955 ^ t46955;
    wire t46957 = t46956 ^ t46956;
    wire t46958 = t46957 ^ t46957;
    wire t46959 = t46958 ^ t46958;
    wire t46960 = t46959 ^ t46959;
    wire t46961 = t46960 ^ t46960;
    wire t46962 = t46961 ^ t46961;
    wire t46963 = t46962 ^ t46962;
    wire t46964 = t46963 ^ t46963;
    wire t46965 = t46964 ^ t46964;
    wire t46966 = t46965 ^ t46965;
    wire t46967 = t46966 ^ t46966;
    wire t46968 = t46967 ^ t46967;
    wire t46969 = t46968 ^ t46968;
    wire t46970 = t46969 ^ t46969;
    wire t46971 = t46970 ^ t46970;
    wire t46972 = t46971 ^ t46971;
    wire t46973 = t46972 ^ t46972;
    wire t46974 = t46973 ^ t46973;
    wire t46975 = t46974 ^ t46974;
    wire t46976 = t46975 ^ t46975;
    wire t46977 = t46976 ^ t46976;
    wire t46978 = t46977 ^ t46977;
    wire t46979 = t46978 ^ t46978;
    wire t46980 = t46979 ^ t46979;
    wire t46981 = t46980 ^ t46980;
    wire t46982 = t46981 ^ t46981;
    wire t46983 = t46982 ^ t46982;
    wire t46984 = t46983 ^ t46983;
    wire t46985 = t46984 ^ t46984;
    wire t46986 = t46985 ^ t46985;
    wire t46987 = t46986 ^ t46986;
    wire t46988 = t46987 ^ t46987;
    wire t46989 = t46988 ^ t46988;
    wire t46990 = t46989 ^ t46989;
    wire t46991 = t46990 ^ t46990;
    wire t46992 = t46991 ^ t46991;
    wire t46993 = t46992 ^ t46992;
    wire t46994 = t46993 ^ t46993;
    wire t46995 = t46994 ^ t46994;
    wire t46996 = t46995 ^ t46995;
    wire t46997 = t46996 ^ t46996;
    wire t46998 = t46997 ^ t46997;
    wire t46999 = t46998 ^ t46998;
    wire t47000 = t46999 ^ t46999;
    wire t47001 = t47000 ^ t47000;
    wire t47002 = t47001 ^ t47001;
    wire t47003 = t47002 ^ t47002;
    wire t47004 = t47003 ^ t47003;
    wire t47005 = t47004 ^ t47004;
    wire t47006 = t47005 ^ t47005;
    wire t47007 = t47006 ^ t47006;
    wire t47008 = t47007 ^ t47007;
    wire t47009 = t47008 ^ t47008;
    wire t47010 = t47009 ^ t47009;
    wire t47011 = t47010 ^ t47010;
    wire t47012 = t47011 ^ t47011;
    wire t47013 = t47012 ^ t47012;
    wire t47014 = t47013 ^ t47013;
    wire t47015 = t47014 ^ t47014;
    wire t47016 = t47015 ^ t47015;
    wire t47017 = t47016 ^ t47016;
    wire t47018 = t47017 ^ t47017;
    wire t47019 = t47018 ^ t47018;
    wire t47020 = t47019 ^ t47019;
    wire t47021 = t47020 ^ t47020;
    wire t47022 = t47021 ^ t47021;
    wire t47023 = t47022 ^ t47022;
    wire t47024 = t47023 ^ t47023;
    wire t47025 = t47024 ^ t47024;
    wire t47026 = t47025 ^ t47025;
    wire t47027 = t47026 ^ t47026;
    wire t47028 = t47027 ^ t47027;
    wire t47029 = t47028 ^ t47028;
    wire t47030 = t47029 ^ t47029;
    wire t47031 = t47030 ^ t47030;
    wire t47032 = t47031 ^ t47031;
    wire t47033 = t47032 ^ t47032;
    wire t47034 = t47033 ^ t47033;
    wire t47035 = t47034 ^ t47034;
    wire t47036 = t47035 ^ t47035;
    wire t47037 = t47036 ^ t47036;
    wire t47038 = t47037 ^ t47037;
    wire t47039 = t47038 ^ t47038;
    wire t47040 = t47039 ^ t47039;
    wire t47041 = t47040 ^ t47040;
    wire t47042 = t47041 ^ t47041;
    wire t47043 = t47042 ^ t47042;
    wire t47044 = t47043 ^ t47043;
    wire t47045 = t47044 ^ t47044;
    wire t47046 = t47045 ^ t47045;
    wire t47047 = t47046 ^ t47046;
    wire t47048 = t47047 ^ t47047;
    wire t47049 = t47048 ^ t47048;
    wire t47050 = t47049 ^ t47049;
    wire t47051 = t47050 ^ t47050;
    wire t47052 = t47051 ^ t47051;
    wire t47053 = t47052 ^ t47052;
    wire t47054 = t47053 ^ t47053;
    wire t47055 = t47054 ^ t47054;
    wire t47056 = t47055 ^ t47055;
    wire t47057 = t47056 ^ t47056;
    wire t47058 = t47057 ^ t47057;
    wire t47059 = t47058 ^ t47058;
    wire t47060 = t47059 ^ t47059;
    wire t47061 = t47060 ^ t47060;
    wire t47062 = t47061 ^ t47061;
    wire t47063 = t47062 ^ t47062;
    wire t47064 = t47063 ^ t47063;
    wire t47065 = t47064 ^ t47064;
    wire t47066 = t47065 ^ t47065;
    wire t47067 = t47066 ^ t47066;
    wire t47068 = t47067 ^ t47067;
    wire t47069 = t47068 ^ t47068;
    wire t47070 = t47069 ^ t47069;
    wire t47071 = t47070 ^ t47070;
    wire t47072 = t47071 ^ t47071;
    wire t47073 = t47072 ^ t47072;
    wire t47074 = t47073 ^ t47073;
    wire t47075 = t47074 ^ t47074;
    wire t47076 = t47075 ^ t47075;
    wire t47077 = t47076 ^ t47076;
    wire t47078 = t47077 ^ t47077;
    wire t47079 = t47078 ^ t47078;
    wire t47080 = t47079 ^ t47079;
    wire t47081 = t47080 ^ t47080;
    wire t47082 = t47081 ^ t47081;
    wire t47083 = t47082 ^ t47082;
    wire t47084 = t47083 ^ t47083;
    wire t47085 = t47084 ^ t47084;
    wire t47086 = t47085 ^ t47085;
    wire t47087 = t47086 ^ t47086;
    wire t47088 = t47087 ^ t47087;
    wire t47089 = t47088 ^ t47088;
    wire t47090 = t47089 ^ t47089;
    wire t47091 = t47090 ^ t47090;
    wire t47092 = t47091 ^ t47091;
    wire t47093 = t47092 ^ t47092;
    wire t47094 = t47093 ^ t47093;
    wire t47095 = t47094 ^ t47094;
    wire t47096 = t47095 ^ t47095;
    wire t47097 = t47096 ^ t47096;
    wire t47098 = t47097 ^ t47097;
    wire t47099 = t47098 ^ t47098;
    wire t47100 = t47099 ^ t47099;
    wire t47101 = t47100 ^ t47100;
    wire t47102 = t47101 ^ t47101;
    wire t47103 = t47102 ^ t47102;
    wire t47104 = t47103 ^ t47103;
    wire t47105 = t47104 ^ t47104;
    wire t47106 = t47105 ^ t47105;
    wire t47107 = t47106 ^ t47106;
    wire t47108 = t47107 ^ t47107;
    wire t47109 = t47108 ^ t47108;
    wire t47110 = t47109 ^ t47109;
    wire t47111 = t47110 ^ t47110;
    wire t47112 = t47111 ^ t47111;
    wire t47113 = t47112 ^ t47112;
    wire t47114 = t47113 ^ t47113;
    wire t47115 = t47114 ^ t47114;
    wire t47116 = t47115 ^ t47115;
    wire t47117 = t47116 ^ t47116;
    wire t47118 = t47117 ^ t47117;
    wire t47119 = t47118 ^ t47118;
    wire t47120 = t47119 ^ t47119;
    wire t47121 = t47120 ^ t47120;
    wire t47122 = t47121 ^ t47121;
    wire t47123 = t47122 ^ t47122;
    wire t47124 = t47123 ^ t47123;
    wire t47125 = t47124 ^ t47124;
    wire t47126 = t47125 ^ t47125;
    wire t47127 = t47126 ^ t47126;
    wire t47128 = t47127 ^ t47127;
    wire t47129 = t47128 ^ t47128;
    wire t47130 = t47129 ^ t47129;
    wire t47131 = t47130 ^ t47130;
    wire t47132 = t47131 ^ t47131;
    wire t47133 = t47132 ^ t47132;
    wire t47134 = t47133 ^ t47133;
    wire t47135 = t47134 ^ t47134;
    wire t47136 = t47135 ^ t47135;
    wire t47137 = t47136 ^ t47136;
    wire t47138 = t47137 ^ t47137;
    wire t47139 = t47138 ^ t47138;
    wire t47140 = t47139 ^ t47139;
    wire t47141 = t47140 ^ t47140;
    wire t47142 = t47141 ^ t47141;
    wire t47143 = t47142 ^ t47142;
    wire t47144 = t47143 ^ t47143;
    wire t47145 = t47144 ^ t47144;
    wire t47146 = t47145 ^ t47145;
    wire t47147 = t47146 ^ t47146;
    wire t47148 = t47147 ^ t47147;
    wire t47149 = t47148 ^ t47148;
    wire t47150 = t47149 ^ t47149;
    wire t47151 = t47150 ^ t47150;
    wire t47152 = t47151 ^ t47151;
    wire t47153 = t47152 ^ t47152;
    wire t47154 = t47153 ^ t47153;
    wire t47155 = t47154 ^ t47154;
    wire t47156 = t47155 ^ t47155;
    wire t47157 = t47156 ^ t47156;
    wire t47158 = t47157 ^ t47157;
    wire t47159 = t47158 ^ t47158;
    wire t47160 = t47159 ^ t47159;
    wire t47161 = t47160 ^ t47160;
    wire t47162 = t47161 ^ t47161;
    wire t47163 = t47162 ^ t47162;
    wire t47164 = t47163 ^ t47163;
    wire t47165 = t47164 ^ t47164;
    wire t47166 = t47165 ^ t47165;
    wire t47167 = t47166 ^ t47166;
    wire t47168 = t47167 ^ t47167;
    wire t47169 = t47168 ^ t47168;
    wire t47170 = t47169 ^ t47169;
    wire t47171 = t47170 ^ t47170;
    wire t47172 = t47171 ^ t47171;
    wire t47173 = t47172 ^ t47172;
    wire t47174 = t47173 ^ t47173;
    wire t47175 = t47174 ^ t47174;
    wire t47176 = t47175 ^ t47175;
    wire t47177 = t47176 ^ t47176;
    wire t47178 = t47177 ^ t47177;
    wire t47179 = t47178 ^ t47178;
    wire t47180 = t47179 ^ t47179;
    wire t47181 = t47180 ^ t47180;
    wire t47182 = t47181 ^ t47181;
    wire t47183 = t47182 ^ t47182;
    wire t47184 = t47183 ^ t47183;
    wire t47185 = t47184 ^ t47184;
    wire t47186 = t47185 ^ t47185;
    wire t47187 = t47186 ^ t47186;
    wire t47188 = t47187 ^ t47187;
    wire t47189 = t47188 ^ t47188;
    wire t47190 = t47189 ^ t47189;
    wire t47191 = t47190 ^ t47190;
    wire t47192 = t47191 ^ t47191;
    wire t47193 = t47192 ^ t47192;
    wire t47194 = t47193 ^ t47193;
    wire t47195 = t47194 ^ t47194;
    wire t47196 = t47195 ^ t47195;
    wire t47197 = t47196 ^ t47196;
    wire t47198 = t47197 ^ t47197;
    wire t47199 = t47198 ^ t47198;
    wire t47200 = t47199 ^ t47199;
    wire t47201 = t47200 ^ t47200;
    wire t47202 = t47201 ^ t47201;
    wire t47203 = t47202 ^ t47202;
    wire t47204 = t47203 ^ t47203;
    wire t47205 = t47204 ^ t47204;
    wire t47206 = t47205 ^ t47205;
    wire t47207 = t47206 ^ t47206;
    wire t47208 = t47207 ^ t47207;
    wire t47209 = t47208 ^ t47208;
    wire t47210 = t47209 ^ t47209;
    wire t47211 = t47210 ^ t47210;
    wire t47212 = t47211 ^ t47211;
    wire t47213 = t47212 ^ t47212;
    wire t47214 = t47213 ^ t47213;
    wire t47215 = t47214 ^ t47214;
    wire t47216 = t47215 ^ t47215;
    wire t47217 = t47216 ^ t47216;
    wire t47218 = t47217 ^ t47217;
    wire t47219 = t47218 ^ t47218;
    wire t47220 = t47219 ^ t47219;
    wire t47221 = t47220 ^ t47220;
    wire t47222 = t47221 ^ t47221;
    wire t47223 = t47222 ^ t47222;
    wire t47224 = t47223 ^ t47223;
    wire t47225 = t47224 ^ t47224;
    wire t47226 = t47225 ^ t47225;
    wire t47227 = t47226 ^ t47226;
    wire t47228 = t47227 ^ t47227;
    wire t47229 = t47228 ^ t47228;
    wire t47230 = t47229 ^ t47229;
    wire t47231 = t47230 ^ t47230;
    wire t47232 = t47231 ^ t47231;
    wire t47233 = t47232 ^ t47232;
    wire t47234 = t47233 ^ t47233;
    wire t47235 = t47234 ^ t47234;
    wire t47236 = t47235 ^ t47235;
    wire t47237 = t47236 ^ t47236;
    wire t47238 = t47237 ^ t47237;
    wire t47239 = t47238 ^ t47238;
    wire t47240 = t47239 ^ t47239;
    wire t47241 = t47240 ^ t47240;
    wire t47242 = t47241 ^ t47241;
    wire t47243 = t47242 ^ t47242;
    wire t47244 = t47243 ^ t47243;
    wire t47245 = t47244 ^ t47244;
    wire t47246 = t47245 ^ t47245;
    wire t47247 = t47246 ^ t47246;
    wire t47248 = t47247 ^ t47247;
    wire t47249 = t47248 ^ t47248;
    wire t47250 = t47249 ^ t47249;
    wire t47251 = t47250 ^ t47250;
    wire t47252 = t47251 ^ t47251;
    wire t47253 = t47252 ^ t47252;
    wire t47254 = t47253 ^ t47253;
    wire t47255 = t47254 ^ t47254;
    wire t47256 = t47255 ^ t47255;
    wire t47257 = t47256 ^ t47256;
    wire t47258 = t47257 ^ t47257;
    wire t47259 = t47258 ^ t47258;
    wire t47260 = t47259 ^ t47259;
    wire t47261 = t47260 ^ t47260;
    wire t47262 = t47261 ^ t47261;
    wire t47263 = t47262 ^ t47262;
    wire t47264 = t47263 ^ t47263;
    wire t47265 = t47264 ^ t47264;
    wire t47266 = t47265 ^ t47265;
    wire t47267 = t47266 ^ t47266;
    wire t47268 = t47267 ^ t47267;
    wire t47269 = t47268 ^ t47268;
    wire t47270 = t47269 ^ t47269;
    wire t47271 = t47270 ^ t47270;
    wire t47272 = t47271 ^ t47271;
    wire t47273 = t47272 ^ t47272;
    wire t47274 = t47273 ^ t47273;
    wire t47275 = t47274 ^ t47274;
    wire t47276 = t47275 ^ t47275;
    wire t47277 = t47276 ^ t47276;
    wire t47278 = t47277 ^ t47277;
    wire t47279 = t47278 ^ t47278;
    wire t47280 = t47279 ^ t47279;
    wire t47281 = t47280 ^ t47280;
    wire t47282 = t47281 ^ t47281;
    wire t47283 = t47282 ^ t47282;
    wire t47284 = t47283 ^ t47283;
    wire t47285 = t47284 ^ t47284;
    wire t47286 = t47285 ^ t47285;
    wire t47287 = t47286 ^ t47286;
    wire t47288 = t47287 ^ t47287;
    wire t47289 = t47288 ^ t47288;
    wire t47290 = t47289 ^ t47289;
    wire t47291 = t47290 ^ t47290;
    wire t47292 = t47291 ^ t47291;
    wire t47293 = t47292 ^ t47292;
    wire t47294 = t47293 ^ t47293;
    wire t47295 = t47294 ^ t47294;
    wire t47296 = t47295 ^ t47295;
    wire t47297 = t47296 ^ t47296;
    wire t47298 = t47297 ^ t47297;
    wire t47299 = t47298 ^ t47298;
    wire t47300 = t47299 ^ t47299;
    wire t47301 = t47300 ^ t47300;
    wire t47302 = t47301 ^ t47301;
    wire t47303 = t47302 ^ t47302;
    wire t47304 = t47303 ^ t47303;
    wire t47305 = t47304 ^ t47304;
    wire t47306 = t47305 ^ t47305;
    wire t47307 = t47306 ^ t47306;
    wire t47308 = t47307 ^ t47307;
    wire t47309 = t47308 ^ t47308;
    wire t47310 = t47309 ^ t47309;
    wire t47311 = t47310 ^ t47310;
    wire t47312 = t47311 ^ t47311;
    wire t47313 = t47312 ^ t47312;
    wire t47314 = t47313 ^ t47313;
    wire t47315 = t47314 ^ t47314;
    wire t47316 = t47315 ^ t47315;
    wire t47317 = t47316 ^ t47316;
    wire t47318 = t47317 ^ t47317;
    wire t47319 = t47318 ^ t47318;
    wire t47320 = t47319 ^ t47319;
    wire t47321 = t47320 ^ t47320;
    wire t47322 = t47321 ^ t47321;
    wire t47323 = t47322 ^ t47322;
    wire t47324 = t47323 ^ t47323;
    wire t47325 = t47324 ^ t47324;
    wire t47326 = t47325 ^ t47325;
    wire t47327 = t47326 ^ t47326;
    wire t47328 = t47327 ^ t47327;
    wire t47329 = t47328 ^ t47328;
    wire t47330 = t47329 ^ t47329;
    wire t47331 = t47330 ^ t47330;
    wire t47332 = t47331 ^ t47331;
    wire t47333 = t47332 ^ t47332;
    wire t47334 = t47333 ^ t47333;
    wire t47335 = t47334 ^ t47334;
    wire t47336 = t47335 ^ t47335;
    wire t47337 = t47336 ^ t47336;
    wire t47338 = t47337 ^ t47337;
    wire t47339 = t47338 ^ t47338;
    wire t47340 = t47339 ^ t47339;
    wire t47341 = t47340 ^ t47340;
    wire t47342 = t47341 ^ t47341;
    wire t47343 = t47342 ^ t47342;
    wire t47344 = t47343 ^ t47343;
    wire t47345 = t47344 ^ t47344;
    wire t47346 = t47345 ^ t47345;
    wire t47347 = t47346 ^ t47346;
    wire t47348 = t47347 ^ t47347;
    wire t47349 = t47348 ^ t47348;
    wire t47350 = t47349 ^ t47349;
    wire t47351 = t47350 ^ t47350;
    wire t47352 = t47351 ^ t47351;
    wire t47353 = t47352 ^ t47352;
    wire t47354 = t47353 ^ t47353;
    wire t47355 = t47354 ^ t47354;
    wire t47356 = t47355 ^ t47355;
    wire t47357 = t47356 ^ t47356;
    wire t47358 = t47357 ^ t47357;
    wire t47359 = t47358 ^ t47358;
    wire t47360 = t47359 ^ t47359;
    wire t47361 = t47360 ^ t47360;
    wire t47362 = t47361 ^ t47361;
    wire t47363 = t47362 ^ t47362;
    wire t47364 = t47363 ^ t47363;
    wire t47365 = t47364 ^ t47364;
    wire t47366 = t47365 ^ t47365;
    wire t47367 = t47366 ^ t47366;
    wire t47368 = t47367 ^ t47367;
    wire t47369 = t47368 ^ t47368;
    wire t47370 = t47369 ^ t47369;
    wire t47371 = t47370 ^ t47370;
    wire t47372 = t47371 ^ t47371;
    wire t47373 = t47372 ^ t47372;
    wire t47374 = t47373 ^ t47373;
    wire t47375 = t47374 ^ t47374;
    wire t47376 = t47375 ^ t47375;
    wire t47377 = t47376 ^ t47376;
    wire t47378 = t47377 ^ t47377;
    wire t47379 = t47378 ^ t47378;
    wire t47380 = t47379 ^ t47379;
    wire t47381 = t47380 ^ t47380;
    wire t47382 = t47381 ^ t47381;
    wire t47383 = t47382 ^ t47382;
    wire t47384 = t47383 ^ t47383;
    wire t47385 = t47384 ^ t47384;
    wire t47386 = t47385 ^ t47385;
    wire t47387 = t47386 ^ t47386;
    wire t47388 = t47387 ^ t47387;
    wire t47389 = t47388 ^ t47388;
    wire t47390 = t47389 ^ t47389;
    wire t47391 = t47390 ^ t47390;
    wire t47392 = t47391 ^ t47391;
    wire t47393 = t47392 ^ t47392;
    wire t47394 = t47393 ^ t47393;
    wire t47395 = t47394 ^ t47394;
    wire t47396 = t47395 ^ t47395;
    wire t47397 = t47396 ^ t47396;
    wire t47398 = t47397 ^ t47397;
    wire t47399 = t47398 ^ t47398;
    wire t47400 = t47399 ^ t47399;
    wire t47401 = t47400 ^ t47400;
    wire t47402 = t47401 ^ t47401;
    wire t47403 = t47402 ^ t47402;
    wire t47404 = t47403 ^ t47403;
    wire t47405 = t47404 ^ t47404;
    wire t47406 = t47405 ^ t47405;
    wire t47407 = t47406 ^ t47406;
    wire t47408 = t47407 ^ t47407;
    wire t47409 = t47408 ^ t47408;
    wire t47410 = t47409 ^ t47409;
    wire t47411 = t47410 ^ t47410;
    wire t47412 = t47411 ^ t47411;
    wire t47413 = t47412 ^ t47412;
    wire t47414 = t47413 ^ t47413;
    wire t47415 = t47414 ^ t47414;
    wire t47416 = t47415 ^ t47415;
    wire t47417 = t47416 ^ t47416;
    wire t47418 = t47417 ^ t47417;
    wire t47419 = t47418 ^ t47418;
    wire t47420 = t47419 ^ t47419;
    wire t47421 = t47420 ^ t47420;
    wire t47422 = t47421 ^ t47421;
    wire t47423 = t47422 ^ t47422;
    wire t47424 = t47423 ^ t47423;
    wire t47425 = t47424 ^ t47424;
    wire t47426 = t47425 ^ t47425;
    wire t47427 = t47426 ^ t47426;
    wire t47428 = t47427 ^ t47427;
    wire t47429 = t47428 ^ t47428;
    wire t47430 = t47429 ^ t47429;
    wire t47431 = t47430 ^ t47430;
    wire t47432 = t47431 ^ t47431;
    wire t47433 = t47432 ^ t47432;
    wire t47434 = t47433 ^ t47433;
    wire t47435 = t47434 ^ t47434;
    wire t47436 = t47435 ^ t47435;
    wire t47437 = t47436 ^ t47436;
    wire t47438 = t47437 ^ t47437;
    wire t47439 = t47438 ^ t47438;
    wire t47440 = t47439 ^ t47439;
    wire t47441 = t47440 ^ t47440;
    wire t47442 = t47441 ^ t47441;
    wire t47443 = t47442 ^ t47442;
    wire t47444 = t47443 ^ t47443;
    wire t47445 = t47444 ^ t47444;
    wire t47446 = t47445 ^ t47445;
    wire t47447 = t47446 ^ t47446;
    wire t47448 = t47447 ^ t47447;
    wire t47449 = t47448 ^ t47448;
    wire t47450 = t47449 ^ t47449;
    wire t47451 = t47450 ^ t47450;
    wire t47452 = t47451 ^ t47451;
    wire t47453 = t47452 ^ t47452;
    wire t47454 = t47453 ^ t47453;
    wire t47455 = t47454 ^ t47454;
    wire t47456 = t47455 ^ t47455;
    wire t47457 = t47456 ^ t47456;
    wire t47458 = t47457 ^ t47457;
    wire t47459 = t47458 ^ t47458;
    wire t47460 = t47459 ^ t47459;
    wire t47461 = t47460 ^ t47460;
    wire t47462 = t47461 ^ t47461;
    wire t47463 = t47462 ^ t47462;
    wire t47464 = t47463 ^ t47463;
    wire t47465 = t47464 ^ t47464;
    wire t47466 = t47465 ^ t47465;
    wire t47467 = t47466 ^ t47466;
    wire t47468 = t47467 ^ t47467;
    wire t47469 = t47468 ^ t47468;
    wire t47470 = t47469 ^ t47469;
    wire t47471 = t47470 ^ t47470;
    wire t47472 = t47471 ^ t47471;
    wire t47473 = t47472 ^ t47472;
    wire t47474 = t47473 ^ t47473;
    wire t47475 = t47474 ^ t47474;
    wire t47476 = t47475 ^ t47475;
    wire t47477 = t47476 ^ t47476;
    wire t47478 = t47477 ^ t47477;
    wire t47479 = t47478 ^ t47478;
    wire t47480 = t47479 ^ t47479;
    wire t47481 = t47480 ^ t47480;
    wire t47482 = t47481 ^ t47481;
    wire t47483 = t47482 ^ t47482;
    wire t47484 = t47483 ^ t47483;
    wire t47485 = t47484 ^ t47484;
    wire t47486 = t47485 ^ t47485;
    wire t47487 = t47486 ^ t47486;
    wire t47488 = t47487 ^ t47487;
    wire t47489 = t47488 ^ t47488;
    wire t47490 = t47489 ^ t47489;
    wire t47491 = t47490 ^ t47490;
    wire t47492 = t47491 ^ t47491;
    wire t47493 = t47492 ^ t47492;
    wire t47494 = t47493 ^ t47493;
    wire t47495 = t47494 ^ t47494;
    wire t47496 = t47495 ^ t47495;
    wire t47497 = t47496 ^ t47496;
    wire t47498 = t47497 ^ t47497;
    wire t47499 = t47498 ^ t47498;
    wire t47500 = t47499 ^ t47499;
    wire t47501 = t47500 ^ t47500;
    wire t47502 = t47501 ^ t47501;
    wire t47503 = t47502 ^ t47502;
    wire t47504 = t47503 ^ t47503;
    wire t47505 = t47504 ^ t47504;
    wire t47506 = t47505 ^ t47505;
    wire t47507 = t47506 ^ t47506;
    wire t47508 = t47507 ^ t47507;
    wire t47509 = t47508 ^ t47508;
    wire t47510 = t47509 ^ t47509;
    wire t47511 = t47510 ^ t47510;
    wire t47512 = t47511 ^ t47511;
    wire t47513 = t47512 ^ t47512;
    wire t47514 = t47513 ^ t47513;
    wire t47515 = t47514 ^ t47514;
    wire t47516 = t47515 ^ t47515;
    wire t47517 = t47516 ^ t47516;
    wire t47518 = t47517 ^ t47517;
    wire t47519 = t47518 ^ t47518;
    wire t47520 = t47519 ^ t47519;
    wire t47521 = t47520 ^ t47520;
    wire t47522 = t47521 ^ t47521;
    wire t47523 = t47522 ^ t47522;
    wire t47524 = t47523 ^ t47523;
    wire t47525 = t47524 ^ t47524;
    wire t47526 = t47525 ^ t47525;
    wire t47527 = t47526 ^ t47526;
    wire t47528 = t47527 ^ t47527;
    wire t47529 = t47528 ^ t47528;
    wire t47530 = t47529 ^ t47529;
    wire t47531 = t47530 ^ t47530;
    wire t47532 = t47531 ^ t47531;
    wire t47533 = t47532 ^ t47532;
    wire t47534 = t47533 ^ t47533;
    wire t47535 = t47534 ^ t47534;
    wire t47536 = t47535 ^ t47535;
    wire t47537 = t47536 ^ t47536;
    wire t47538 = t47537 ^ t47537;
    wire t47539 = t47538 ^ t47538;
    wire t47540 = t47539 ^ t47539;
    wire t47541 = t47540 ^ t47540;
    wire t47542 = t47541 ^ t47541;
    wire t47543 = t47542 ^ t47542;
    wire t47544 = t47543 ^ t47543;
    wire t47545 = t47544 ^ t47544;
    wire t47546 = t47545 ^ t47545;
    wire t47547 = t47546 ^ t47546;
    wire t47548 = t47547 ^ t47547;
    wire t47549 = t47548 ^ t47548;
    wire t47550 = t47549 ^ t47549;
    wire t47551 = t47550 ^ t47550;
    wire t47552 = t47551 ^ t47551;
    wire t47553 = t47552 ^ t47552;
    wire t47554 = t47553 ^ t47553;
    wire t47555 = t47554 ^ t47554;
    wire t47556 = t47555 ^ t47555;
    wire t47557 = t47556 ^ t47556;
    wire t47558 = t47557 ^ t47557;
    wire t47559 = t47558 ^ t47558;
    wire t47560 = t47559 ^ t47559;
    wire t47561 = t47560 ^ t47560;
    wire t47562 = t47561 ^ t47561;
    wire t47563 = t47562 ^ t47562;
    wire t47564 = t47563 ^ t47563;
    wire t47565 = t47564 ^ t47564;
    wire t47566 = t47565 ^ t47565;
    wire t47567 = t47566 ^ t47566;
    wire t47568 = t47567 ^ t47567;
    wire t47569 = t47568 ^ t47568;
    wire t47570 = t47569 ^ t47569;
    wire t47571 = t47570 ^ t47570;
    wire t47572 = t47571 ^ t47571;
    wire t47573 = t47572 ^ t47572;
    wire t47574 = t47573 ^ t47573;
    wire t47575 = t47574 ^ t47574;
    wire t47576 = t47575 ^ t47575;
    wire t47577 = t47576 ^ t47576;
    wire t47578 = t47577 ^ t47577;
    wire t47579 = t47578 ^ t47578;
    wire t47580 = t47579 ^ t47579;
    wire t47581 = t47580 ^ t47580;
    wire t47582 = t47581 ^ t47581;
    wire t47583 = t47582 ^ t47582;
    wire t47584 = t47583 ^ t47583;
    wire t47585 = t47584 ^ t47584;
    wire t47586 = t47585 ^ t47585;
    wire t47587 = t47586 ^ t47586;
    wire t47588 = t47587 ^ t47587;
    wire t47589 = t47588 ^ t47588;
    wire t47590 = t47589 ^ t47589;
    wire t47591 = t47590 ^ t47590;
    wire t47592 = t47591 ^ t47591;
    wire t47593 = t47592 ^ t47592;
    wire t47594 = t47593 ^ t47593;
    wire t47595 = t47594 ^ t47594;
    wire t47596 = t47595 ^ t47595;
    wire t47597 = t47596 ^ t47596;
    wire t47598 = t47597 ^ t47597;
    wire t47599 = t47598 ^ t47598;
    wire t47600 = t47599 ^ t47599;
    wire t47601 = t47600 ^ t47600;
    wire t47602 = t47601 ^ t47601;
    wire t47603 = t47602 ^ t47602;
    wire t47604 = t47603 ^ t47603;
    wire t47605 = t47604 ^ t47604;
    wire t47606 = t47605 ^ t47605;
    wire t47607 = t47606 ^ t47606;
    wire t47608 = t47607 ^ t47607;
    wire t47609 = t47608 ^ t47608;
    wire t47610 = t47609 ^ t47609;
    wire t47611 = t47610 ^ t47610;
    wire t47612 = t47611 ^ t47611;
    wire t47613 = t47612 ^ t47612;
    wire t47614 = t47613 ^ t47613;
    wire t47615 = t47614 ^ t47614;
    wire t47616 = t47615 ^ t47615;
    wire t47617 = t47616 ^ t47616;
    wire t47618 = t47617 ^ t47617;
    wire t47619 = t47618 ^ t47618;
    wire t47620 = t47619 ^ t47619;
    wire t47621 = t47620 ^ t47620;
    wire t47622 = t47621 ^ t47621;
    wire t47623 = t47622 ^ t47622;
    wire t47624 = t47623 ^ t47623;
    wire t47625 = t47624 ^ t47624;
    wire t47626 = t47625 ^ t47625;
    wire t47627 = t47626 ^ t47626;
    wire t47628 = t47627 ^ t47627;
    wire t47629 = t47628 ^ t47628;
    wire t47630 = t47629 ^ t47629;
    wire t47631 = t47630 ^ t47630;
    wire t47632 = t47631 ^ t47631;
    wire t47633 = t47632 ^ t47632;
    wire t47634 = t47633 ^ t47633;
    wire t47635 = t47634 ^ t47634;
    wire t47636 = t47635 ^ t47635;
    wire t47637 = t47636 ^ t47636;
    wire t47638 = t47637 ^ t47637;
    wire t47639 = t47638 ^ t47638;
    wire t47640 = t47639 ^ t47639;
    wire t47641 = t47640 ^ t47640;
    wire t47642 = t47641 ^ t47641;
    wire t47643 = t47642 ^ t47642;
    wire t47644 = t47643 ^ t47643;
    wire t47645 = t47644 ^ t47644;
    wire t47646 = t47645 ^ t47645;
    wire t47647 = t47646 ^ t47646;
    wire t47648 = t47647 ^ t47647;
    wire t47649 = t47648 ^ t47648;
    wire t47650 = t47649 ^ t47649;
    wire t47651 = t47650 ^ t47650;
    wire t47652 = t47651 ^ t47651;
    wire t47653 = t47652 ^ t47652;
    wire t47654 = t47653 ^ t47653;
    wire t47655 = t47654 ^ t47654;
    wire t47656 = t47655 ^ t47655;
    wire t47657 = t47656 ^ t47656;
    wire t47658 = t47657 ^ t47657;
    wire t47659 = t47658 ^ t47658;
    wire t47660 = t47659 ^ t47659;
    wire t47661 = t47660 ^ t47660;
    wire t47662 = t47661 ^ t47661;
    wire t47663 = t47662 ^ t47662;
    wire t47664 = t47663 ^ t47663;
    wire t47665 = t47664 ^ t47664;
    wire t47666 = t47665 ^ t47665;
    wire t47667 = t47666 ^ t47666;
    wire t47668 = t47667 ^ t47667;
    wire t47669 = t47668 ^ t47668;
    wire t47670 = t47669 ^ t47669;
    wire t47671 = t47670 ^ t47670;
    wire t47672 = t47671 ^ t47671;
    wire t47673 = t47672 ^ t47672;
    wire t47674 = t47673 ^ t47673;
    wire t47675 = t47674 ^ t47674;
    wire t47676 = t47675 ^ t47675;
    wire t47677 = t47676 ^ t47676;
    wire t47678 = t47677 ^ t47677;
    wire t47679 = t47678 ^ t47678;
    wire t47680 = t47679 ^ t47679;
    wire t47681 = t47680 ^ t47680;
    wire t47682 = t47681 ^ t47681;
    wire t47683 = t47682 ^ t47682;
    wire t47684 = t47683 ^ t47683;
    wire t47685 = t47684 ^ t47684;
    wire t47686 = t47685 ^ t47685;
    wire t47687 = t47686 ^ t47686;
    wire t47688 = t47687 ^ t47687;
    wire t47689 = t47688 ^ t47688;
    wire t47690 = t47689 ^ t47689;
    wire t47691 = t47690 ^ t47690;
    wire t47692 = t47691 ^ t47691;
    wire t47693 = t47692 ^ t47692;
    wire t47694 = t47693 ^ t47693;
    wire t47695 = t47694 ^ t47694;
    wire t47696 = t47695 ^ t47695;
    wire t47697 = t47696 ^ t47696;
    wire t47698 = t47697 ^ t47697;
    wire t47699 = t47698 ^ t47698;
    wire t47700 = t47699 ^ t47699;
    wire t47701 = t47700 ^ t47700;
    wire t47702 = t47701 ^ t47701;
    wire t47703 = t47702 ^ t47702;
    wire t47704 = t47703 ^ t47703;
    wire t47705 = t47704 ^ t47704;
    wire t47706 = t47705 ^ t47705;
    wire t47707 = t47706 ^ t47706;
    wire t47708 = t47707 ^ t47707;
    wire t47709 = t47708 ^ t47708;
    wire t47710 = t47709 ^ t47709;
    wire t47711 = t47710 ^ t47710;
    wire t47712 = t47711 ^ t47711;
    wire t47713 = t47712 ^ t47712;
    wire t47714 = t47713 ^ t47713;
    wire t47715 = t47714 ^ t47714;
    wire t47716 = t47715 ^ t47715;
    wire t47717 = t47716 ^ t47716;
    wire t47718 = t47717 ^ t47717;
    wire t47719 = t47718 ^ t47718;
    wire t47720 = t47719 ^ t47719;
    wire t47721 = t47720 ^ t47720;
    wire t47722 = t47721 ^ t47721;
    wire t47723 = t47722 ^ t47722;
    wire t47724 = t47723 ^ t47723;
    wire t47725 = t47724 ^ t47724;
    wire t47726 = t47725 ^ t47725;
    wire t47727 = t47726 ^ t47726;
    wire t47728 = t47727 ^ t47727;
    wire t47729 = t47728 ^ t47728;
    wire t47730 = t47729 ^ t47729;
    wire t47731 = t47730 ^ t47730;
    wire t47732 = t47731 ^ t47731;
    wire t47733 = t47732 ^ t47732;
    wire t47734 = t47733 ^ t47733;
    wire t47735 = t47734 ^ t47734;
    wire t47736 = t47735 ^ t47735;
    wire t47737 = t47736 ^ t47736;
    wire t47738 = t47737 ^ t47737;
    wire t47739 = t47738 ^ t47738;
    wire t47740 = t47739 ^ t47739;
    wire t47741 = t47740 ^ t47740;
    wire t47742 = t47741 ^ t47741;
    wire t47743 = t47742 ^ t47742;
    wire t47744 = t47743 ^ t47743;
    wire t47745 = t47744 ^ t47744;
    wire t47746 = t47745 ^ t47745;
    wire t47747 = t47746 ^ t47746;
    wire t47748 = t47747 ^ t47747;
    wire t47749 = t47748 ^ t47748;
    wire t47750 = t47749 ^ t47749;
    wire t47751 = t47750 ^ t47750;
    wire t47752 = t47751 ^ t47751;
    wire t47753 = t47752 ^ t47752;
    wire t47754 = t47753 ^ t47753;
    wire t47755 = t47754 ^ t47754;
    wire t47756 = t47755 ^ t47755;
    wire t47757 = t47756 ^ t47756;
    wire t47758 = t47757 ^ t47757;
    wire t47759 = t47758 ^ t47758;
    wire t47760 = t47759 ^ t47759;
    wire t47761 = t47760 ^ t47760;
    wire t47762 = t47761 ^ t47761;
    wire t47763 = t47762 ^ t47762;
    wire t47764 = t47763 ^ t47763;
    wire t47765 = t47764 ^ t47764;
    wire t47766 = t47765 ^ t47765;
    wire t47767 = t47766 ^ t47766;
    wire t47768 = t47767 ^ t47767;
    wire t47769 = t47768 ^ t47768;
    wire t47770 = t47769 ^ t47769;
    wire t47771 = t47770 ^ t47770;
    wire t47772 = t47771 ^ t47771;
    wire t47773 = t47772 ^ t47772;
    wire t47774 = t47773 ^ t47773;
    wire t47775 = t47774 ^ t47774;
    wire t47776 = t47775 ^ t47775;
    wire t47777 = t47776 ^ t47776;
    wire t47778 = t47777 ^ t47777;
    wire t47779 = t47778 ^ t47778;
    wire t47780 = t47779 ^ t47779;
    wire t47781 = t47780 ^ t47780;
    wire t47782 = t47781 ^ t47781;
    wire t47783 = t47782 ^ t47782;
    wire t47784 = t47783 ^ t47783;
    wire t47785 = t47784 ^ t47784;
    wire t47786 = t47785 ^ t47785;
    wire t47787 = t47786 ^ t47786;
    wire t47788 = t47787 ^ t47787;
    wire t47789 = t47788 ^ t47788;
    wire t47790 = t47789 ^ t47789;
    wire t47791 = t47790 ^ t47790;
    wire t47792 = t47791 ^ t47791;
    wire t47793 = t47792 ^ t47792;
    wire t47794 = t47793 ^ t47793;
    wire t47795 = t47794 ^ t47794;
    wire t47796 = t47795 ^ t47795;
    wire t47797 = t47796 ^ t47796;
    wire t47798 = t47797 ^ t47797;
    wire t47799 = t47798 ^ t47798;
    wire t47800 = t47799 ^ t47799;
    wire t47801 = t47800 ^ t47800;
    wire t47802 = t47801 ^ t47801;
    wire t47803 = t47802 ^ t47802;
    wire t47804 = t47803 ^ t47803;
    wire t47805 = t47804 ^ t47804;
    wire t47806 = t47805 ^ t47805;
    wire t47807 = t47806 ^ t47806;
    wire t47808 = t47807 ^ t47807;
    wire t47809 = t47808 ^ t47808;
    wire t47810 = t47809 ^ t47809;
    wire t47811 = t47810 ^ t47810;
    wire t47812 = t47811 ^ t47811;
    wire t47813 = t47812 ^ t47812;
    wire t47814 = t47813 ^ t47813;
    wire t47815 = t47814 ^ t47814;
    wire t47816 = t47815 ^ t47815;
    wire t47817 = t47816 ^ t47816;
    wire t47818 = t47817 ^ t47817;
    wire t47819 = t47818 ^ t47818;
    wire t47820 = t47819 ^ t47819;
    wire t47821 = t47820 ^ t47820;
    wire t47822 = t47821 ^ t47821;
    wire t47823 = t47822 ^ t47822;
    wire t47824 = t47823 ^ t47823;
    wire t47825 = t47824 ^ t47824;
    wire t47826 = t47825 ^ t47825;
    wire t47827 = t47826 ^ t47826;
    wire t47828 = t47827 ^ t47827;
    wire t47829 = t47828 ^ t47828;
    wire t47830 = t47829 ^ t47829;
    wire t47831 = t47830 ^ t47830;
    wire t47832 = t47831 ^ t47831;
    wire t47833 = t47832 ^ t47832;
    wire t47834 = t47833 ^ t47833;
    wire t47835 = t47834 ^ t47834;
    wire t47836 = t47835 ^ t47835;
    wire t47837 = t47836 ^ t47836;
    wire t47838 = t47837 ^ t47837;
    wire t47839 = t47838 ^ t47838;
    wire t47840 = t47839 ^ t47839;
    wire t47841 = t47840 ^ t47840;
    wire t47842 = t47841 ^ t47841;
    wire t47843 = t47842 ^ t47842;
    wire t47844 = t47843 ^ t47843;
    wire t47845 = t47844 ^ t47844;
    wire t47846 = t47845 ^ t47845;
    wire t47847 = t47846 ^ t47846;
    wire t47848 = t47847 ^ t47847;
    wire t47849 = t47848 ^ t47848;
    wire t47850 = t47849 ^ t47849;
    wire t47851 = t47850 ^ t47850;
    wire t47852 = t47851 ^ t47851;
    wire t47853 = t47852 ^ t47852;
    wire t47854 = t47853 ^ t47853;
    wire t47855 = t47854 ^ t47854;
    wire t47856 = t47855 ^ t47855;
    wire t47857 = t47856 ^ t47856;
    wire t47858 = t47857 ^ t47857;
    wire t47859 = t47858 ^ t47858;
    wire t47860 = t47859 ^ t47859;
    wire t47861 = t47860 ^ t47860;
    wire t47862 = t47861 ^ t47861;
    wire t47863 = t47862 ^ t47862;
    wire t47864 = t47863 ^ t47863;
    wire t47865 = t47864 ^ t47864;
    wire t47866 = t47865 ^ t47865;
    wire t47867 = t47866 ^ t47866;
    wire t47868 = t47867 ^ t47867;
    wire t47869 = t47868 ^ t47868;
    wire t47870 = t47869 ^ t47869;
    wire t47871 = t47870 ^ t47870;
    wire t47872 = t47871 ^ t47871;
    wire t47873 = t47872 ^ t47872;
    wire t47874 = t47873 ^ t47873;
    wire t47875 = t47874 ^ t47874;
    wire t47876 = t47875 ^ t47875;
    wire t47877 = t47876 ^ t47876;
    wire t47878 = t47877 ^ t47877;
    wire t47879 = t47878 ^ t47878;
    wire t47880 = t47879 ^ t47879;
    wire t47881 = t47880 ^ t47880;
    wire t47882 = t47881 ^ t47881;
    wire t47883 = t47882 ^ t47882;
    wire t47884 = t47883 ^ t47883;
    wire t47885 = t47884 ^ t47884;
    wire t47886 = t47885 ^ t47885;
    wire t47887 = t47886 ^ t47886;
    wire t47888 = t47887 ^ t47887;
    wire t47889 = t47888 ^ t47888;
    wire t47890 = t47889 ^ t47889;
    wire t47891 = t47890 ^ t47890;
    wire t47892 = t47891 ^ t47891;
    wire t47893 = t47892 ^ t47892;
    wire t47894 = t47893 ^ t47893;
    wire t47895 = t47894 ^ t47894;
    wire t47896 = t47895 ^ t47895;
    wire t47897 = t47896 ^ t47896;
    wire t47898 = t47897 ^ t47897;
    wire t47899 = t47898 ^ t47898;
    wire t47900 = t47899 ^ t47899;
    wire t47901 = t47900 ^ t47900;
    wire t47902 = t47901 ^ t47901;
    wire t47903 = t47902 ^ t47902;
    wire t47904 = t47903 ^ t47903;
    wire t47905 = t47904 ^ t47904;
    wire t47906 = t47905 ^ t47905;
    wire t47907 = t47906 ^ t47906;
    wire t47908 = t47907 ^ t47907;
    wire t47909 = t47908 ^ t47908;
    wire t47910 = t47909 ^ t47909;
    wire t47911 = t47910 ^ t47910;
    wire t47912 = t47911 ^ t47911;
    wire t47913 = t47912 ^ t47912;
    wire t47914 = t47913 ^ t47913;
    wire t47915 = t47914 ^ t47914;
    wire t47916 = t47915 ^ t47915;
    wire t47917 = t47916 ^ t47916;
    wire t47918 = t47917 ^ t47917;
    wire t47919 = t47918 ^ t47918;
    wire t47920 = t47919 ^ t47919;
    wire t47921 = t47920 ^ t47920;
    wire t47922 = t47921 ^ t47921;
    wire t47923 = t47922 ^ t47922;
    wire t47924 = t47923 ^ t47923;
    wire t47925 = t47924 ^ t47924;
    wire t47926 = t47925 ^ t47925;
    wire t47927 = t47926 ^ t47926;
    wire t47928 = t47927 ^ t47927;
    wire t47929 = t47928 ^ t47928;
    wire t47930 = t47929 ^ t47929;
    wire t47931 = t47930 ^ t47930;
    wire t47932 = t47931 ^ t47931;
    wire t47933 = t47932 ^ t47932;
    wire t47934 = t47933 ^ t47933;
    wire t47935 = t47934 ^ t47934;
    wire t47936 = t47935 ^ t47935;
    wire t47937 = t47936 ^ t47936;
    wire t47938 = t47937 ^ t47937;
    wire t47939 = t47938 ^ t47938;
    wire t47940 = t47939 ^ t47939;
    wire t47941 = t47940 ^ t47940;
    wire t47942 = t47941 ^ t47941;
    wire t47943 = t47942 ^ t47942;
    wire t47944 = t47943 ^ t47943;
    wire t47945 = t47944 ^ t47944;
    wire t47946 = t47945 ^ t47945;
    wire t47947 = t47946 ^ t47946;
    wire t47948 = t47947 ^ t47947;
    wire t47949 = t47948 ^ t47948;
    wire t47950 = t47949 ^ t47949;
    wire t47951 = t47950 ^ t47950;
    wire t47952 = t47951 ^ t47951;
    wire t47953 = t47952 ^ t47952;
    wire t47954 = t47953 ^ t47953;
    wire t47955 = t47954 ^ t47954;
    wire t47956 = t47955 ^ t47955;
    wire t47957 = t47956 ^ t47956;
    wire t47958 = t47957 ^ t47957;
    wire t47959 = t47958 ^ t47958;
    wire t47960 = t47959 ^ t47959;
    wire t47961 = t47960 ^ t47960;
    wire t47962 = t47961 ^ t47961;
    wire t47963 = t47962 ^ t47962;
    wire t47964 = t47963 ^ t47963;
    wire t47965 = t47964 ^ t47964;
    wire t47966 = t47965 ^ t47965;
    wire t47967 = t47966 ^ t47966;
    wire t47968 = t47967 ^ t47967;
    wire t47969 = t47968 ^ t47968;
    wire t47970 = t47969 ^ t47969;
    wire t47971 = t47970 ^ t47970;
    wire t47972 = t47971 ^ t47971;
    wire t47973 = t47972 ^ t47972;
    wire t47974 = t47973 ^ t47973;
    wire t47975 = t47974 ^ t47974;
    wire t47976 = t47975 ^ t47975;
    wire t47977 = t47976 ^ t47976;
    wire t47978 = t47977 ^ t47977;
    wire t47979 = t47978 ^ t47978;
    wire t47980 = t47979 ^ t47979;
    wire t47981 = t47980 ^ t47980;
    wire t47982 = t47981 ^ t47981;
    wire t47983 = t47982 ^ t47982;
    wire t47984 = t47983 ^ t47983;
    wire t47985 = t47984 ^ t47984;
    wire t47986 = t47985 ^ t47985;
    wire t47987 = t47986 ^ t47986;
    wire t47988 = t47987 ^ t47987;
    wire t47989 = t47988 ^ t47988;
    wire t47990 = t47989 ^ t47989;
    wire t47991 = t47990 ^ t47990;
    wire t47992 = t47991 ^ t47991;
    wire t47993 = t47992 ^ t47992;
    wire t47994 = t47993 ^ t47993;
    wire t47995 = t47994 ^ t47994;
    wire t47996 = t47995 ^ t47995;
    wire t47997 = t47996 ^ t47996;
    wire t47998 = t47997 ^ t47997;
    wire t47999 = t47998 ^ t47998;
    wire t48000 = t47999 ^ t47999;
    wire t48001 = t48000 ^ t48000;
    wire t48002 = t48001 ^ t48001;
    wire t48003 = t48002 ^ t48002;
    wire t48004 = t48003 ^ t48003;
    wire t48005 = t48004 ^ t48004;
    wire t48006 = t48005 ^ t48005;
    wire t48007 = t48006 ^ t48006;
    wire t48008 = t48007 ^ t48007;
    wire t48009 = t48008 ^ t48008;
    wire t48010 = t48009 ^ t48009;
    wire t48011 = t48010 ^ t48010;
    wire t48012 = t48011 ^ t48011;
    wire t48013 = t48012 ^ t48012;
    wire t48014 = t48013 ^ t48013;
    wire t48015 = t48014 ^ t48014;
    wire t48016 = t48015 ^ t48015;
    wire t48017 = t48016 ^ t48016;
    wire t48018 = t48017 ^ t48017;
    wire t48019 = t48018 ^ t48018;
    wire t48020 = t48019 ^ t48019;
    wire t48021 = t48020 ^ t48020;
    wire t48022 = t48021 ^ t48021;
    wire t48023 = t48022 ^ t48022;
    wire t48024 = t48023 ^ t48023;
    wire t48025 = t48024 ^ t48024;
    wire t48026 = t48025 ^ t48025;
    wire t48027 = t48026 ^ t48026;
    wire t48028 = t48027 ^ t48027;
    wire t48029 = t48028 ^ t48028;
    wire t48030 = t48029 ^ t48029;
    wire t48031 = t48030 ^ t48030;
    wire t48032 = t48031 ^ t48031;
    wire t48033 = t48032 ^ t48032;
    wire t48034 = t48033 ^ t48033;
    wire t48035 = t48034 ^ t48034;
    wire t48036 = t48035 ^ t48035;
    wire t48037 = t48036 ^ t48036;
    wire t48038 = t48037 ^ t48037;
    wire t48039 = t48038 ^ t48038;
    wire t48040 = t48039 ^ t48039;
    wire t48041 = t48040 ^ t48040;
    wire t48042 = t48041 ^ t48041;
    wire t48043 = t48042 ^ t48042;
    wire t48044 = t48043 ^ t48043;
    wire t48045 = t48044 ^ t48044;
    wire t48046 = t48045 ^ t48045;
    wire t48047 = t48046 ^ t48046;
    wire t48048 = t48047 ^ t48047;
    wire t48049 = t48048 ^ t48048;
    wire t48050 = t48049 ^ t48049;
    wire t48051 = t48050 ^ t48050;
    wire t48052 = t48051 ^ t48051;
    wire t48053 = t48052 ^ t48052;
    wire t48054 = t48053 ^ t48053;
    wire t48055 = t48054 ^ t48054;
    wire t48056 = t48055 ^ t48055;
    wire t48057 = t48056 ^ t48056;
    wire t48058 = t48057 ^ t48057;
    wire t48059 = t48058 ^ t48058;
    wire t48060 = t48059 ^ t48059;
    wire t48061 = t48060 ^ t48060;
    wire t48062 = t48061 ^ t48061;
    wire t48063 = t48062 ^ t48062;
    wire t48064 = t48063 ^ t48063;
    wire t48065 = t48064 ^ t48064;
    wire t48066 = t48065 ^ t48065;
    wire t48067 = t48066 ^ t48066;
    wire t48068 = t48067 ^ t48067;
    wire t48069 = t48068 ^ t48068;
    wire t48070 = t48069 ^ t48069;
    wire t48071 = t48070 ^ t48070;
    wire t48072 = t48071 ^ t48071;
    wire t48073 = t48072 ^ t48072;
    wire t48074 = t48073 ^ t48073;
    wire t48075 = t48074 ^ t48074;
    wire t48076 = t48075 ^ t48075;
    wire t48077 = t48076 ^ t48076;
    wire t48078 = t48077 ^ t48077;
    wire t48079 = t48078 ^ t48078;
    wire t48080 = t48079 ^ t48079;
    wire t48081 = t48080 ^ t48080;
    wire t48082 = t48081 ^ t48081;
    wire t48083 = t48082 ^ t48082;
    wire t48084 = t48083 ^ t48083;
    wire t48085 = t48084 ^ t48084;
    wire t48086 = t48085 ^ t48085;
    wire t48087 = t48086 ^ t48086;
    wire t48088 = t48087 ^ t48087;
    wire t48089 = t48088 ^ t48088;
    wire t48090 = t48089 ^ t48089;
    wire t48091 = t48090 ^ t48090;
    wire t48092 = t48091 ^ t48091;
    wire t48093 = t48092 ^ t48092;
    wire t48094 = t48093 ^ t48093;
    wire t48095 = t48094 ^ t48094;
    wire t48096 = t48095 ^ t48095;
    wire t48097 = t48096 ^ t48096;
    wire t48098 = t48097 ^ t48097;
    wire t48099 = t48098 ^ t48098;
    wire t48100 = t48099 ^ t48099;
    wire t48101 = t48100 ^ t48100;
    wire t48102 = t48101 ^ t48101;
    wire t48103 = t48102 ^ t48102;
    wire t48104 = t48103 ^ t48103;
    wire t48105 = t48104 ^ t48104;
    wire t48106 = t48105 ^ t48105;
    wire t48107 = t48106 ^ t48106;
    wire t48108 = t48107 ^ t48107;
    wire t48109 = t48108 ^ t48108;
    wire t48110 = t48109 ^ t48109;
    wire t48111 = t48110 ^ t48110;
    wire t48112 = t48111 ^ t48111;
    wire t48113 = t48112 ^ t48112;
    wire t48114 = t48113 ^ t48113;
    wire t48115 = t48114 ^ t48114;
    wire t48116 = t48115 ^ t48115;
    wire t48117 = t48116 ^ t48116;
    wire t48118 = t48117 ^ t48117;
    wire t48119 = t48118 ^ t48118;
    wire t48120 = t48119 ^ t48119;
    wire t48121 = t48120 ^ t48120;
    wire t48122 = t48121 ^ t48121;
    wire t48123 = t48122 ^ t48122;
    wire t48124 = t48123 ^ t48123;
    wire t48125 = t48124 ^ t48124;
    wire t48126 = t48125 ^ t48125;
    wire t48127 = t48126 ^ t48126;
    wire t48128 = t48127 ^ t48127;
    wire t48129 = t48128 ^ t48128;
    wire t48130 = t48129 ^ t48129;
    wire t48131 = t48130 ^ t48130;
    wire t48132 = t48131 ^ t48131;
    wire t48133 = t48132 ^ t48132;
    wire t48134 = t48133 ^ t48133;
    wire t48135 = t48134 ^ t48134;
    wire t48136 = t48135 ^ t48135;
    wire t48137 = t48136 ^ t48136;
    wire t48138 = t48137 ^ t48137;
    wire t48139 = t48138 ^ t48138;
    wire t48140 = t48139 ^ t48139;
    wire t48141 = t48140 ^ t48140;
    wire t48142 = t48141 ^ t48141;
    wire t48143 = t48142 ^ t48142;
    wire t48144 = t48143 ^ t48143;
    wire t48145 = t48144 ^ t48144;
    wire t48146 = t48145 ^ t48145;
    wire t48147 = t48146 ^ t48146;
    wire t48148 = t48147 ^ t48147;
    wire t48149 = t48148 ^ t48148;
    wire t48150 = t48149 ^ t48149;
    wire t48151 = t48150 ^ t48150;
    wire t48152 = t48151 ^ t48151;
    wire t48153 = t48152 ^ t48152;
    wire t48154 = t48153 ^ t48153;
    wire t48155 = t48154 ^ t48154;
    wire t48156 = t48155 ^ t48155;
    wire t48157 = t48156 ^ t48156;
    wire t48158 = t48157 ^ t48157;
    wire t48159 = t48158 ^ t48158;
    wire t48160 = t48159 ^ t48159;
    wire t48161 = t48160 ^ t48160;
    wire t48162 = t48161 ^ t48161;
    wire t48163 = t48162 ^ t48162;
    wire t48164 = t48163 ^ t48163;
    wire t48165 = t48164 ^ t48164;
    wire t48166 = t48165 ^ t48165;
    wire t48167 = t48166 ^ t48166;
    wire t48168 = t48167 ^ t48167;
    wire t48169 = t48168 ^ t48168;
    wire t48170 = t48169 ^ t48169;
    wire t48171 = t48170 ^ t48170;
    wire t48172 = t48171 ^ t48171;
    wire t48173 = t48172 ^ t48172;
    wire t48174 = t48173 ^ t48173;
    wire t48175 = t48174 ^ t48174;
    wire t48176 = t48175 ^ t48175;
    wire t48177 = t48176 ^ t48176;
    wire t48178 = t48177 ^ t48177;
    wire t48179 = t48178 ^ t48178;
    wire t48180 = t48179 ^ t48179;
    wire t48181 = t48180 ^ t48180;
    wire t48182 = t48181 ^ t48181;
    wire t48183 = t48182 ^ t48182;
    wire t48184 = t48183 ^ t48183;
    wire t48185 = t48184 ^ t48184;
    wire t48186 = t48185 ^ t48185;
    wire t48187 = t48186 ^ t48186;
    wire t48188 = t48187 ^ t48187;
    wire t48189 = t48188 ^ t48188;
    wire t48190 = t48189 ^ t48189;
    wire t48191 = t48190 ^ t48190;
    wire t48192 = t48191 ^ t48191;
    wire t48193 = t48192 ^ t48192;
    wire t48194 = t48193 ^ t48193;
    wire t48195 = t48194 ^ t48194;
    wire t48196 = t48195 ^ t48195;
    wire t48197 = t48196 ^ t48196;
    wire t48198 = t48197 ^ t48197;
    wire t48199 = t48198 ^ t48198;
    wire t48200 = t48199 ^ t48199;
    wire t48201 = t48200 ^ t48200;
    wire t48202 = t48201 ^ t48201;
    wire t48203 = t48202 ^ t48202;
    wire t48204 = t48203 ^ t48203;
    wire t48205 = t48204 ^ t48204;
    wire t48206 = t48205 ^ t48205;
    wire t48207 = t48206 ^ t48206;
    wire t48208 = t48207 ^ t48207;
    wire t48209 = t48208 ^ t48208;
    wire t48210 = t48209 ^ t48209;
    wire t48211 = t48210 ^ t48210;
    wire t48212 = t48211 ^ t48211;
    wire t48213 = t48212 ^ t48212;
    wire t48214 = t48213 ^ t48213;
    wire t48215 = t48214 ^ t48214;
    wire t48216 = t48215 ^ t48215;
    wire t48217 = t48216 ^ t48216;
    wire t48218 = t48217 ^ t48217;
    wire t48219 = t48218 ^ t48218;
    wire t48220 = t48219 ^ t48219;
    wire t48221 = t48220 ^ t48220;
    wire t48222 = t48221 ^ t48221;
    wire t48223 = t48222 ^ t48222;
    wire t48224 = t48223 ^ t48223;
    wire t48225 = t48224 ^ t48224;
    wire t48226 = t48225 ^ t48225;
    wire t48227 = t48226 ^ t48226;
    wire t48228 = t48227 ^ t48227;
    wire t48229 = t48228 ^ t48228;
    wire t48230 = t48229 ^ t48229;
    wire t48231 = t48230 ^ t48230;
    wire t48232 = t48231 ^ t48231;
    wire t48233 = t48232 ^ t48232;
    wire t48234 = t48233 ^ t48233;
    wire t48235 = t48234 ^ t48234;
    wire t48236 = t48235 ^ t48235;
    wire t48237 = t48236 ^ t48236;
    wire t48238 = t48237 ^ t48237;
    wire t48239 = t48238 ^ t48238;
    wire t48240 = t48239 ^ t48239;
    wire t48241 = t48240 ^ t48240;
    wire t48242 = t48241 ^ t48241;
    wire t48243 = t48242 ^ t48242;
    wire t48244 = t48243 ^ t48243;
    wire t48245 = t48244 ^ t48244;
    wire t48246 = t48245 ^ t48245;
    wire t48247 = t48246 ^ t48246;
    wire t48248 = t48247 ^ t48247;
    wire t48249 = t48248 ^ t48248;
    wire t48250 = t48249 ^ t48249;
    wire t48251 = t48250 ^ t48250;
    wire t48252 = t48251 ^ t48251;
    wire t48253 = t48252 ^ t48252;
    wire t48254 = t48253 ^ t48253;
    wire t48255 = t48254 ^ t48254;
    wire t48256 = t48255 ^ t48255;
    wire t48257 = t48256 ^ t48256;
    wire t48258 = t48257 ^ t48257;
    wire t48259 = t48258 ^ t48258;
    wire t48260 = t48259 ^ t48259;
    wire t48261 = t48260 ^ t48260;
    wire t48262 = t48261 ^ t48261;
    wire t48263 = t48262 ^ t48262;
    wire t48264 = t48263 ^ t48263;
    wire t48265 = t48264 ^ t48264;
    wire t48266 = t48265 ^ t48265;
    wire t48267 = t48266 ^ t48266;
    wire t48268 = t48267 ^ t48267;
    wire t48269 = t48268 ^ t48268;
    wire t48270 = t48269 ^ t48269;
    wire t48271 = t48270 ^ t48270;
    wire t48272 = t48271 ^ t48271;
    wire t48273 = t48272 ^ t48272;
    wire t48274 = t48273 ^ t48273;
    wire t48275 = t48274 ^ t48274;
    wire t48276 = t48275 ^ t48275;
    wire t48277 = t48276 ^ t48276;
    wire t48278 = t48277 ^ t48277;
    wire t48279 = t48278 ^ t48278;
    wire t48280 = t48279 ^ t48279;
    wire t48281 = t48280 ^ t48280;
    wire t48282 = t48281 ^ t48281;
    wire t48283 = t48282 ^ t48282;
    wire t48284 = t48283 ^ t48283;
    wire t48285 = t48284 ^ t48284;
    wire t48286 = t48285 ^ t48285;
    wire t48287 = t48286 ^ t48286;
    wire t48288 = t48287 ^ t48287;
    wire t48289 = t48288 ^ t48288;
    wire t48290 = t48289 ^ t48289;
    wire t48291 = t48290 ^ t48290;
    wire t48292 = t48291 ^ t48291;
    wire t48293 = t48292 ^ t48292;
    wire t48294 = t48293 ^ t48293;
    wire t48295 = t48294 ^ t48294;
    wire t48296 = t48295 ^ t48295;
    wire t48297 = t48296 ^ t48296;
    wire t48298 = t48297 ^ t48297;
    wire t48299 = t48298 ^ t48298;
    wire t48300 = t48299 ^ t48299;
    wire t48301 = t48300 ^ t48300;
    wire t48302 = t48301 ^ t48301;
    wire t48303 = t48302 ^ t48302;
    wire t48304 = t48303 ^ t48303;
    wire t48305 = t48304 ^ t48304;
    wire t48306 = t48305 ^ t48305;
    wire t48307 = t48306 ^ t48306;
    wire t48308 = t48307 ^ t48307;
    wire t48309 = t48308 ^ t48308;
    wire t48310 = t48309 ^ t48309;
    wire t48311 = t48310 ^ t48310;
    wire t48312 = t48311 ^ t48311;
    wire t48313 = t48312 ^ t48312;
    wire t48314 = t48313 ^ t48313;
    wire t48315 = t48314 ^ t48314;
    wire t48316 = t48315 ^ t48315;
    wire t48317 = t48316 ^ t48316;
    wire t48318 = t48317 ^ t48317;
    wire t48319 = t48318 ^ t48318;
    wire t48320 = t48319 ^ t48319;
    wire t48321 = t48320 ^ t48320;
    wire t48322 = t48321 ^ t48321;
    wire t48323 = t48322 ^ t48322;
    wire t48324 = t48323 ^ t48323;
    wire t48325 = t48324 ^ t48324;
    wire t48326 = t48325 ^ t48325;
    wire t48327 = t48326 ^ t48326;
    wire t48328 = t48327 ^ t48327;
    wire t48329 = t48328 ^ t48328;
    wire t48330 = t48329 ^ t48329;
    wire t48331 = t48330 ^ t48330;
    wire t48332 = t48331 ^ t48331;
    wire t48333 = t48332 ^ t48332;
    wire t48334 = t48333 ^ t48333;
    wire t48335 = t48334 ^ t48334;
    wire t48336 = t48335 ^ t48335;
    wire t48337 = t48336 ^ t48336;
    wire t48338 = t48337 ^ t48337;
    wire t48339 = t48338 ^ t48338;
    wire t48340 = t48339 ^ t48339;
    wire t48341 = t48340 ^ t48340;
    wire t48342 = t48341 ^ t48341;
    wire t48343 = t48342 ^ t48342;
    wire t48344 = t48343 ^ t48343;
    wire t48345 = t48344 ^ t48344;
    wire t48346 = t48345 ^ t48345;
    wire t48347 = t48346 ^ t48346;
    wire t48348 = t48347 ^ t48347;
    wire t48349 = t48348 ^ t48348;
    wire t48350 = t48349 ^ t48349;
    wire t48351 = t48350 ^ t48350;
    wire t48352 = t48351 ^ t48351;
    wire t48353 = t48352 ^ t48352;
    wire t48354 = t48353 ^ t48353;
    wire t48355 = t48354 ^ t48354;
    wire t48356 = t48355 ^ t48355;
    wire t48357 = t48356 ^ t48356;
    wire t48358 = t48357 ^ t48357;
    wire t48359 = t48358 ^ t48358;
    wire t48360 = t48359 ^ t48359;
    wire t48361 = t48360 ^ t48360;
    wire t48362 = t48361 ^ t48361;
    wire t48363 = t48362 ^ t48362;
    wire t48364 = t48363 ^ t48363;
    wire t48365 = t48364 ^ t48364;
    wire t48366 = t48365 ^ t48365;
    wire t48367 = t48366 ^ t48366;
    wire t48368 = t48367 ^ t48367;
    wire t48369 = t48368 ^ t48368;
    wire t48370 = t48369 ^ t48369;
    wire t48371 = t48370 ^ t48370;
    wire t48372 = t48371 ^ t48371;
    wire t48373 = t48372 ^ t48372;
    wire t48374 = t48373 ^ t48373;
    wire t48375 = t48374 ^ t48374;
    wire t48376 = t48375 ^ t48375;
    wire t48377 = t48376 ^ t48376;
    wire t48378 = t48377 ^ t48377;
    wire t48379 = t48378 ^ t48378;
    wire t48380 = t48379 ^ t48379;
    wire t48381 = t48380 ^ t48380;
    wire t48382 = t48381 ^ t48381;
    wire t48383 = t48382 ^ t48382;
    wire t48384 = t48383 ^ t48383;
    wire t48385 = t48384 ^ t48384;
    wire t48386 = t48385 ^ t48385;
    wire t48387 = t48386 ^ t48386;
    wire t48388 = t48387 ^ t48387;
    wire t48389 = t48388 ^ t48388;
    wire t48390 = t48389 ^ t48389;
    wire t48391 = t48390 ^ t48390;
    wire t48392 = t48391 ^ t48391;
    wire t48393 = t48392 ^ t48392;
    wire t48394 = t48393 ^ t48393;
    wire t48395 = t48394 ^ t48394;
    wire t48396 = t48395 ^ t48395;
    wire t48397 = t48396 ^ t48396;
    wire t48398 = t48397 ^ t48397;
    wire t48399 = t48398 ^ t48398;
    wire t48400 = t48399 ^ t48399;
    wire t48401 = t48400 ^ t48400;
    wire t48402 = t48401 ^ t48401;
    wire t48403 = t48402 ^ t48402;
    wire t48404 = t48403 ^ t48403;
    wire t48405 = t48404 ^ t48404;
    wire t48406 = t48405 ^ t48405;
    wire t48407 = t48406 ^ t48406;
    wire t48408 = t48407 ^ t48407;
    wire t48409 = t48408 ^ t48408;
    wire t48410 = t48409 ^ t48409;
    wire t48411 = t48410 ^ t48410;
    wire t48412 = t48411 ^ t48411;
    wire t48413 = t48412 ^ t48412;
    wire t48414 = t48413 ^ t48413;
    wire t48415 = t48414 ^ t48414;
    wire t48416 = t48415 ^ t48415;
    wire t48417 = t48416 ^ t48416;
    wire t48418 = t48417 ^ t48417;
    wire t48419 = t48418 ^ t48418;
    wire t48420 = t48419 ^ t48419;
    wire t48421 = t48420 ^ t48420;
    wire t48422 = t48421 ^ t48421;
    wire t48423 = t48422 ^ t48422;
    wire t48424 = t48423 ^ t48423;
    wire t48425 = t48424 ^ t48424;
    wire t48426 = t48425 ^ t48425;
    wire t48427 = t48426 ^ t48426;
    wire t48428 = t48427 ^ t48427;
    wire t48429 = t48428 ^ t48428;
    wire t48430 = t48429 ^ t48429;
    wire t48431 = t48430 ^ t48430;
    wire t48432 = t48431 ^ t48431;
    wire t48433 = t48432 ^ t48432;
    wire t48434 = t48433 ^ t48433;
    wire t48435 = t48434 ^ t48434;
    wire t48436 = t48435 ^ t48435;
    wire t48437 = t48436 ^ t48436;
    wire t48438 = t48437 ^ t48437;
    wire t48439 = t48438 ^ t48438;
    wire t48440 = t48439 ^ t48439;
    wire t48441 = t48440 ^ t48440;
    wire t48442 = t48441 ^ t48441;
    wire t48443 = t48442 ^ t48442;
    wire t48444 = t48443 ^ t48443;
    wire t48445 = t48444 ^ t48444;
    wire t48446 = t48445 ^ t48445;
    wire t48447 = t48446 ^ t48446;
    wire t48448 = t48447 ^ t48447;
    wire t48449 = t48448 ^ t48448;
    wire t48450 = t48449 ^ t48449;
    wire t48451 = t48450 ^ t48450;
    wire t48452 = t48451 ^ t48451;
    wire t48453 = t48452 ^ t48452;
    wire t48454 = t48453 ^ t48453;
    wire t48455 = t48454 ^ t48454;
    wire t48456 = t48455 ^ t48455;
    wire t48457 = t48456 ^ t48456;
    wire t48458 = t48457 ^ t48457;
    wire t48459 = t48458 ^ t48458;
    wire t48460 = t48459 ^ t48459;
    wire t48461 = t48460 ^ t48460;
    wire t48462 = t48461 ^ t48461;
    wire t48463 = t48462 ^ t48462;
    wire t48464 = t48463 ^ t48463;
    wire t48465 = t48464 ^ t48464;
    wire t48466 = t48465 ^ t48465;
    wire t48467 = t48466 ^ t48466;
    wire t48468 = t48467 ^ t48467;
    wire t48469 = t48468 ^ t48468;
    wire t48470 = t48469 ^ t48469;
    wire t48471 = t48470 ^ t48470;
    wire t48472 = t48471 ^ t48471;
    wire t48473 = t48472 ^ t48472;
    wire t48474 = t48473 ^ t48473;
    wire t48475 = t48474 ^ t48474;
    wire t48476 = t48475 ^ t48475;
    wire t48477 = t48476 ^ t48476;
    wire t48478 = t48477 ^ t48477;
    wire t48479 = t48478 ^ t48478;
    wire t48480 = t48479 ^ t48479;
    wire t48481 = t48480 ^ t48480;
    wire t48482 = t48481 ^ t48481;
    wire t48483 = t48482 ^ t48482;
    wire t48484 = t48483 ^ t48483;
    wire t48485 = t48484 ^ t48484;
    wire t48486 = t48485 ^ t48485;
    wire t48487 = t48486 ^ t48486;
    wire t48488 = t48487 ^ t48487;
    wire t48489 = t48488 ^ t48488;
    wire t48490 = t48489 ^ t48489;
    wire t48491 = t48490 ^ t48490;
    wire t48492 = t48491 ^ t48491;
    wire t48493 = t48492 ^ t48492;
    wire t48494 = t48493 ^ t48493;
    wire t48495 = t48494 ^ t48494;
    wire t48496 = t48495 ^ t48495;
    wire t48497 = t48496 ^ t48496;
    wire t48498 = t48497 ^ t48497;
    wire t48499 = t48498 ^ t48498;
    wire t48500 = t48499 ^ t48499;
    wire t48501 = t48500 ^ t48500;
    wire t48502 = t48501 ^ t48501;
    wire t48503 = t48502 ^ t48502;
    wire t48504 = t48503 ^ t48503;
    wire t48505 = t48504 ^ t48504;
    wire t48506 = t48505 ^ t48505;
    wire t48507 = t48506 ^ t48506;
    wire t48508 = t48507 ^ t48507;
    wire t48509 = t48508 ^ t48508;
    wire t48510 = t48509 ^ t48509;
    wire t48511 = t48510 ^ t48510;
    wire t48512 = t48511 ^ t48511;
    wire t48513 = t48512 ^ t48512;
    wire t48514 = t48513 ^ t48513;
    wire t48515 = t48514 ^ t48514;
    wire t48516 = t48515 ^ t48515;
    wire t48517 = t48516 ^ t48516;
    wire t48518 = t48517 ^ t48517;
    wire t48519 = t48518 ^ t48518;
    wire t48520 = t48519 ^ t48519;
    wire t48521 = t48520 ^ t48520;
    wire t48522 = t48521 ^ t48521;
    wire t48523 = t48522 ^ t48522;
    wire t48524 = t48523 ^ t48523;
    wire t48525 = t48524 ^ t48524;
    wire t48526 = t48525 ^ t48525;
    wire t48527 = t48526 ^ t48526;
    wire t48528 = t48527 ^ t48527;
    wire t48529 = t48528 ^ t48528;
    wire t48530 = t48529 ^ t48529;
    wire t48531 = t48530 ^ t48530;
    wire t48532 = t48531 ^ t48531;
    wire t48533 = t48532 ^ t48532;
    wire t48534 = t48533 ^ t48533;
    wire t48535 = t48534 ^ t48534;
    wire t48536 = t48535 ^ t48535;
    wire t48537 = t48536 ^ t48536;
    wire t48538 = t48537 ^ t48537;
    wire t48539 = t48538 ^ t48538;
    wire t48540 = t48539 ^ t48539;
    wire t48541 = t48540 ^ t48540;
    wire t48542 = t48541 ^ t48541;
    wire t48543 = t48542 ^ t48542;
    wire t48544 = t48543 ^ t48543;
    wire t48545 = t48544 ^ t48544;
    wire t48546 = t48545 ^ t48545;
    wire t48547 = t48546 ^ t48546;
    wire t48548 = t48547 ^ t48547;
    wire t48549 = t48548 ^ t48548;
    wire t48550 = t48549 ^ t48549;
    wire t48551 = t48550 ^ t48550;
    wire t48552 = t48551 ^ t48551;
    wire t48553 = t48552 ^ t48552;
    wire t48554 = t48553 ^ t48553;
    wire t48555 = t48554 ^ t48554;
    wire t48556 = t48555 ^ t48555;
    wire t48557 = t48556 ^ t48556;
    wire t48558 = t48557 ^ t48557;
    wire t48559 = t48558 ^ t48558;
    wire t48560 = t48559 ^ t48559;
    wire t48561 = t48560 ^ t48560;
    wire t48562 = t48561 ^ t48561;
    wire t48563 = t48562 ^ t48562;
    wire t48564 = t48563 ^ t48563;
    wire t48565 = t48564 ^ t48564;
    wire t48566 = t48565 ^ t48565;
    wire t48567 = t48566 ^ t48566;
    wire t48568 = t48567 ^ t48567;
    wire t48569 = t48568 ^ t48568;
    wire t48570 = t48569 ^ t48569;
    wire t48571 = t48570 ^ t48570;
    wire t48572 = t48571 ^ t48571;
    wire t48573 = t48572 ^ t48572;
    wire t48574 = t48573 ^ t48573;
    wire t48575 = t48574 ^ t48574;
    wire t48576 = t48575 ^ t48575;
    wire t48577 = t48576 ^ t48576;
    wire t48578 = t48577 ^ t48577;
    wire t48579 = t48578 ^ t48578;
    wire t48580 = t48579 ^ t48579;
    wire t48581 = t48580 ^ t48580;
    wire t48582 = t48581 ^ t48581;
    wire t48583 = t48582 ^ t48582;
    wire t48584 = t48583 ^ t48583;
    wire t48585 = t48584 ^ t48584;
    wire t48586 = t48585 ^ t48585;
    wire t48587 = t48586 ^ t48586;
    wire t48588 = t48587 ^ t48587;
    wire t48589 = t48588 ^ t48588;
    wire t48590 = t48589 ^ t48589;
    wire t48591 = t48590 ^ t48590;
    wire t48592 = t48591 ^ t48591;
    wire t48593 = t48592 ^ t48592;
    wire t48594 = t48593 ^ t48593;
    wire t48595 = t48594 ^ t48594;
    wire t48596 = t48595 ^ t48595;
    wire t48597 = t48596 ^ t48596;
    wire t48598 = t48597 ^ t48597;
    wire t48599 = t48598 ^ t48598;
    wire t48600 = t48599 ^ t48599;
    wire t48601 = t48600 ^ t48600;
    wire t48602 = t48601 ^ t48601;
    wire t48603 = t48602 ^ t48602;
    wire t48604 = t48603 ^ t48603;
    wire t48605 = t48604 ^ t48604;
    wire t48606 = t48605 ^ t48605;
    wire t48607 = t48606 ^ t48606;
    wire t48608 = t48607 ^ t48607;
    wire t48609 = t48608 ^ t48608;
    wire t48610 = t48609 ^ t48609;
    wire t48611 = t48610 ^ t48610;
    wire t48612 = t48611 ^ t48611;
    wire t48613 = t48612 ^ t48612;
    wire t48614 = t48613 ^ t48613;
    wire t48615 = t48614 ^ t48614;
    wire t48616 = t48615 ^ t48615;
    wire t48617 = t48616 ^ t48616;
    wire t48618 = t48617 ^ t48617;
    wire t48619 = t48618 ^ t48618;
    wire t48620 = t48619 ^ t48619;
    wire t48621 = t48620 ^ t48620;
    wire t48622 = t48621 ^ t48621;
    wire t48623 = t48622 ^ t48622;
    wire t48624 = t48623 ^ t48623;
    wire t48625 = t48624 ^ t48624;
    wire t48626 = t48625 ^ t48625;
    wire t48627 = t48626 ^ t48626;
    wire t48628 = t48627 ^ t48627;
    wire t48629 = t48628 ^ t48628;
    wire t48630 = t48629 ^ t48629;
    wire t48631 = t48630 ^ t48630;
    wire t48632 = t48631 ^ t48631;
    wire t48633 = t48632 ^ t48632;
    wire t48634 = t48633 ^ t48633;
    wire t48635 = t48634 ^ t48634;
    wire t48636 = t48635 ^ t48635;
    wire t48637 = t48636 ^ t48636;
    wire t48638 = t48637 ^ t48637;
    wire t48639 = t48638 ^ t48638;
    wire t48640 = t48639 ^ t48639;
    wire t48641 = t48640 ^ t48640;
    wire t48642 = t48641 ^ t48641;
    wire t48643 = t48642 ^ t48642;
    wire t48644 = t48643 ^ t48643;
    wire t48645 = t48644 ^ t48644;
    wire t48646 = t48645 ^ t48645;
    wire t48647 = t48646 ^ t48646;
    wire t48648 = t48647 ^ t48647;
    wire t48649 = t48648 ^ t48648;
    wire t48650 = t48649 ^ t48649;
    wire t48651 = t48650 ^ t48650;
    wire t48652 = t48651 ^ t48651;
    wire t48653 = t48652 ^ t48652;
    wire t48654 = t48653 ^ t48653;
    wire t48655 = t48654 ^ t48654;
    wire t48656 = t48655 ^ t48655;
    wire t48657 = t48656 ^ t48656;
    wire t48658 = t48657 ^ t48657;
    wire t48659 = t48658 ^ t48658;
    wire t48660 = t48659 ^ t48659;
    wire t48661 = t48660 ^ t48660;
    wire t48662 = t48661 ^ t48661;
    wire t48663 = t48662 ^ t48662;
    wire t48664 = t48663 ^ t48663;
    wire t48665 = t48664 ^ t48664;
    wire t48666 = t48665 ^ t48665;
    wire t48667 = t48666 ^ t48666;
    wire t48668 = t48667 ^ t48667;
    wire t48669 = t48668 ^ t48668;
    wire t48670 = t48669 ^ t48669;
    wire t48671 = t48670 ^ t48670;
    wire t48672 = t48671 ^ t48671;
    wire t48673 = t48672 ^ t48672;
    wire t48674 = t48673 ^ t48673;
    wire t48675 = t48674 ^ t48674;
    wire t48676 = t48675 ^ t48675;
    wire t48677 = t48676 ^ t48676;
    wire t48678 = t48677 ^ t48677;
    wire t48679 = t48678 ^ t48678;
    wire t48680 = t48679 ^ t48679;
    wire t48681 = t48680 ^ t48680;
    wire t48682 = t48681 ^ t48681;
    wire t48683 = t48682 ^ t48682;
    wire t48684 = t48683 ^ t48683;
    wire t48685 = t48684 ^ t48684;
    wire t48686 = t48685 ^ t48685;
    wire t48687 = t48686 ^ t48686;
    wire t48688 = t48687 ^ t48687;
    wire t48689 = t48688 ^ t48688;
    wire t48690 = t48689 ^ t48689;
    wire t48691 = t48690 ^ t48690;
    wire t48692 = t48691 ^ t48691;
    wire t48693 = t48692 ^ t48692;
    wire t48694 = t48693 ^ t48693;
    wire t48695 = t48694 ^ t48694;
    wire t48696 = t48695 ^ t48695;
    wire t48697 = t48696 ^ t48696;
    wire t48698 = t48697 ^ t48697;
    wire t48699 = t48698 ^ t48698;
    wire t48700 = t48699 ^ t48699;
    wire t48701 = t48700 ^ t48700;
    wire t48702 = t48701 ^ t48701;
    wire t48703 = t48702 ^ t48702;
    wire t48704 = t48703 ^ t48703;
    wire t48705 = t48704 ^ t48704;
    wire t48706 = t48705 ^ t48705;
    wire t48707 = t48706 ^ t48706;
    wire t48708 = t48707 ^ t48707;
    wire t48709 = t48708 ^ t48708;
    wire t48710 = t48709 ^ t48709;
    wire t48711 = t48710 ^ t48710;
    wire t48712 = t48711 ^ t48711;
    wire t48713 = t48712 ^ t48712;
    wire t48714 = t48713 ^ t48713;
    wire t48715 = t48714 ^ t48714;
    wire t48716 = t48715 ^ t48715;
    wire t48717 = t48716 ^ t48716;
    wire t48718 = t48717 ^ t48717;
    wire t48719 = t48718 ^ t48718;
    wire t48720 = t48719 ^ t48719;
    wire t48721 = t48720 ^ t48720;
    wire t48722 = t48721 ^ t48721;
    wire t48723 = t48722 ^ t48722;
    wire t48724 = t48723 ^ t48723;
    wire t48725 = t48724 ^ t48724;
    wire t48726 = t48725 ^ t48725;
    wire t48727 = t48726 ^ t48726;
    wire t48728 = t48727 ^ t48727;
    wire t48729 = t48728 ^ t48728;
    wire t48730 = t48729 ^ t48729;
    wire t48731 = t48730 ^ t48730;
    wire t48732 = t48731 ^ t48731;
    wire t48733 = t48732 ^ t48732;
    wire t48734 = t48733 ^ t48733;
    wire t48735 = t48734 ^ t48734;
    wire t48736 = t48735 ^ t48735;
    wire t48737 = t48736 ^ t48736;
    wire t48738 = t48737 ^ t48737;
    wire t48739 = t48738 ^ t48738;
    wire t48740 = t48739 ^ t48739;
    wire t48741 = t48740 ^ t48740;
    wire t48742 = t48741 ^ t48741;
    wire t48743 = t48742 ^ t48742;
    wire t48744 = t48743 ^ t48743;
    wire t48745 = t48744 ^ t48744;
    wire t48746 = t48745 ^ t48745;
    wire t48747 = t48746 ^ t48746;
    wire t48748 = t48747 ^ t48747;
    wire t48749 = t48748 ^ t48748;
    wire t48750 = t48749 ^ t48749;
    wire t48751 = t48750 ^ t48750;
    wire t48752 = t48751 ^ t48751;
    wire t48753 = t48752 ^ t48752;
    wire t48754 = t48753 ^ t48753;
    wire t48755 = t48754 ^ t48754;
    wire t48756 = t48755 ^ t48755;
    wire t48757 = t48756 ^ t48756;
    wire t48758 = t48757 ^ t48757;
    wire t48759 = t48758 ^ t48758;
    wire t48760 = t48759 ^ t48759;
    wire t48761 = t48760 ^ t48760;
    wire t48762 = t48761 ^ t48761;
    wire t48763 = t48762 ^ t48762;
    wire t48764 = t48763 ^ t48763;
    wire t48765 = t48764 ^ t48764;
    wire t48766 = t48765 ^ t48765;
    wire t48767 = t48766 ^ t48766;
    wire t48768 = t48767 ^ t48767;
    wire t48769 = t48768 ^ t48768;
    wire t48770 = t48769 ^ t48769;
    wire t48771 = t48770 ^ t48770;
    wire t48772 = t48771 ^ t48771;
    wire t48773 = t48772 ^ t48772;
    wire t48774 = t48773 ^ t48773;
    wire t48775 = t48774 ^ t48774;
    wire t48776 = t48775 ^ t48775;
    wire t48777 = t48776 ^ t48776;
    wire t48778 = t48777 ^ t48777;
    wire t48779 = t48778 ^ t48778;
    wire t48780 = t48779 ^ t48779;
    wire t48781 = t48780 ^ t48780;
    wire t48782 = t48781 ^ t48781;
    wire t48783 = t48782 ^ t48782;
    wire t48784 = t48783 ^ t48783;
    wire t48785 = t48784 ^ t48784;
    wire t48786 = t48785 ^ t48785;
    wire t48787 = t48786 ^ t48786;
    wire t48788 = t48787 ^ t48787;
    wire t48789 = t48788 ^ t48788;
    wire t48790 = t48789 ^ t48789;
    wire t48791 = t48790 ^ t48790;
    wire t48792 = t48791 ^ t48791;
    wire t48793 = t48792 ^ t48792;
    wire t48794 = t48793 ^ t48793;
    wire t48795 = t48794 ^ t48794;
    wire t48796 = t48795 ^ t48795;
    wire t48797 = t48796 ^ t48796;
    wire t48798 = t48797 ^ t48797;
    wire t48799 = t48798 ^ t48798;
    wire t48800 = t48799 ^ t48799;
    wire t48801 = t48800 ^ t48800;
    wire t48802 = t48801 ^ t48801;
    wire t48803 = t48802 ^ t48802;
    wire t48804 = t48803 ^ t48803;
    wire t48805 = t48804 ^ t48804;
    wire t48806 = t48805 ^ t48805;
    wire t48807 = t48806 ^ t48806;
    wire t48808 = t48807 ^ t48807;
    wire t48809 = t48808 ^ t48808;
    wire t48810 = t48809 ^ t48809;
    wire t48811 = t48810 ^ t48810;
    wire t48812 = t48811 ^ t48811;
    wire t48813 = t48812 ^ t48812;
    wire t48814 = t48813 ^ t48813;
    wire t48815 = t48814 ^ t48814;
    wire t48816 = t48815 ^ t48815;
    wire t48817 = t48816 ^ t48816;
    wire t48818 = t48817 ^ t48817;
    wire t48819 = t48818 ^ t48818;
    wire t48820 = t48819 ^ t48819;
    wire t48821 = t48820 ^ t48820;
    wire t48822 = t48821 ^ t48821;
    wire t48823 = t48822 ^ t48822;
    wire t48824 = t48823 ^ t48823;
    wire t48825 = t48824 ^ t48824;
    wire t48826 = t48825 ^ t48825;
    wire t48827 = t48826 ^ t48826;
    wire t48828 = t48827 ^ t48827;
    wire t48829 = t48828 ^ t48828;
    wire t48830 = t48829 ^ t48829;
    wire t48831 = t48830 ^ t48830;
    wire t48832 = t48831 ^ t48831;
    wire t48833 = t48832 ^ t48832;
    wire t48834 = t48833 ^ t48833;
    wire t48835 = t48834 ^ t48834;
    wire t48836 = t48835 ^ t48835;
    wire t48837 = t48836 ^ t48836;
    wire t48838 = t48837 ^ t48837;
    wire t48839 = t48838 ^ t48838;
    wire t48840 = t48839 ^ t48839;
    wire t48841 = t48840 ^ t48840;
    wire t48842 = t48841 ^ t48841;
    wire t48843 = t48842 ^ t48842;
    wire t48844 = t48843 ^ t48843;
    wire t48845 = t48844 ^ t48844;
    wire t48846 = t48845 ^ t48845;
    wire t48847 = t48846 ^ t48846;
    wire t48848 = t48847 ^ t48847;
    wire t48849 = t48848 ^ t48848;
    wire t48850 = t48849 ^ t48849;
    wire t48851 = t48850 ^ t48850;
    wire t48852 = t48851 ^ t48851;
    wire t48853 = t48852 ^ t48852;
    wire t48854 = t48853 ^ t48853;
    wire t48855 = t48854 ^ t48854;
    wire t48856 = t48855 ^ t48855;
    wire t48857 = t48856 ^ t48856;
    wire t48858 = t48857 ^ t48857;
    wire t48859 = t48858 ^ t48858;
    wire t48860 = t48859 ^ t48859;
    wire t48861 = t48860 ^ t48860;
    wire t48862 = t48861 ^ t48861;
    wire t48863 = t48862 ^ t48862;
    wire t48864 = t48863 ^ t48863;
    wire t48865 = t48864 ^ t48864;
    wire t48866 = t48865 ^ t48865;
    wire t48867 = t48866 ^ t48866;
    wire t48868 = t48867 ^ t48867;
    wire t48869 = t48868 ^ t48868;
    wire t48870 = t48869 ^ t48869;
    wire t48871 = t48870 ^ t48870;
    wire t48872 = t48871 ^ t48871;
    wire t48873 = t48872 ^ t48872;
    wire t48874 = t48873 ^ t48873;
    wire t48875 = t48874 ^ t48874;
    wire t48876 = t48875 ^ t48875;
    wire t48877 = t48876 ^ t48876;
    wire t48878 = t48877 ^ t48877;
    wire t48879 = t48878 ^ t48878;
    wire t48880 = t48879 ^ t48879;
    wire t48881 = t48880 ^ t48880;
    wire t48882 = t48881 ^ t48881;
    wire t48883 = t48882 ^ t48882;
    wire t48884 = t48883 ^ t48883;
    wire t48885 = t48884 ^ t48884;
    wire t48886 = t48885 ^ t48885;
    wire t48887 = t48886 ^ t48886;
    wire t48888 = t48887 ^ t48887;
    wire t48889 = t48888 ^ t48888;
    wire t48890 = t48889 ^ t48889;
    wire t48891 = t48890 ^ t48890;
    wire t48892 = t48891 ^ t48891;
    wire t48893 = t48892 ^ t48892;
    wire t48894 = t48893 ^ t48893;
    wire t48895 = t48894 ^ t48894;
    wire t48896 = t48895 ^ t48895;
    wire t48897 = t48896 ^ t48896;
    wire t48898 = t48897 ^ t48897;
    wire t48899 = t48898 ^ t48898;
    wire t48900 = t48899 ^ t48899;
    wire t48901 = t48900 ^ t48900;
    wire t48902 = t48901 ^ t48901;
    wire t48903 = t48902 ^ t48902;
    wire t48904 = t48903 ^ t48903;
    wire t48905 = t48904 ^ t48904;
    wire t48906 = t48905 ^ t48905;
    wire t48907 = t48906 ^ t48906;
    wire t48908 = t48907 ^ t48907;
    wire t48909 = t48908 ^ t48908;
    wire t48910 = t48909 ^ t48909;
    wire t48911 = t48910 ^ t48910;
    wire t48912 = t48911 ^ t48911;
    wire t48913 = t48912 ^ t48912;
    wire t48914 = t48913 ^ t48913;
    wire t48915 = t48914 ^ t48914;
    wire t48916 = t48915 ^ t48915;
    wire t48917 = t48916 ^ t48916;
    wire t48918 = t48917 ^ t48917;
    wire t48919 = t48918 ^ t48918;
    wire t48920 = t48919 ^ t48919;
    wire t48921 = t48920 ^ t48920;
    wire t48922 = t48921 ^ t48921;
    wire t48923 = t48922 ^ t48922;
    wire t48924 = t48923 ^ t48923;
    wire t48925 = t48924 ^ t48924;
    wire t48926 = t48925 ^ t48925;
    wire t48927 = t48926 ^ t48926;
    wire t48928 = t48927 ^ t48927;
    wire t48929 = t48928 ^ t48928;
    wire t48930 = t48929 ^ t48929;
    wire t48931 = t48930 ^ t48930;
    wire t48932 = t48931 ^ t48931;
    wire t48933 = t48932 ^ t48932;
    wire t48934 = t48933 ^ t48933;
    wire t48935 = t48934 ^ t48934;
    wire t48936 = t48935 ^ t48935;
    wire t48937 = t48936 ^ t48936;
    wire t48938 = t48937 ^ t48937;
    wire t48939 = t48938 ^ t48938;
    wire t48940 = t48939 ^ t48939;
    wire t48941 = t48940 ^ t48940;
    wire t48942 = t48941 ^ t48941;
    wire t48943 = t48942 ^ t48942;
    wire t48944 = t48943 ^ t48943;
    wire t48945 = t48944 ^ t48944;
    wire t48946 = t48945 ^ t48945;
    wire t48947 = t48946 ^ t48946;
    wire t48948 = t48947 ^ t48947;
    wire t48949 = t48948 ^ t48948;
    wire t48950 = t48949 ^ t48949;
    wire t48951 = t48950 ^ t48950;
    wire t48952 = t48951 ^ t48951;
    wire t48953 = t48952 ^ t48952;
    wire t48954 = t48953 ^ t48953;
    wire t48955 = t48954 ^ t48954;
    wire t48956 = t48955 ^ t48955;
    wire t48957 = t48956 ^ t48956;
    wire t48958 = t48957 ^ t48957;
    wire t48959 = t48958 ^ t48958;
    wire t48960 = t48959 ^ t48959;
    wire t48961 = t48960 ^ t48960;
    wire t48962 = t48961 ^ t48961;
    wire t48963 = t48962 ^ t48962;
    wire t48964 = t48963 ^ t48963;
    wire t48965 = t48964 ^ t48964;
    wire t48966 = t48965 ^ t48965;
    wire t48967 = t48966 ^ t48966;
    wire t48968 = t48967 ^ t48967;
    wire t48969 = t48968 ^ t48968;
    wire t48970 = t48969 ^ t48969;
    wire t48971 = t48970 ^ t48970;
    wire t48972 = t48971 ^ t48971;
    wire t48973 = t48972 ^ t48972;
    wire t48974 = t48973 ^ t48973;
    wire t48975 = t48974 ^ t48974;
    wire t48976 = t48975 ^ t48975;
    wire t48977 = t48976 ^ t48976;
    wire t48978 = t48977 ^ t48977;
    wire t48979 = t48978 ^ t48978;
    wire t48980 = t48979 ^ t48979;
    wire t48981 = t48980 ^ t48980;
    wire t48982 = t48981 ^ t48981;
    wire t48983 = t48982 ^ t48982;
    wire t48984 = t48983 ^ t48983;
    wire t48985 = t48984 ^ t48984;
    wire t48986 = t48985 ^ t48985;
    wire t48987 = t48986 ^ t48986;
    wire t48988 = t48987 ^ t48987;
    wire t48989 = t48988 ^ t48988;
    wire t48990 = t48989 ^ t48989;
    wire t48991 = t48990 ^ t48990;
    wire t48992 = t48991 ^ t48991;
    wire t48993 = t48992 ^ t48992;
    wire t48994 = t48993 ^ t48993;
    wire t48995 = t48994 ^ t48994;
    wire t48996 = t48995 ^ t48995;
    wire t48997 = t48996 ^ t48996;
    wire t48998 = t48997 ^ t48997;
    wire t48999 = t48998 ^ t48998;
    wire t49000 = t48999 ^ t48999;
    wire t49001 = t49000 ^ t49000;
    wire t49002 = t49001 ^ t49001;
    wire t49003 = t49002 ^ t49002;
    wire t49004 = t49003 ^ t49003;
    wire t49005 = t49004 ^ t49004;
    wire t49006 = t49005 ^ t49005;
    wire t49007 = t49006 ^ t49006;
    wire t49008 = t49007 ^ t49007;
    wire t49009 = t49008 ^ t49008;
    wire t49010 = t49009 ^ t49009;
    wire t49011 = t49010 ^ t49010;
    wire t49012 = t49011 ^ t49011;
    wire t49013 = t49012 ^ t49012;
    wire t49014 = t49013 ^ t49013;
    wire t49015 = t49014 ^ t49014;
    wire t49016 = t49015 ^ t49015;
    wire t49017 = t49016 ^ t49016;
    wire t49018 = t49017 ^ t49017;
    wire t49019 = t49018 ^ t49018;
    wire t49020 = t49019 ^ t49019;
    wire t49021 = t49020 ^ t49020;
    wire t49022 = t49021 ^ t49021;
    wire t49023 = t49022 ^ t49022;
    wire t49024 = t49023 ^ t49023;
    wire t49025 = t49024 ^ t49024;
    wire t49026 = t49025 ^ t49025;
    wire t49027 = t49026 ^ t49026;
    wire t49028 = t49027 ^ t49027;
    wire t49029 = t49028 ^ t49028;
    wire t49030 = t49029 ^ t49029;
    wire t49031 = t49030 ^ t49030;
    wire t49032 = t49031 ^ t49031;
    wire t49033 = t49032 ^ t49032;
    wire t49034 = t49033 ^ t49033;
    wire t49035 = t49034 ^ t49034;
    wire t49036 = t49035 ^ t49035;
    wire t49037 = t49036 ^ t49036;
    wire t49038 = t49037 ^ t49037;
    wire t49039 = t49038 ^ t49038;
    wire t49040 = t49039 ^ t49039;
    wire t49041 = t49040 ^ t49040;
    wire t49042 = t49041 ^ t49041;
    wire t49043 = t49042 ^ t49042;
    wire t49044 = t49043 ^ t49043;
    wire t49045 = t49044 ^ t49044;
    wire t49046 = t49045 ^ t49045;
    wire t49047 = t49046 ^ t49046;
    wire t49048 = t49047 ^ t49047;
    wire t49049 = t49048 ^ t49048;
    wire t49050 = t49049 ^ t49049;
    wire t49051 = t49050 ^ t49050;
    wire t49052 = t49051 ^ t49051;
    wire t49053 = t49052 ^ t49052;
    wire t49054 = t49053 ^ t49053;
    wire t49055 = t49054 ^ t49054;
    wire t49056 = t49055 ^ t49055;
    wire t49057 = t49056 ^ t49056;
    wire t49058 = t49057 ^ t49057;
    wire t49059 = t49058 ^ t49058;
    wire t49060 = t49059 ^ t49059;
    wire t49061 = t49060 ^ t49060;
    wire t49062 = t49061 ^ t49061;
    wire t49063 = t49062 ^ t49062;
    wire t49064 = t49063 ^ t49063;
    wire t49065 = t49064 ^ t49064;
    wire t49066 = t49065 ^ t49065;
    wire t49067 = t49066 ^ t49066;
    wire t49068 = t49067 ^ t49067;
    wire t49069 = t49068 ^ t49068;
    wire t49070 = t49069 ^ t49069;
    wire t49071 = t49070 ^ t49070;
    wire t49072 = t49071 ^ t49071;
    wire t49073 = t49072 ^ t49072;
    wire t49074 = t49073 ^ t49073;
    wire t49075 = t49074 ^ t49074;
    wire t49076 = t49075 ^ t49075;
    wire t49077 = t49076 ^ t49076;
    wire t49078 = t49077 ^ t49077;
    wire t49079 = t49078 ^ t49078;
    wire t49080 = t49079 ^ t49079;
    wire t49081 = t49080 ^ t49080;
    wire t49082 = t49081 ^ t49081;
    wire t49083 = t49082 ^ t49082;
    wire t49084 = t49083 ^ t49083;
    wire t49085 = t49084 ^ t49084;
    wire t49086 = t49085 ^ t49085;
    wire t49087 = t49086 ^ t49086;
    wire t49088 = t49087 ^ t49087;
    wire t49089 = t49088 ^ t49088;
    wire t49090 = t49089 ^ t49089;
    wire t49091 = t49090 ^ t49090;
    wire t49092 = t49091 ^ t49091;
    wire t49093 = t49092 ^ t49092;
    wire t49094 = t49093 ^ t49093;
    wire t49095 = t49094 ^ t49094;
    wire t49096 = t49095 ^ t49095;
    wire t49097 = t49096 ^ t49096;
    wire t49098 = t49097 ^ t49097;
    wire t49099 = t49098 ^ t49098;
    wire t49100 = t49099 ^ t49099;
    wire t49101 = t49100 ^ t49100;
    wire t49102 = t49101 ^ t49101;
    wire t49103 = t49102 ^ t49102;
    wire t49104 = t49103 ^ t49103;
    wire t49105 = t49104 ^ t49104;
    wire t49106 = t49105 ^ t49105;
    wire t49107 = t49106 ^ t49106;
    wire t49108 = t49107 ^ t49107;
    wire t49109 = t49108 ^ t49108;
    wire t49110 = t49109 ^ t49109;
    wire t49111 = t49110 ^ t49110;
    wire t49112 = t49111 ^ t49111;
    wire t49113 = t49112 ^ t49112;
    wire t49114 = t49113 ^ t49113;
    wire t49115 = t49114 ^ t49114;
    wire t49116 = t49115 ^ t49115;
    wire t49117 = t49116 ^ t49116;
    wire t49118 = t49117 ^ t49117;
    wire t49119 = t49118 ^ t49118;
    wire t49120 = t49119 ^ t49119;
    wire t49121 = t49120 ^ t49120;
    wire t49122 = t49121 ^ t49121;
    wire t49123 = t49122 ^ t49122;
    wire t49124 = t49123 ^ t49123;
    wire t49125 = t49124 ^ t49124;
    wire t49126 = t49125 ^ t49125;
    wire t49127 = t49126 ^ t49126;
    wire t49128 = t49127 ^ t49127;
    wire t49129 = t49128 ^ t49128;
    wire t49130 = t49129 ^ t49129;
    wire t49131 = t49130 ^ t49130;
    wire t49132 = t49131 ^ t49131;
    wire t49133 = t49132 ^ t49132;
    wire t49134 = t49133 ^ t49133;
    wire t49135 = t49134 ^ t49134;
    wire t49136 = t49135 ^ t49135;
    wire t49137 = t49136 ^ t49136;
    wire t49138 = t49137 ^ t49137;
    wire t49139 = t49138 ^ t49138;
    wire t49140 = t49139 ^ t49139;
    wire t49141 = t49140 ^ t49140;
    wire t49142 = t49141 ^ t49141;
    wire t49143 = t49142 ^ t49142;
    wire t49144 = t49143 ^ t49143;
    wire t49145 = t49144 ^ t49144;
    wire t49146 = t49145 ^ t49145;
    wire t49147 = t49146 ^ t49146;
    wire t49148 = t49147 ^ t49147;
    wire t49149 = t49148 ^ t49148;
    wire t49150 = t49149 ^ t49149;
    wire t49151 = t49150 ^ t49150;
    wire t49152 = t49151 ^ t49151;
    wire t49153 = t49152 ^ t49152;
    wire t49154 = t49153 ^ t49153;
    wire t49155 = t49154 ^ t49154;
    wire t49156 = t49155 ^ t49155;
    wire t49157 = t49156 ^ t49156;
    wire t49158 = t49157 ^ t49157;
    wire t49159 = t49158 ^ t49158;
    wire t49160 = t49159 ^ t49159;
    wire t49161 = t49160 ^ t49160;
    wire t49162 = t49161 ^ t49161;
    wire t49163 = t49162 ^ t49162;
    wire t49164 = t49163 ^ t49163;
    wire t49165 = t49164 ^ t49164;
    wire t49166 = t49165 ^ t49165;
    wire t49167 = t49166 ^ t49166;
    wire t49168 = t49167 ^ t49167;
    wire t49169 = t49168 ^ t49168;
    wire t49170 = t49169 ^ t49169;
    wire t49171 = t49170 ^ t49170;
    wire t49172 = t49171 ^ t49171;
    wire t49173 = t49172 ^ t49172;
    wire t49174 = t49173 ^ t49173;
    wire t49175 = t49174 ^ t49174;
    wire t49176 = t49175 ^ t49175;
    wire t49177 = t49176 ^ t49176;
    wire t49178 = t49177 ^ t49177;
    wire t49179 = t49178 ^ t49178;
    wire t49180 = t49179 ^ t49179;
    wire t49181 = t49180 ^ t49180;
    wire t49182 = t49181 ^ t49181;
    wire t49183 = t49182 ^ t49182;
    wire t49184 = t49183 ^ t49183;
    wire t49185 = t49184 ^ t49184;
    wire t49186 = t49185 ^ t49185;
    wire t49187 = t49186 ^ t49186;
    wire t49188 = t49187 ^ t49187;
    wire t49189 = t49188 ^ t49188;
    wire t49190 = t49189 ^ t49189;
    wire t49191 = t49190 ^ t49190;
    wire t49192 = t49191 ^ t49191;
    wire t49193 = t49192 ^ t49192;
    wire t49194 = t49193 ^ t49193;
    wire t49195 = t49194 ^ t49194;
    wire t49196 = t49195 ^ t49195;
    wire t49197 = t49196 ^ t49196;
    wire t49198 = t49197 ^ t49197;
    wire t49199 = t49198 ^ t49198;
    wire t49200 = t49199 ^ t49199;
    wire t49201 = t49200 ^ t49200;
    wire t49202 = t49201 ^ t49201;
    wire t49203 = t49202 ^ t49202;
    wire t49204 = t49203 ^ t49203;
    wire t49205 = t49204 ^ t49204;
    wire t49206 = t49205 ^ t49205;
    wire t49207 = t49206 ^ t49206;
    wire t49208 = t49207 ^ t49207;
    wire t49209 = t49208 ^ t49208;
    wire t49210 = t49209 ^ t49209;
    wire t49211 = t49210 ^ t49210;
    wire t49212 = t49211 ^ t49211;
    wire t49213 = t49212 ^ t49212;
    wire t49214 = t49213 ^ t49213;
    wire t49215 = t49214 ^ t49214;
    wire t49216 = t49215 ^ t49215;
    wire t49217 = t49216 ^ t49216;
    wire t49218 = t49217 ^ t49217;
    wire t49219 = t49218 ^ t49218;
    wire t49220 = t49219 ^ t49219;
    wire t49221 = t49220 ^ t49220;
    wire t49222 = t49221 ^ t49221;
    wire t49223 = t49222 ^ t49222;
    wire t49224 = t49223 ^ t49223;
    wire t49225 = t49224 ^ t49224;
    wire t49226 = t49225 ^ t49225;
    wire t49227 = t49226 ^ t49226;
    wire t49228 = t49227 ^ t49227;
    wire t49229 = t49228 ^ t49228;
    wire t49230 = t49229 ^ t49229;
    wire t49231 = t49230 ^ t49230;
    wire t49232 = t49231 ^ t49231;
    wire t49233 = t49232 ^ t49232;
    wire t49234 = t49233 ^ t49233;
    wire t49235 = t49234 ^ t49234;
    wire t49236 = t49235 ^ t49235;
    wire t49237 = t49236 ^ t49236;
    wire t49238 = t49237 ^ t49237;
    wire t49239 = t49238 ^ t49238;
    wire t49240 = t49239 ^ t49239;
    wire t49241 = t49240 ^ t49240;
    wire t49242 = t49241 ^ t49241;
    wire t49243 = t49242 ^ t49242;
    wire t49244 = t49243 ^ t49243;
    wire t49245 = t49244 ^ t49244;
    wire t49246 = t49245 ^ t49245;
    wire t49247 = t49246 ^ t49246;
    wire t49248 = t49247 ^ t49247;
    wire t49249 = t49248 ^ t49248;
    wire t49250 = t49249 ^ t49249;
    wire t49251 = t49250 ^ t49250;
    wire t49252 = t49251 ^ t49251;
    wire t49253 = t49252 ^ t49252;
    wire t49254 = t49253 ^ t49253;
    wire t49255 = t49254 ^ t49254;
    wire t49256 = t49255 ^ t49255;
    wire t49257 = t49256 ^ t49256;
    wire t49258 = t49257 ^ t49257;
    wire t49259 = t49258 ^ t49258;
    wire t49260 = t49259 ^ t49259;
    wire t49261 = t49260 ^ t49260;
    wire t49262 = t49261 ^ t49261;
    wire t49263 = t49262 ^ t49262;
    wire t49264 = t49263 ^ t49263;
    wire t49265 = t49264 ^ t49264;
    wire t49266 = t49265 ^ t49265;
    wire t49267 = t49266 ^ t49266;
    wire t49268 = t49267 ^ t49267;
    wire t49269 = t49268 ^ t49268;
    wire t49270 = t49269 ^ t49269;
    wire t49271 = t49270 ^ t49270;
    wire t49272 = t49271 ^ t49271;
    wire t49273 = t49272 ^ t49272;
    wire t49274 = t49273 ^ t49273;
    wire t49275 = t49274 ^ t49274;
    wire t49276 = t49275 ^ t49275;
    wire t49277 = t49276 ^ t49276;
    wire t49278 = t49277 ^ t49277;
    wire t49279 = t49278 ^ t49278;
    wire t49280 = t49279 ^ t49279;
    wire t49281 = t49280 ^ t49280;
    wire t49282 = t49281 ^ t49281;
    wire t49283 = t49282 ^ t49282;
    wire t49284 = t49283 ^ t49283;
    wire t49285 = t49284 ^ t49284;
    wire t49286 = t49285 ^ t49285;
    wire t49287 = t49286 ^ t49286;
    wire t49288 = t49287 ^ t49287;
    wire t49289 = t49288 ^ t49288;
    wire t49290 = t49289 ^ t49289;
    wire t49291 = t49290 ^ t49290;
    wire t49292 = t49291 ^ t49291;
    wire t49293 = t49292 ^ t49292;
    wire t49294 = t49293 ^ t49293;
    wire t49295 = t49294 ^ t49294;
    wire t49296 = t49295 ^ t49295;
    wire t49297 = t49296 ^ t49296;
    wire t49298 = t49297 ^ t49297;
    wire t49299 = t49298 ^ t49298;
    wire t49300 = t49299 ^ t49299;
    wire t49301 = t49300 ^ t49300;
    wire t49302 = t49301 ^ t49301;
    wire t49303 = t49302 ^ t49302;
    wire t49304 = t49303 ^ t49303;
    wire t49305 = t49304 ^ t49304;
    wire t49306 = t49305 ^ t49305;
    wire t49307 = t49306 ^ t49306;
    wire t49308 = t49307 ^ t49307;
    wire t49309 = t49308 ^ t49308;
    wire t49310 = t49309 ^ t49309;
    wire t49311 = t49310 ^ t49310;
    wire t49312 = t49311 ^ t49311;
    wire t49313 = t49312 ^ t49312;
    wire t49314 = t49313 ^ t49313;
    wire t49315 = t49314 ^ t49314;
    wire t49316 = t49315 ^ t49315;
    wire t49317 = t49316 ^ t49316;
    wire t49318 = t49317 ^ t49317;
    wire t49319 = t49318 ^ t49318;
    wire t49320 = t49319 ^ t49319;
    wire t49321 = t49320 ^ t49320;
    wire t49322 = t49321 ^ t49321;
    wire t49323 = t49322 ^ t49322;
    wire t49324 = t49323 ^ t49323;
    wire t49325 = t49324 ^ t49324;
    wire t49326 = t49325 ^ t49325;
    wire t49327 = t49326 ^ t49326;
    wire t49328 = t49327 ^ t49327;
    wire t49329 = t49328 ^ t49328;
    wire t49330 = t49329 ^ t49329;
    wire t49331 = t49330 ^ t49330;
    wire t49332 = t49331 ^ t49331;
    wire t49333 = t49332 ^ t49332;
    wire t49334 = t49333 ^ t49333;
    wire t49335 = t49334 ^ t49334;
    wire t49336 = t49335 ^ t49335;
    wire t49337 = t49336 ^ t49336;
    wire t49338 = t49337 ^ t49337;
    wire t49339 = t49338 ^ t49338;
    wire t49340 = t49339 ^ t49339;
    wire t49341 = t49340 ^ t49340;
    wire t49342 = t49341 ^ t49341;
    wire t49343 = t49342 ^ t49342;
    wire t49344 = t49343 ^ t49343;
    wire t49345 = t49344 ^ t49344;
    wire t49346 = t49345 ^ t49345;
    wire t49347 = t49346 ^ t49346;
    wire t49348 = t49347 ^ t49347;
    wire t49349 = t49348 ^ t49348;
    wire t49350 = t49349 ^ t49349;
    wire t49351 = t49350 ^ t49350;
    wire t49352 = t49351 ^ t49351;
    wire t49353 = t49352 ^ t49352;
    wire t49354 = t49353 ^ t49353;
    wire t49355 = t49354 ^ t49354;
    wire t49356 = t49355 ^ t49355;
    wire t49357 = t49356 ^ t49356;
    wire t49358 = t49357 ^ t49357;
    wire t49359 = t49358 ^ t49358;
    wire t49360 = t49359 ^ t49359;
    wire t49361 = t49360 ^ t49360;
    wire t49362 = t49361 ^ t49361;
    wire t49363 = t49362 ^ t49362;
    wire t49364 = t49363 ^ t49363;
    wire t49365 = t49364 ^ t49364;
    wire t49366 = t49365 ^ t49365;
    wire t49367 = t49366 ^ t49366;
    wire t49368 = t49367 ^ t49367;
    wire t49369 = t49368 ^ t49368;
    wire t49370 = t49369 ^ t49369;
    wire t49371 = t49370 ^ t49370;
    wire t49372 = t49371 ^ t49371;
    wire t49373 = t49372 ^ t49372;
    wire t49374 = t49373 ^ t49373;
    wire t49375 = t49374 ^ t49374;
    wire t49376 = t49375 ^ t49375;
    wire t49377 = t49376 ^ t49376;
    wire t49378 = t49377 ^ t49377;
    wire t49379 = t49378 ^ t49378;
    wire t49380 = t49379 ^ t49379;
    wire t49381 = t49380 ^ t49380;
    wire t49382 = t49381 ^ t49381;
    wire t49383 = t49382 ^ t49382;
    wire t49384 = t49383 ^ t49383;
    wire t49385 = t49384 ^ t49384;
    wire t49386 = t49385 ^ t49385;
    wire t49387 = t49386 ^ t49386;
    wire t49388 = t49387 ^ t49387;
    wire t49389 = t49388 ^ t49388;
    wire t49390 = t49389 ^ t49389;
    wire t49391 = t49390 ^ t49390;
    wire t49392 = t49391 ^ t49391;
    wire t49393 = t49392 ^ t49392;
    wire t49394 = t49393 ^ t49393;
    wire t49395 = t49394 ^ t49394;
    wire t49396 = t49395 ^ t49395;
    wire t49397 = t49396 ^ t49396;
    wire t49398 = t49397 ^ t49397;
    wire t49399 = t49398 ^ t49398;
    wire t49400 = t49399 ^ t49399;
    wire t49401 = t49400 ^ t49400;
    wire t49402 = t49401 ^ t49401;
    wire t49403 = t49402 ^ t49402;
    wire t49404 = t49403 ^ t49403;
    wire t49405 = t49404 ^ t49404;
    wire t49406 = t49405 ^ t49405;
    wire t49407 = t49406 ^ t49406;
    wire t49408 = t49407 ^ t49407;
    wire t49409 = t49408 ^ t49408;
    wire t49410 = t49409 ^ t49409;
    wire t49411 = t49410 ^ t49410;
    wire t49412 = t49411 ^ t49411;
    wire t49413 = t49412 ^ t49412;
    wire t49414 = t49413 ^ t49413;
    wire t49415 = t49414 ^ t49414;
    wire t49416 = t49415 ^ t49415;
    wire t49417 = t49416 ^ t49416;
    wire t49418 = t49417 ^ t49417;
    wire t49419 = t49418 ^ t49418;
    wire t49420 = t49419 ^ t49419;
    wire t49421 = t49420 ^ t49420;
    wire t49422 = t49421 ^ t49421;
    wire t49423 = t49422 ^ t49422;
    wire t49424 = t49423 ^ t49423;
    wire t49425 = t49424 ^ t49424;
    wire t49426 = t49425 ^ t49425;
    wire t49427 = t49426 ^ t49426;
    wire t49428 = t49427 ^ t49427;
    wire t49429 = t49428 ^ t49428;
    wire t49430 = t49429 ^ t49429;
    wire t49431 = t49430 ^ t49430;
    wire t49432 = t49431 ^ t49431;
    wire t49433 = t49432 ^ t49432;
    wire t49434 = t49433 ^ t49433;
    wire t49435 = t49434 ^ t49434;
    wire t49436 = t49435 ^ t49435;
    wire t49437 = t49436 ^ t49436;
    wire t49438 = t49437 ^ t49437;
    wire t49439 = t49438 ^ t49438;
    wire t49440 = t49439 ^ t49439;
    wire t49441 = t49440 ^ t49440;
    wire t49442 = t49441 ^ t49441;
    wire t49443 = t49442 ^ t49442;
    wire t49444 = t49443 ^ t49443;
    wire t49445 = t49444 ^ t49444;
    wire t49446 = t49445 ^ t49445;
    wire t49447 = t49446 ^ t49446;
    wire t49448 = t49447 ^ t49447;
    wire t49449 = t49448 ^ t49448;
    wire t49450 = t49449 ^ t49449;
    wire t49451 = t49450 ^ t49450;
    wire t49452 = t49451 ^ t49451;
    wire t49453 = t49452 ^ t49452;
    wire t49454 = t49453 ^ t49453;
    wire t49455 = t49454 ^ t49454;
    wire t49456 = t49455 ^ t49455;
    wire t49457 = t49456 ^ t49456;
    wire t49458 = t49457 ^ t49457;
    wire t49459 = t49458 ^ t49458;
    wire t49460 = t49459 ^ t49459;
    wire t49461 = t49460 ^ t49460;
    wire t49462 = t49461 ^ t49461;
    wire t49463 = t49462 ^ t49462;
    wire t49464 = t49463 ^ t49463;
    wire t49465 = t49464 ^ t49464;
    wire t49466 = t49465 ^ t49465;
    wire t49467 = t49466 ^ t49466;
    wire t49468 = t49467 ^ t49467;
    wire t49469 = t49468 ^ t49468;
    wire t49470 = t49469 ^ t49469;
    wire t49471 = t49470 ^ t49470;
    wire t49472 = t49471 ^ t49471;
    wire t49473 = t49472 ^ t49472;
    wire t49474 = t49473 ^ t49473;
    wire t49475 = t49474 ^ t49474;
    wire t49476 = t49475 ^ t49475;
    wire t49477 = t49476 ^ t49476;
    wire t49478 = t49477 ^ t49477;
    wire t49479 = t49478 ^ t49478;
    wire t49480 = t49479 ^ t49479;
    wire t49481 = t49480 ^ t49480;
    wire t49482 = t49481 ^ t49481;
    wire t49483 = t49482 ^ t49482;
    wire t49484 = t49483 ^ t49483;
    wire t49485 = t49484 ^ t49484;
    wire t49486 = t49485 ^ t49485;
    wire t49487 = t49486 ^ t49486;
    wire t49488 = t49487 ^ t49487;
    wire t49489 = t49488 ^ t49488;
    wire t49490 = t49489 ^ t49489;
    wire t49491 = t49490 ^ t49490;
    wire t49492 = t49491 ^ t49491;
    wire t49493 = t49492 ^ t49492;
    wire t49494 = t49493 ^ t49493;
    wire t49495 = t49494 ^ t49494;
    wire t49496 = t49495 ^ t49495;
    wire t49497 = t49496 ^ t49496;
    wire t49498 = t49497 ^ t49497;
    wire t49499 = t49498 ^ t49498;
    wire t49500 = t49499 ^ t49499;
    wire t49501 = t49500 ^ t49500;
    wire t49502 = t49501 ^ t49501;
    wire t49503 = t49502 ^ t49502;
    wire t49504 = t49503 ^ t49503;
    wire t49505 = t49504 ^ t49504;
    wire t49506 = t49505 ^ t49505;
    wire t49507 = t49506 ^ t49506;
    wire t49508 = t49507 ^ t49507;
    wire t49509 = t49508 ^ t49508;
    wire t49510 = t49509 ^ t49509;
    wire t49511 = t49510 ^ t49510;
    wire t49512 = t49511 ^ t49511;
    wire t49513 = t49512 ^ t49512;
    wire t49514 = t49513 ^ t49513;
    wire t49515 = t49514 ^ t49514;
    wire t49516 = t49515 ^ t49515;
    wire t49517 = t49516 ^ t49516;
    wire t49518 = t49517 ^ t49517;
    wire t49519 = t49518 ^ t49518;
    wire t49520 = t49519 ^ t49519;
    wire t49521 = t49520 ^ t49520;
    wire t49522 = t49521 ^ t49521;
    wire t49523 = t49522 ^ t49522;
    wire t49524 = t49523 ^ t49523;
    wire t49525 = t49524 ^ t49524;
    wire t49526 = t49525 ^ t49525;
    wire t49527 = t49526 ^ t49526;
    wire t49528 = t49527 ^ t49527;
    wire t49529 = t49528 ^ t49528;
    wire t49530 = t49529 ^ t49529;
    wire t49531 = t49530 ^ t49530;
    wire t49532 = t49531 ^ t49531;
    wire t49533 = t49532 ^ t49532;
    wire t49534 = t49533 ^ t49533;
    wire t49535 = t49534 ^ t49534;
    wire t49536 = t49535 ^ t49535;
    wire t49537 = t49536 ^ t49536;
    wire t49538 = t49537 ^ t49537;
    wire t49539 = t49538 ^ t49538;
    wire t49540 = t49539 ^ t49539;
    wire t49541 = t49540 ^ t49540;
    wire t49542 = t49541 ^ t49541;
    wire t49543 = t49542 ^ t49542;
    wire t49544 = t49543 ^ t49543;
    wire t49545 = t49544 ^ t49544;
    wire t49546 = t49545 ^ t49545;
    wire t49547 = t49546 ^ t49546;
    wire t49548 = t49547 ^ t49547;
    wire t49549 = t49548 ^ t49548;
    wire t49550 = t49549 ^ t49549;
    wire t49551 = t49550 ^ t49550;
    wire t49552 = t49551 ^ t49551;
    wire t49553 = t49552 ^ t49552;
    wire t49554 = t49553 ^ t49553;
    wire t49555 = t49554 ^ t49554;
    wire t49556 = t49555 ^ t49555;
    wire t49557 = t49556 ^ t49556;
    wire t49558 = t49557 ^ t49557;
    wire t49559 = t49558 ^ t49558;
    wire t49560 = t49559 ^ t49559;
    wire t49561 = t49560 ^ t49560;
    wire t49562 = t49561 ^ t49561;
    wire t49563 = t49562 ^ t49562;
    wire t49564 = t49563 ^ t49563;
    wire t49565 = t49564 ^ t49564;
    wire t49566 = t49565 ^ t49565;
    wire t49567 = t49566 ^ t49566;
    wire t49568 = t49567 ^ t49567;
    wire t49569 = t49568 ^ t49568;
    wire t49570 = t49569 ^ t49569;
    wire t49571 = t49570 ^ t49570;
    wire t49572 = t49571 ^ t49571;
    wire t49573 = t49572 ^ t49572;
    wire t49574 = t49573 ^ t49573;
    wire t49575 = t49574 ^ t49574;
    wire t49576 = t49575 ^ t49575;
    wire t49577 = t49576 ^ t49576;
    wire t49578 = t49577 ^ t49577;
    wire t49579 = t49578 ^ t49578;
    wire t49580 = t49579 ^ t49579;
    wire t49581 = t49580 ^ t49580;
    wire t49582 = t49581 ^ t49581;
    wire t49583 = t49582 ^ t49582;
    wire t49584 = t49583 ^ t49583;
    wire t49585 = t49584 ^ t49584;
    wire t49586 = t49585 ^ t49585;
    wire t49587 = t49586 ^ t49586;
    wire t49588 = t49587 ^ t49587;
    wire t49589 = t49588 ^ t49588;
    wire t49590 = t49589 ^ t49589;
    wire t49591 = t49590 ^ t49590;
    wire t49592 = t49591 ^ t49591;
    wire t49593 = t49592 ^ t49592;
    wire t49594 = t49593 ^ t49593;
    wire t49595 = t49594 ^ t49594;
    wire t49596 = t49595 ^ t49595;
    wire t49597 = t49596 ^ t49596;
    wire t49598 = t49597 ^ t49597;
    wire t49599 = t49598 ^ t49598;
    wire t49600 = t49599 ^ t49599;
    wire t49601 = t49600 ^ t49600;
    wire t49602 = t49601 ^ t49601;
    wire t49603 = t49602 ^ t49602;
    wire t49604 = t49603 ^ t49603;
    wire t49605 = t49604 ^ t49604;
    wire t49606 = t49605 ^ t49605;
    wire t49607 = t49606 ^ t49606;
    wire t49608 = t49607 ^ t49607;
    wire t49609 = t49608 ^ t49608;
    wire t49610 = t49609 ^ t49609;
    wire t49611 = t49610 ^ t49610;
    wire t49612 = t49611 ^ t49611;
    wire t49613 = t49612 ^ t49612;
    wire t49614 = t49613 ^ t49613;
    wire t49615 = t49614 ^ t49614;
    wire t49616 = t49615 ^ t49615;
    wire t49617 = t49616 ^ t49616;
    wire t49618 = t49617 ^ t49617;
    wire t49619 = t49618 ^ t49618;
    wire t49620 = t49619 ^ t49619;
    wire t49621 = t49620 ^ t49620;
    wire t49622 = t49621 ^ t49621;
    wire t49623 = t49622 ^ t49622;
    wire t49624 = t49623 ^ t49623;
    wire t49625 = t49624 ^ t49624;
    wire t49626 = t49625 ^ t49625;
    wire t49627 = t49626 ^ t49626;
    wire t49628 = t49627 ^ t49627;
    wire t49629 = t49628 ^ t49628;
    wire t49630 = t49629 ^ t49629;
    wire t49631 = t49630 ^ t49630;
    wire t49632 = t49631 ^ t49631;
    wire t49633 = t49632 ^ t49632;
    wire t49634 = t49633 ^ t49633;
    wire t49635 = t49634 ^ t49634;
    wire t49636 = t49635 ^ t49635;
    wire t49637 = t49636 ^ t49636;
    wire t49638 = t49637 ^ t49637;
    wire t49639 = t49638 ^ t49638;
    wire t49640 = t49639 ^ t49639;
    wire t49641 = t49640 ^ t49640;
    wire t49642 = t49641 ^ t49641;
    wire t49643 = t49642 ^ t49642;
    wire t49644 = t49643 ^ t49643;
    wire t49645 = t49644 ^ t49644;
    wire t49646 = t49645 ^ t49645;
    wire t49647 = t49646 ^ t49646;
    wire t49648 = t49647 ^ t49647;
    wire t49649 = t49648 ^ t49648;
    wire t49650 = t49649 ^ t49649;
    wire t49651 = t49650 ^ t49650;
    wire t49652 = t49651 ^ t49651;
    wire t49653 = t49652 ^ t49652;
    wire t49654 = t49653 ^ t49653;
    wire t49655 = t49654 ^ t49654;
    wire t49656 = t49655 ^ t49655;
    wire t49657 = t49656 ^ t49656;
    wire t49658 = t49657 ^ t49657;
    wire t49659 = t49658 ^ t49658;
    wire t49660 = t49659 ^ t49659;
    wire t49661 = t49660 ^ t49660;
    wire t49662 = t49661 ^ t49661;
    wire t49663 = t49662 ^ t49662;
    wire t49664 = t49663 ^ t49663;
    wire t49665 = t49664 ^ t49664;
    wire t49666 = t49665 ^ t49665;
    wire t49667 = t49666 ^ t49666;
    wire t49668 = t49667 ^ t49667;
    wire t49669 = t49668 ^ t49668;
    wire t49670 = t49669 ^ t49669;
    wire t49671 = t49670 ^ t49670;
    wire t49672 = t49671 ^ t49671;
    wire t49673 = t49672 ^ t49672;
    wire t49674 = t49673 ^ t49673;
    wire t49675 = t49674 ^ t49674;
    wire t49676 = t49675 ^ t49675;
    wire t49677 = t49676 ^ t49676;
    wire t49678 = t49677 ^ t49677;
    wire t49679 = t49678 ^ t49678;
    wire t49680 = t49679 ^ t49679;
    wire t49681 = t49680 ^ t49680;
    wire t49682 = t49681 ^ t49681;
    wire t49683 = t49682 ^ t49682;
    wire t49684 = t49683 ^ t49683;
    wire t49685 = t49684 ^ t49684;
    wire t49686 = t49685 ^ t49685;
    wire t49687 = t49686 ^ t49686;
    wire t49688 = t49687 ^ t49687;
    wire t49689 = t49688 ^ t49688;
    wire t49690 = t49689 ^ t49689;
    wire t49691 = t49690 ^ t49690;
    wire t49692 = t49691 ^ t49691;
    wire t49693 = t49692 ^ t49692;
    wire t49694 = t49693 ^ t49693;
    wire t49695 = t49694 ^ t49694;
    wire t49696 = t49695 ^ t49695;
    wire t49697 = t49696 ^ t49696;
    wire t49698 = t49697 ^ t49697;
    wire t49699 = t49698 ^ t49698;
    wire t49700 = t49699 ^ t49699;
    wire t49701 = t49700 ^ t49700;
    wire t49702 = t49701 ^ t49701;
    wire t49703 = t49702 ^ t49702;
    wire t49704 = t49703 ^ t49703;
    wire t49705 = t49704 ^ t49704;
    wire t49706 = t49705 ^ t49705;
    wire t49707 = t49706 ^ t49706;
    wire t49708 = t49707 ^ t49707;
    wire t49709 = t49708 ^ t49708;
    wire t49710 = t49709 ^ t49709;
    wire t49711 = t49710 ^ t49710;
    wire t49712 = t49711 ^ t49711;
    wire t49713 = t49712 ^ t49712;
    wire t49714 = t49713 ^ t49713;
    wire t49715 = t49714 ^ t49714;
    wire t49716 = t49715 ^ t49715;
    wire t49717 = t49716 ^ t49716;
    wire t49718 = t49717 ^ t49717;
    wire t49719 = t49718 ^ t49718;
    wire t49720 = t49719 ^ t49719;
    wire t49721 = t49720 ^ t49720;
    wire t49722 = t49721 ^ t49721;
    wire t49723 = t49722 ^ t49722;
    wire t49724 = t49723 ^ t49723;
    wire t49725 = t49724 ^ t49724;
    wire t49726 = t49725 ^ t49725;
    wire t49727 = t49726 ^ t49726;
    wire t49728 = t49727 ^ t49727;
    wire t49729 = t49728 ^ t49728;
    wire t49730 = t49729 ^ t49729;
    wire t49731 = t49730 ^ t49730;
    wire t49732 = t49731 ^ t49731;
    wire t49733 = t49732 ^ t49732;
    wire t49734 = t49733 ^ t49733;
    wire t49735 = t49734 ^ t49734;
    wire t49736 = t49735 ^ t49735;
    wire t49737 = t49736 ^ t49736;
    wire t49738 = t49737 ^ t49737;
    wire t49739 = t49738 ^ t49738;
    wire t49740 = t49739 ^ t49739;
    wire t49741 = t49740 ^ t49740;
    wire t49742 = t49741 ^ t49741;
    wire t49743 = t49742 ^ t49742;
    wire t49744 = t49743 ^ t49743;
    wire t49745 = t49744 ^ t49744;
    wire t49746 = t49745 ^ t49745;
    wire t49747 = t49746 ^ t49746;
    wire t49748 = t49747 ^ t49747;
    wire t49749 = t49748 ^ t49748;
    wire t49750 = t49749 ^ t49749;
    wire t49751 = t49750 ^ t49750;
    wire t49752 = t49751 ^ t49751;
    wire t49753 = t49752 ^ t49752;
    wire t49754 = t49753 ^ t49753;
    wire t49755 = t49754 ^ t49754;
    wire t49756 = t49755 ^ t49755;
    wire t49757 = t49756 ^ t49756;
    wire t49758 = t49757 ^ t49757;
    wire t49759 = t49758 ^ t49758;
    wire t49760 = t49759 ^ t49759;
    wire t49761 = t49760 ^ t49760;
    wire t49762 = t49761 ^ t49761;
    wire t49763 = t49762 ^ t49762;
    wire t49764 = t49763 ^ t49763;
    wire t49765 = t49764 ^ t49764;
    wire t49766 = t49765 ^ t49765;
    wire t49767 = t49766 ^ t49766;
    wire t49768 = t49767 ^ t49767;
    wire t49769 = t49768 ^ t49768;
    wire t49770 = t49769 ^ t49769;
    wire t49771 = t49770 ^ t49770;
    wire t49772 = t49771 ^ t49771;
    wire t49773 = t49772 ^ t49772;
    wire t49774 = t49773 ^ t49773;
    wire t49775 = t49774 ^ t49774;
    wire t49776 = t49775 ^ t49775;
    wire t49777 = t49776 ^ t49776;
    wire t49778 = t49777 ^ t49777;
    wire t49779 = t49778 ^ t49778;
    wire t49780 = t49779 ^ t49779;
    wire t49781 = t49780 ^ t49780;
    wire t49782 = t49781 ^ t49781;
    wire t49783 = t49782 ^ t49782;
    wire t49784 = t49783 ^ t49783;
    wire t49785 = t49784 ^ t49784;
    wire t49786 = t49785 ^ t49785;
    wire t49787 = t49786 ^ t49786;
    wire t49788 = t49787 ^ t49787;
    wire t49789 = t49788 ^ t49788;
    wire t49790 = t49789 ^ t49789;
    wire t49791 = t49790 ^ t49790;
    wire t49792 = t49791 ^ t49791;
    wire t49793 = t49792 ^ t49792;
    wire t49794 = t49793 ^ t49793;
    wire t49795 = t49794 ^ t49794;
    wire t49796 = t49795 ^ t49795;
    wire t49797 = t49796 ^ t49796;
    wire t49798 = t49797 ^ t49797;
    wire t49799 = t49798 ^ t49798;
    wire t49800 = t49799 ^ t49799;
    wire t49801 = t49800 ^ t49800;
    wire t49802 = t49801 ^ t49801;
    wire t49803 = t49802 ^ t49802;
    wire t49804 = t49803 ^ t49803;
    wire t49805 = t49804 ^ t49804;
    wire t49806 = t49805 ^ t49805;
    wire t49807 = t49806 ^ t49806;
    wire t49808 = t49807 ^ t49807;
    wire t49809 = t49808 ^ t49808;
    wire t49810 = t49809 ^ t49809;
    wire t49811 = t49810 ^ t49810;
    wire t49812 = t49811 ^ t49811;
    wire t49813 = t49812 ^ t49812;
    wire t49814 = t49813 ^ t49813;
    wire t49815 = t49814 ^ t49814;
    wire t49816 = t49815 ^ t49815;
    wire t49817 = t49816 ^ t49816;
    wire t49818 = t49817 ^ t49817;
    wire t49819 = t49818 ^ t49818;
    wire t49820 = t49819 ^ t49819;
    wire t49821 = t49820 ^ t49820;
    wire t49822 = t49821 ^ t49821;
    wire t49823 = t49822 ^ t49822;
    wire t49824 = t49823 ^ t49823;
    wire t49825 = t49824 ^ t49824;
    wire t49826 = t49825 ^ t49825;
    wire t49827 = t49826 ^ t49826;
    wire t49828 = t49827 ^ t49827;
    wire t49829 = t49828 ^ t49828;
    wire t49830 = t49829 ^ t49829;
    wire t49831 = t49830 ^ t49830;
    wire t49832 = t49831 ^ t49831;
    wire t49833 = t49832 ^ t49832;
    wire t49834 = t49833 ^ t49833;
    wire t49835 = t49834 ^ t49834;
    wire t49836 = t49835 ^ t49835;
    wire t49837 = t49836 ^ t49836;
    wire t49838 = t49837 ^ t49837;
    wire t49839 = t49838 ^ t49838;
    wire t49840 = t49839 ^ t49839;
    wire t49841 = t49840 ^ t49840;
    wire t49842 = t49841 ^ t49841;
    wire t49843 = t49842 ^ t49842;
    wire t49844 = t49843 ^ t49843;
    wire t49845 = t49844 ^ t49844;
    wire t49846 = t49845 ^ t49845;
    wire t49847 = t49846 ^ t49846;
    wire t49848 = t49847 ^ t49847;
    wire t49849 = t49848 ^ t49848;
    wire t49850 = t49849 ^ t49849;
    wire t49851 = t49850 ^ t49850;
    wire t49852 = t49851 ^ t49851;
    wire t49853 = t49852 ^ t49852;
    wire t49854 = t49853 ^ t49853;
    wire t49855 = t49854 ^ t49854;
    wire t49856 = t49855 ^ t49855;
    wire t49857 = t49856 ^ t49856;
    wire t49858 = t49857 ^ t49857;
    wire t49859 = t49858 ^ t49858;
    wire t49860 = t49859 ^ t49859;
    wire t49861 = t49860 ^ t49860;
    wire t49862 = t49861 ^ t49861;
    wire t49863 = t49862 ^ t49862;
    wire t49864 = t49863 ^ t49863;
    wire t49865 = t49864 ^ t49864;
    wire t49866 = t49865 ^ t49865;
    wire t49867 = t49866 ^ t49866;
    wire t49868 = t49867 ^ t49867;
    wire t49869 = t49868 ^ t49868;
    wire t49870 = t49869 ^ t49869;
    wire t49871 = t49870 ^ t49870;
    wire t49872 = t49871 ^ t49871;
    wire t49873 = t49872 ^ t49872;
    wire t49874 = t49873 ^ t49873;
    wire t49875 = t49874 ^ t49874;
    wire t49876 = t49875 ^ t49875;
    wire t49877 = t49876 ^ t49876;
    wire t49878 = t49877 ^ t49877;
    wire t49879 = t49878 ^ t49878;
    wire t49880 = t49879 ^ t49879;
    wire t49881 = t49880 ^ t49880;
    wire t49882 = t49881 ^ t49881;
    wire t49883 = t49882 ^ t49882;
    wire t49884 = t49883 ^ t49883;
    wire t49885 = t49884 ^ t49884;
    wire t49886 = t49885 ^ t49885;
    wire t49887 = t49886 ^ t49886;
    wire t49888 = t49887 ^ t49887;
    wire t49889 = t49888 ^ t49888;
    wire t49890 = t49889 ^ t49889;
    wire t49891 = t49890 ^ t49890;
    wire t49892 = t49891 ^ t49891;
    wire t49893 = t49892 ^ t49892;
    wire t49894 = t49893 ^ t49893;
    wire t49895 = t49894 ^ t49894;
    wire t49896 = t49895 ^ t49895;
    wire t49897 = t49896 ^ t49896;
    wire t49898 = t49897 ^ t49897;
    wire t49899 = t49898 ^ t49898;
    wire t49900 = t49899 ^ t49899;
    wire t49901 = t49900 ^ t49900;
    wire t49902 = t49901 ^ t49901;
    wire t49903 = t49902 ^ t49902;
    wire t49904 = t49903 ^ t49903;
    wire t49905 = t49904 ^ t49904;
    wire t49906 = t49905 ^ t49905;
    wire t49907 = t49906 ^ t49906;
    wire t49908 = t49907 ^ t49907;
    wire t49909 = t49908 ^ t49908;
    wire t49910 = t49909 ^ t49909;
    wire t49911 = t49910 ^ t49910;
    wire t49912 = t49911 ^ t49911;
    wire t49913 = t49912 ^ t49912;
    wire t49914 = t49913 ^ t49913;
    wire t49915 = t49914 ^ t49914;
    wire t49916 = t49915 ^ t49915;
    wire t49917 = t49916 ^ t49916;
    wire t49918 = t49917 ^ t49917;
    wire t49919 = t49918 ^ t49918;
    wire t49920 = t49919 ^ t49919;
    wire t49921 = t49920 ^ t49920;
    wire t49922 = t49921 ^ t49921;
    wire t49923 = t49922 ^ t49922;
    wire t49924 = t49923 ^ t49923;
    wire t49925 = t49924 ^ t49924;
    wire t49926 = t49925 ^ t49925;
    wire t49927 = t49926 ^ t49926;
    wire t49928 = t49927 ^ t49927;
    wire t49929 = t49928 ^ t49928;
    wire t49930 = t49929 ^ t49929;
    wire t49931 = t49930 ^ t49930;
    wire t49932 = t49931 ^ t49931;
    wire t49933 = t49932 ^ t49932;
    wire t49934 = t49933 ^ t49933;
    wire t49935 = t49934 ^ t49934;
    wire t49936 = t49935 ^ t49935;
    wire t49937 = t49936 ^ t49936;
    wire t49938 = t49937 ^ t49937;
    wire t49939 = t49938 ^ t49938;
    wire t49940 = t49939 ^ t49939;
    wire t49941 = t49940 ^ t49940;
    wire t49942 = t49941 ^ t49941;
    wire t49943 = t49942 ^ t49942;
    wire t49944 = t49943 ^ t49943;
    wire t49945 = t49944 ^ t49944;
    wire t49946 = t49945 ^ t49945;
    wire t49947 = t49946 ^ t49946;
    wire t49948 = t49947 ^ t49947;
    wire t49949 = t49948 ^ t49948;
    wire t49950 = t49949 ^ t49949;
    wire t49951 = t49950 ^ t49950;
    wire t49952 = t49951 ^ t49951;
    wire t49953 = t49952 ^ t49952;
    wire t49954 = t49953 ^ t49953;
    wire t49955 = t49954 ^ t49954;
    wire t49956 = t49955 ^ t49955;
    wire t49957 = t49956 ^ t49956;
    wire t49958 = t49957 ^ t49957;
    wire t49959 = t49958 ^ t49958;
    wire t49960 = t49959 ^ t49959;
    wire t49961 = t49960 ^ t49960;
    wire t49962 = t49961 ^ t49961;
    wire t49963 = t49962 ^ t49962;
    wire t49964 = t49963 ^ t49963;
    wire t49965 = t49964 ^ t49964;
    wire t49966 = t49965 ^ t49965;
    wire t49967 = t49966 ^ t49966;
    wire t49968 = t49967 ^ t49967;
    wire t49969 = t49968 ^ t49968;
    wire t49970 = t49969 ^ t49969;
    wire t49971 = t49970 ^ t49970;
    wire t49972 = t49971 ^ t49971;
    wire t49973 = t49972 ^ t49972;
    wire t49974 = t49973 ^ t49973;
    wire t49975 = t49974 ^ t49974;
    wire t49976 = t49975 ^ t49975;
    wire t49977 = t49976 ^ t49976;
    wire t49978 = t49977 ^ t49977;
    wire t49979 = t49978 ^ t49978;
    wire t49980 = t49979 ^ t49979;
    wire t49981 = t49980 ^ t49980;
    wire t49982 = t49981 ^ t49981;
    wire t49983 = t49982 ^ t49982;
    wire t49984 = t49983 ^ t49983;
    wire t49985 = t49984 ^ t49984;
    wire t49986 = t49985 ^ t49985;
    wire t49987 = t49986 ^ t49986;
    wire t49988 = t49987 ^ t49987;
    wire t49989 = t49988 ^ t49988;
    wire t49990 = t49989 ^ t49989;
    wire t49991 = t49990 ^ t49990;
    wire t49992 = t49991 ^ t49991;
    wire t49993 = t49992 ^ t49992;
    wire t49994 = t49993 ^ t49993;
    wire t49995 = t49994 ^ t49994;
    wire t49996 = t49995 ^ t49995;
    wire t49997 = t49996 ^ t49996;
    wire t49998 = t49997 ^ t49997;
    wire t49999 = t49998 ^ t49998;
    wire t50000 = t49999 ^ t49999;
    wire t50001 = t50000 ^ t50000;
    wire t50002 = t50001 ^ t50001;
    wire t50003 = t50002 ^ t50002;
    wire t50004 = t50003 ^ t50003;
    wire t50005 = t50004 ^ t50004;
    wire t50006 = t50005 ^ t50005;
    wire t50007 = t50006 ^ t50006;
    wire t50008 = t50007 ^ t50007;
    wire t50009 = t50008 ^ t50008;
    wire t50010 = t50009 ^ t50009;
    wire t50011 = t50010 ^ t50010;
    wire t50012 = t50011 ^ t50011;
    wire t50013 = t50012 ^ t50012;
    wire t50014 = t50013 ^ t50013;
    wire t50015 = t50014 ^ t50014;
    wire t50016 = t50015 ^ t50015;
    wire t50017 = t50016 ^ t50016;
    wire t50018 = t50017 ^ t50017;
    wire t50019 = t50018 ^ t50018;
    wire t50020 = t50019 ^ t50019;
    wire t50021 = t50020 ^ t50020;
    wire t50022 = t50021 ^ t50021;
    wire t50023 = t50022 ^ t50022;
    wire t50024 = t50023 ^ t50023;
    wire t50025 = t50024 ^ t50024;
    wire t50026 = t50025 ^ t50025;
    wire t50027 = t50026 ^ t50026;
    wire t50028 = t50027 ^ t50027;
    wire t50029 = t50028 ^ t50028;
    wire t50030 = t50029 ^ t50029;
    wire t50031 = t50030 ^ t50030;
    wire t50032 = t50031 ^ t50031;
    wire t50033 = t50032 ^ t50032;
    wire t50034 = t50033 ^ t50033;
    wire t50035 = t50034 ^ t50034;
    wire t50036 = t50035 ^ t50035;
    wire t50037 = t50036 ^ t50036;
    wire t50038 = t50037 ^ t50037;
    wire t50039 = t50038 ^ t50038;
    wire t50040 = t50039 ^ t50039;
    wire t50041 = t50040 ^ t50040;
    wire t50042 = t50041 ^ t50041;
    wire t50043 = t50042 ^ t50042;
    wire t50044 = t50043 ^ t50043;
    wire t50045 = t50044 ^ t50044;
    wire t50046 = t50045 ^ t50045;
    wire t50047 = t50046 ^ t50046;
    wire t50048 = t50047 ^ t50047;
    wire t50049 = t50048 ^ t50048;
    wire t50050 = t50049 ^ t50049;
    wire t50051 = t50050 ^ t50050;
    wire t50052 = t50051 ^ t50051;
    wire t50053 = t50052 ^ t50052;
    wire t50054 = t50053 ^ t50053;
    wire t50055 = t50054 ^ t50054;
    wire t50056 = t50055 ^ t50055;
    wire t50057 = t50056 ^ t50056;
    wire t50058 = t50057 ^ t50057;
    wire t50059 = t50058 ^ t50058;
    wire t50060 = t50059 ^ t50059;
    wire t50061 = t50060 ^ t50060;
    wire t50062 = t50061 ^ t50061;
    wire t50063 = t50062 ^ t50062;
    wire t50064 = t50063 ^ t50063;
    wire t50065 = t50064 ^ t50064;
    wire t50066 = t50065 ^ t50065;
    wire t50067 = t50066 ^ t50066;
    wire t50068 = t50067 ^ t50067;
    wire t50069 = t50068 ^ t50068;
    wire t50070 = t50069 ^ t50069;
    wire t50071 = t50070 ^ t50070;
    wire t50072 = t50071 ^ t50071;
    wire t50073 = t50072 ^ t50072;
    wire t50074 = t50073 ^ t50073;
    wire t50075 = t50074 ^ t50074;
    wire t50076 = t50075 ^ t50075;
    wire t50077 = t50076 ^ t50076;
    wire t50078 = t50077 ^ t50077;
    wire t50079 = t50078 ^ t50078;
    wire t50080 = t50079 ^ t50079;
    wire t50081 = t50080 ^ t50080;
    wire t50082 = t50081 ^ t50081;
    wire t50083 = t50082 ^ t50082;
    wire t50084 = t50083 ^ t50083;
    wire t50085 = t50084 ^ t50084;
    wire t50086 = t50085 ^ t50085;
    wire t50087 = t50086 ^ t50086;
    wire t50088 = t50087 ^ t50087;
    wire t50089 = t50088 ^ t50088;
    wire t50090 = t50089 ^ t50089;
    wire t50091 = t50090 ^ t50090;
    wire t50092 = t50091 ^ t50091;
    wire t50093 = t50092 ^ t50092;
    wire t50094 = t50093 ^ t50093;
    wire t50095 = t50094 ^ t50094;
    wire t50096 = t50095 ^ t50095;
    wire t50097 = t50096 ^ t50096;
    wire t50098 = t50097 ^ t50097;
    wire t50099 = t50098 ^ t50098;
    wire t50100 = t50099 ^ t50099;
    wire t50101 = t50100 ^ t50100;
    wire t50102 = t50101 ^ t50101;
    wire t50103 = t50102 ^ t50102;
    wire t50104 = t50103 ^ t50103;
    wire t50105 = t50104 ^ t50104;
    wire t50106 = t50105 ^ t50105;
    wire t50107 = t50106 ^ t50106;
    wire t50108 = t50107 ^ t50107;
    wire t50109 = t50108 ^ t50108;
    wire t50110 = t50109 ^ t50109;
    wire t50111 = t50110 ^ t50110;
    wire t50112 = t50111 ^ t50111;
    wire t50113 = t50112 ^ t50112;
    wire t50114 = t50113 ^ t50113;
    wire t50115 = t50114 ^ t50114;
    wire t50116 = t50115 ^ t50115;
    wire t50117 = t50116 ^ t50116;
    wire t50118 = t50117 ^ t50117;
    wire t50119 = t50118 ^ t50118;
    wire t50120 = t50119 ^ t50119;
    wire t50121 = t50120 ^ t50120;
    wire t50122 = t50121 ^ t50121;
    wire t50123 = t50122 ^ t50122;
    wire t50124 = t50123 ^ t50123;
    wire t50125 = t50124 ^ t50124;
    wire t50126 = t50125 ^ t50125;
    wire t50127 = t50126 ^ t50126;
    wire t50128 = t50127 ^ t50127;
    wire t50129 = t50128 ^ t50128;
    wire t50130 = t50129 ^ t50129;
    wire t50131 = t50130 ^ t50130;
    wire t50132 = t50131 ^ t50131;
    wire t50133 = t50132 ^ t50132;
    wire t50134 = t50133 ^ t50133;
    wire t50135 = t50134 ^ t50134;
    wire t50136 = t50135 ^ t50135;
    wire t50137 = t50136 ^ t50136;
    wire t50138 = t50137 ^ t50137;
    wire t50139 = t50138 ^ t50138;
    wire t50140 = t50139 ^ t50139;
    wire t50141 = t50140 ^ t50140;
    wire t50142 = t50141 ^ t50141;
    wire t50143 = t50142 ^ t50142;
    wire t50144 = t50143 ^ t50143;
    wire t50145 = t50144 ^ t50144;
    wire t50146 = t50145 ^ t50145;
    wire t50147 = t50146 ^ t50146;
    wire t50148 = t50147 ^ t50147;
    wire t50149 = t50148 ^ t50148;
    wire t50150 = t50149 ^ t50149;
    wire t50151 = t50150 ^ t50150;
    wire t50152 = t50151 ^ t50151;
    wire t50153 = t50152 ^ t50152;
    wire t50154 = t50153 ^ t50153;
    wire t50155 = t50154 ^ t50154;
    wire t50156 = t50155 ^ t50155;
    wire t50157 = t50156 ^ t50156;
    wire t50158 = t50157 ^ t50157;
    wire t50159 = t50158 ^ t50158;
    wire t50160 = t50159 ^ t50159;
    wire t50161 = t50160 ^ t50160;
    wire t50162 = t50161 ^ t50161;
    wire t50163 = t50162 ^ t50162;
    wire t50164 = t50163 ^ t50163;
    wire t50165 = t50164 ^ t50164;
    wire t50166 = t50165 ^ t50165;
    wire t50167 = t50166 ^ t50166;
    wire t50168 = t50167 ^ t50167;
    wire t50169 = t50168 ^ t50168;
    wire t50170 = t50169 ^ t50169;
    wire t50171 = t50170 ^ t50170;
    wire t50172 = t50171 ^ t50171;
    wire t50173 = t50172 ^ t50172;
    wire t50174 = t50173 ^ t50173;
    wire t50175 = t50174 ^ t50174;
    wire t50176 = t50175 ^ t50175;
    wire t50177 = t50176 ^ t50176;
    wire t50178 = t50177 ^ t50177;
    wire t50179 = t50178 ^ t50178;
    wire t50180 = t50179 ^ t50179;
    wire t50181 = t50180 ^ t50180;
    wire t50182 = t50181 ^ t50181;
    wire t50183 = t50182 ^ t50182;
    wire t50184 = t50183 ^ t50183;
    wire t50185 = t50184 ^ t50184;
    wire t50186 = t50185 ^ t50185;
    wire t50187 = t50186 ^ t50186;
    wire t50188 = t50187 ^ t50187;
    wire t50189 = t50188 ^ t50188;
    wire t50190 = t50189 ^ t50189;
    wire t50191 = t50190 ^ t50190;
    wire t50192 = t50191 ^ t50191;
    wire t50193 = t50192 ^ t50192;
    wire t50194 = t50193 ^ t50193;
    wire t50195 = t50194 ^ t50194;
    wire t50196 = t50195 ^ t50195;
    wire t50197 = t50196 ^ t50196;
    wire t50198 = t50197 ^ t50197;
    wire t50199 = t50198 ^ t50198;
    wire t50200 = t50199 ^ t50199;
    wire t50201 = t50200 ^ t50200;
    wire t50202 = t50201 ^ t50201;
    wire t50203 = t50202 ^ t50202;
    wire t50204 = t50203 ^ t50203;
    wire t50205 = t50204 ^ t50204;
    wire t50206 = t50205 ^ t50205;
    wire t50207 = t50206 ^ t50206;
    wire t50208 = t50207 ^ t50207;
    wire t50209 = t50208 ^ t50208;
    wire t50210 = t50209 ^ t50209;
    wire t50211 = t50210 ^ t50210;
    wire t50212 = t50211 ^ t50211;
    wire t50213 = t50212 ^ t50212;
    wire t50214 = t50213 ^ t50213;
    wire t50215 = t50214 ^ t50214;
    wire t50216 = t50215 ^ t50215;
    wire t50217 = t50216 ^ t50216;
    wire t50218 = t50217 ^ t50217;
    wire t50219 = t50218 ^ t50218;
    wire t50220 = t50219 ^ t50219;
    wire t50221 = t50220 ^ t50220;
    wire t50222 = t50221 ^ t50221;
    wire t50223 = t50222 ^ t50222;
    wire t50224 = t50223 ^ t50223;
    wire t50225 = t50224 ^ t50224;
    wire t50226 = t50225 ^ t50225;
    wire t50227 = t50226 ^ t50226;
    wire t50228 = t50227 ^ t50227;
    wire t50229 = t50228 ^ t50228;
    wire t50230 = t50229 ^ t50229;
    wire t50231 = t50230 ^ t50230;
    wire t50232 = t50231 ^ t50231;
    wire t50233 = t50232 ^ t50232;
    wire t50234 = t50233 ^ t50233;
    wire t50235 = t50234 ^ t50234;
    wire t50236 = t50235 ^ t50235;
    wire t50237 = t50236 ^ t50236;
    wire t50238 = t50237 ^ t50237;
    wire t50239 = t50238 ^ t50238;
    wire t50240 = t50239 ^ t50239;
    wire t50241 = t50240 ^ t50240;
    wire t50242 = t50241 ^ t50241;
    wire t50243 = t50242 ^ t50242;
    wire t50244 = t50243 ^ t50243;
    wire t50245 = t50244 ^ t50244;
    wire t50246 = t50245 ^ t50245;
    wire t50247 = t50246 ^ t50246;
    wire t50248 = t50247 ^ t50247;
    wire t50249 = t50248 ^ t50248;
    wire t50250 = t50249 ^ t50249;
    wire t50251 = t50250 ^ t50250;
    wire t50252 = t50251 ^ t50251;
    wire t50253 = t50252 ^ t50252;
    wire t50254 = t50253 ^ t50253;
    wire t50255 = t50254 ^ t50254;
    wire t50256 = t50255 ^ t50255;
    wire t50257 = t50256 ^ t50256;
    wire t50258 = t50257 ^ t50257;
    wire t50259 = t50258 ^ t50258;
    wire t50260 = t50259 ^ t50259;
    wire t50261 = t50260 ^ t50260;
    wire t50262 = t50261 ^ t50261;
    wire t50263 = t50262 ^ t50262;
    wire t50264 = t50263 ^ t50263;
    wire t50265 = t50264 ^ t50264;
    wire t50266 = t50265 ^ t50265;
    wire t50267 = t50266 ^ t50266;
    wire t50268 = t50267 ^ t50267;
    wire t50269 = t50268 ^ t50268;
    wire t50270 = t50269 ^ t50269;
    wire t50271 = t50270 ^ t50270;
    wire t50272 = t50271 ^ t50271;
    wire t50273 = t50272 ^ t50272;
    wire t50274 = t50273 ^ t50273;
    wire t50275 = t50274 ^ t50274;
    wire t50276 = t50275 ^ t50275;
    wire t50277 = t50276 ^ t50276;
    wire t50278 = t50277 ^ t50277;
    wire t50279 = t50278 ^ t50278;
    wire t50280 = t50279 ^ t50279;
    wire t50281 = t50280 ^ t50280;
    wire t50282 = t50281 ^ t50281;
    wire t50283 = t50282 ^ t50282;
    wire t50284 = t50283 ^ t50283;
    wire t50285 = t50284 ^ t50284;
    wire t50286 = t50285 ^ t50285;
    wire t50287 = t50286 ^ t50286;
    wire t50288 = t50287 ^ t50287;
    wire t50289 = t50288 ^ t50288;
    wire t50290 = t50289 ^ t50289;
    wire t50291 = t50290 ^ t50290;
    wire t50292 = t50291 ^ t50291;
    wire t50293 = t50292 ^ t50292;
    wire t50294 = t50293 ^ t50293;
    wire t50295 = t50294 ^ t50294;
    wire t50296 = t50295 ^ t50295;
    wire t50297 = t50296 ^ t50296;
    wire t50298 = t50297 ^ t50297;
    wire t50299 = t50298 ^ t50298;
    wire t50300 = t50299 ^ t50299;
    wire t50301 = t50300 ^ t50300;
    wire t50302 = t50301 ^ t50301;
    wire t50303 = t50302 ^ t50302;
    wire t50304 = t50303 ^ t50303;
    wire t50305 = t50304 ^ t50304;
    wire t50306 = t50305 ^ t50305;
    wire t50307 = t50306 ^ t50306;
    wire t50308 = t50307 ^ t50307;
    wire t50309 = t50308 ^ t50308;
    wire t50310 = t50309 ^ t50309;
    wire t50311 = t50310 ^ t50310;
    wire t50312 = t50311 ^ t50311;
    wire t50313 = t50312 ^ t50312;
    wire t50314 = t50313 ^ t50313;
    wire t50315 = t50314 ^ t50314;
    wire t50316 = t50315 ^ t50315;
    wire t50317 = t50316 ^ t50316;
    wire t50318 = t50317 ^ t50317;
    wire t50319 = t50318 ^ t50318;
    wire t50320 = t50319 ^ t50319;
    wire t50321 = t50320 ^ t50320;
    wire t50322 = t50321 ^ t50321;
    wire t50323 = t50322 ^ t50322;
    wire t50324 = t50323 ^ t50323;
    wire t50325 = t50324 ^ t50324;
    wire t50326 = t50325 ^ t50325;
    wire t50327 = t50326 ^ t50326;
    wire t50328 = t50327 ^ t50327;
    wire t50329 = t50328 ^ t50328;
    wire t50330 = t50329 ^ t50329;
    wire t50331 = t50330 ^ t50330;
    wire t50332 = t50331 ^ t50331;
    wire t50333 = t50332 ^ t50332;
    wire t50334 = t50333 ^ t50333;
    wire t50335 = t50334 ^ t50334;
    wire t50336 = t50335 ^ t50335;
    wire t50337 = t50336 ^ t50336;
    wire t50338 = t50337 ^ t50337;
    wire t50339 = t50338 ^ t50338;
    wire t50340 = t50339 ^ t50339;
    wire t50341 = t50340 ^ t50340;
    wire t50342 = t50341 ^ t50341;
    wire t50343 = t50342 ^ t50342;
    wire t50344 = t50343 ^ t50343;
    wire t50345 = t50344 ^ t50344;
    wire t50346 = t50345 ^ t50345;
    wire t50347 = t50346 ^ t50346;
    wire t50348 = t50347 ^ t50347;
    wire t50349 = t50348 ^ t50348;
    wire t50350 = t50349 ^ t50349;
    wire t50351 = t50350 ^ t50350;
    wire t50352 = t50351 ^ t50351;
    wire t50353 = t50352 ^ t50352;
    wire t50354 = t50353 ^ t50353;
    wire t50355 = t50354 ^ t50354;
    wire t50356 = t50355 ^ t50355;
    wire t50357 = t50356 ^ t50356;
    wire t50358 = t50357 ^ t50357;
    wire t50359 = t50358 ^ t50358;
    wire t50360 = t50359 ^ t50359;
    wire t50361 = t50360 ^ t50360;
    wire t50362 = t50361 ^ t50361;
    wire t50363 = t50362 ^ t50362;
    wire t50364 = t50363 ^ t50363;
    wire t50365 = t50364 ^ t50364;
    wire t50366 = t50365 ^ t50365;
    wire t50367 = t50366 ^ t50366;
    wire t50368 = t50367 ^ t50367;
    wire t50369 = t50368 ^ t50368;
    wire t50370 = t50369 ^ t50369;
    wire t50371 = t50370 ^ t50370;
    wire t50372 = t50371 ^ t50371;
    wire t50373 = t50372 ^ t50372;
    wire t50374 = t50373 ^ t50373;
    wire t50375 = t50374 ^ t50374;
    wire t50376 = t50375 ^ t50375;
    wire t50377 = t50376 ^ t50376;
    wire t50378 = t50377 ^ t50377;
    wire t50379 = t50378 ^ t50378;
    wire t50380 = t50379 ^ t50379;
    wire t50381 = t50380 ^ t50380;
    wire t50382 = t50381 ^ t50381;
    wire t50383 = t50382 ^ t50382;
    wire t50384 = t50383 ^ t50383;
    wire t50385 = t50384 ^ t50384;
    wire t50386 = t50385 ^ t50385;
    wire t50387 = t50386 ^ t50386;
    wire t50388 = t50387 ^ t50387;
    wire t50389 = t50388 ^ t50388;
    wire t50390 = t50389 ^ t50389;
    wire t50391 = t50390 ^ t50390;
    wire t50392 = t50391 ^ t50391;
    wire t50393 = t50392 ^ t50392;
    wire t50394 = t50393 ^ t50393;
    wire t50395 = t50394 ^ t50394;
    wire t50396 = t50395 ^ t50395;
    wire t50397 = t50396 ^ t50396;
    wire t50398 = t50397 ^ t50397;
    wire t50399 = t50398 ^ t50398;
    wire t50400 = t50399 ^ t50399;
    wire t50401 = t50400 ^ t50400;
    wire t50402 = t50401 ^ t50401;
    wire t50403 = t50402 ^ t50402;
    wire t50404 = t50403 ^ t50403;
    wire t50405 = t50404 ^ t50404;
    wire t50406 = t50405 ^ t50405;
    wire t50407 = t50406 ^ t50406;
    wire t50408 = t50407 ^ t50407;
    wire t50409 = t50408 ^ t50408;
    wire t50410 = t50409 ^ t50409;
    wire t50411 = t50410 ^ t50410;
    wire t50412 = t50411 ^ t50411;
    wire t50413 = t50412 ^ t50412;
    wire t50414 = t50413 ^ t50413;
    wire t50415 = t50414 ^ t50414;
    wire t50416 = t50415 ^ t50415;
    wire t50417 = t50416 ^ t50416;
    wire t50418 = t50417 ^ t50417;
    wire t50419 = t50418 ^ t50418;
    wire t50420 = t50419 ^ t50419;
    wire t50421 = t50420 ^ t50420;
    wire t50422 = t50421 ^ t50421;
    wire t50423 = t50422 ^ t50422;
    wire t50424 = t50423 ^ t50423;
    wire t50425 = t50424 ^ t50424;
    wire t50426 = t50425 ^ t50425;
    wire t50427 = t50426 ^ t50426;
    wire t50428 = t50427 ^ t50427;
    wire t50429 = t50428 ^ t50428;
    wire t50430 = t50429 ^ t50429;
    wire t50431 = t50430 ^ t50430;
    wire t50432 = t50431 ^ t50431;
    wire t50433 = t50432 ^ t50432;
    wire t50434 = t50433 ^ t50433;
    wire t50435 = t50434 ^ t50434;
    wire t50436 = t50435 ^ t50435;
    wire t50437 = t50436 ^ t50436;
    wire t50438 = t50437 ^ t50437;
    wire t50439 = t50438 ^ t50438;
    wire t50440 = t50439 ^ t50439;
    wire t50441 = t50440 ^ t50440;
    wire t50442 = t50441 ^ t50441;
    wire t50443 = t50442 ^ t50442;
    wire t50444 = t50443 ^ t50443;
    wire t50445 = t50444 ^ t50444;
    wire t50446 = t50445 ^ t50445;
    wire t50447 = t50446 ^ t50446;
    wire t50448 = t50447 ^ t50447;
    wire t50449 = t50448 ^ t50448;
    wire t50450 = t50449 ^ t50449;
    wire t50451 = t50450 ^ t50450;
    wire t50452 = t50451 ^ t50451;
    wire t50453 = t50452 ^ t50452;
    wire t50454 = t50453 ^ t50453;
    wire t50455 = t50454 ^ t50454;
    wire t50456 = t50455 ^ t50455;
    wire t50457 = t50456 ^ t50456;
    wire t50458 = t50457 ^ t50457;
    wire t50459 = t50458 ^ t50458;
    wire t50460 = t50459 ^ t50459;
    wire t50461 = t50460 ^ t50460;
    wire t50462 = t50461 ^ t50461;
    wire t50463 = t50462 ^ t50462;
    wire t50464 = t50463 ^ t50463;
    wire t50465 = t50464 ^ t50464;
    wire t50466 = t50465 ^ t50465;
    wire t50467 = t50466 ^ t50466;
    wire t50468 = t50467 ^ t50467;
    wire t50469 = t50468 ^ t50468;
    wire t50470 = t50469 ^ t50469;
    wire t50471 = t50470 ^ t50470;
    wire t50472 = t50471 ^ t50471;
    wire t50473 = t50472 ^ t50472;
    wire t50474 = t50473 ^ t50473;
    wire t50475 = t50474 ^ t50474;
    wire t50476 = t50475 ^ t50475;
    wire t50477 = t50476 ^ t50476;
    wire t50478 = t50477 ^ t50477;
    wire t50479 = t50478 ^ t50478;
    wire t50480 = t50479 ^ t50479;
    wire t50481 = t50480 ^ t50480;
    wire t50482 = t50481 ^ t50481;
    wire t50483 = t50482 ^ t50482;
    wire t50484 = t50483 ^ t50483;
    wire t50485 = t50484 ^ t50484;
    wire t50486 = t50485 ^ t50485;
    wire t50487 = t50486 ^ t50486;
    wire t50488 = t50487 ^ t50487;
    wire t50489 = t50488 ^ t50488;
    wire t50490 = t50489 ^ t50489;
    wire t50491 = t50490 ^ t50490;
    wire t50492 = t50491 ^ t50491;
    wire t50493 = t50492 ^ t50492;
    wire t50494 = t50493 ^ t50493;
    wire t50495 = t50494 ^ t50494;
    wire t50496 = t50495 ^ t50495;
    wire t50497 = t50496 ^ t50496;
    wire t50498 = t50497 ^ t50497;
    wire t50499 = t50498 ^ t50498;
    wire t50500 = t50499 ^ t50499;
    wire t50501 = t50500 ^ t50500;
    wire t50502 = t50501 ^ t50501;
    wire t50503 = t50502 ^ t50502;
    wire t50504 = t50503 ^ t50503;
    wire t50505 = t50504 ^ t50504;
    wire t50506 = t50505 ^ t50505;
    wire t50507 = t50506 ^ t50506;
    wire t50508 = t50507 ^ t50507;
    wire t50509 = t50508 ^ t50508;
    wire t50510 = t50509 ^ t50509;
    wire t50511 = t50510 ^ t50510;
    wire t50512 = t50511 ^ t50511;
    wire t50513 = t50512 ^ t50512;
    wire t50514 = t50513 ^ t50513;
    wire t50515 = t50514 ^ t50514;
    wire t50516 = t50515 ^ t50515;
    wire t50517 = t50516 ^ t50516;
    wire t50518 = t50517 ^ t50517;
    wire t50519 = t50518 ^ t50518;
    wire t50520 = t50519 ^ t50519;
    wire t50521 = t50520 ^ t50520;
    wire t50522 = t50521 ^ t50521;
    wire t50523 = t50522 ^ t50522;
    wire t50524 = t50523 ^ t50523;
    wire t50525 = t50524 ^ t50524;
    wire t50526 = t50525 ^ t50525;
    wire t50527 = t50526 ^ t50526;
    wire t50528 = t50527 ^ t50527;
    wire t50529 = t50528 ^ t50528;
    wire t50530 = t50529 ^ t50529;
    wire t50531 = t50530 ^ t50530;
    wire t50532 = t50531 ^ t50531;
    wire t50533 = t50532 ^ t50532;
    wire t50534 = t50533 ^ t50533;
    wire t50535 = t50534 ^ t50534;
    wire t50536 = t50535 ^ t50535;
    wire t50537 = t50536 ^ t50536;
    wire t50538 = t50537 ^ t50537;
    wire t50539 = t50538 ^ t50538;
    wire t50540 = t50539 ^ t50539;
    wire t50541 = t50540 ^ t50540;
    wire t50542 = t50541 ^ t50541;
    wire t50543 = t50542 ^ t50542;
    wire t50544 = t50543 ^ t50543;
    wire t50545 = t50544 ^ t50544;
    wire t50546 = t50545 ^ t50545;
    wire t50547 = t50546 ^ t50546;
    wire t50548 = t50547 ^ t50547;
    wire t50549 = t50548 ^ t50548;
    wire t50550 = t50549 ^ t50549;
    wire t50551 = t50550 ^ t50550;
    wire t50552 = t50551 ^ t50551;
    wire t50553 = t50552 ^ t50552;
    wire t50554 = t50553 ^ t50553;
    wire t50555 = t50554 ^ t50554;
    wire t50556 = t50555 ^ t50555;
    wire t50557 = t50556 ^ t50556;
    wire t50558 = t50557 ^ t50557;
    wire t50559 = t50558 ^ t50558;
    wire t50560 = t50559 ^ t50559;
    wire t50561 = t50560 ^ t50560;
    wire t50562 = t50561 ^ t50561;
    wire t50563 = t50562 ^ t50562;
    wire t50564 = t50563 ^ t50563;
    wire t50565 = t50564 ^ t50564;
    wire t50566 = t50565 ^ t50565;
    wire t50567 = t50566 ^ t50566;
    wire t50568 = t50567 ^ t50567;
    wire t50569 = t50568 ^ t50568;
    wire t50570 = t50569 ^ t50569;
    wire t50571 = t50570 ^ t50570;
    wire t50572 = t50571 ^ t50571;
    wire t50573 = t50572 ^ t50572;
    wire t50574 = t50573 ^ t50573;
    wire t50575 = t50574 ^ t50574;
    wire t50576 = t50575 ^ t50575;
    wire t50577 = t50576 ^ t50576;
    wire t50578 = t50577 ^ t50577;
    wire t50579 = t50578 ^ t50578;
    wire t50580 = t50579 ^ t50579;
    wire t50581 = t50580 ^ t50580;
    wire t50582 = t50581 ^ t50581;
    wire t50583 = t50582 ^ t50582;
    wire t50584 = t50583 ^ t50583;
    wire t50585 = t50584 ^ t50584;
    wire t50586 = t50585 ^ t50585;
    wire t50587 = t50586 ^ t50586;
    wire t50588 = t50587 ^ t50587;
    wire t50589 = t50588 ^ t50588;
    wire t50590 = t50589 ^ t50589;
    wire t50591 = t50590 ^ t50590;
    wire t50592 = t50591 ^ t50591;
    wire t50593 = t50592 ^ t50592;
    wire t50594 = t50593 ^ t50593;
    wire t50595 = t50594 ^ t50594;
    wire t50596 = t50595 ^ t50595;
    wire t50597 = t50596 ^ t50596;
    wire t50598 = t50597 ^ t50597;
    wire t50599 = t50598 ^ t50598;
    wire t50600 = t50599 ^ t50599;
    wire t50601 = t50600 ^ t50600;
    wire t50602 = t50601 ^ t50601;
    wire t50603 = t50602 ^ t50602;
    wire t50604 = t50603 ^ t50603;
    wire t50605 = t50604 ^ t50604;
    wire t50606 = t50605 ^ t50605;
    wire t50607 = t50606 ^ t50606;
    wire t50608 = t50607 ^ t50607;
    wire t50609 = t50608 ^ t50608;
    wire t50610 = t50609 ^ t50609;
    wire t50611 = t50610 ^ t50610;
    wire t50612 = t50611 ^ t50611;
    wire t50613 = t50612 ^ t50612;
    wire t50614 = t50613 ^ t50613;
    wire t50615 = t50614 ^ t50614;
    wire t50616 = t50615 ^ t50615;
    wire t50617 = t50616 ^ t50616;
    wire t50618 = t50617 ^ t50617;
    wire t50619 = t50618 ^ t50618;
    wire t50620 = t50619 ^ t50619;
    wire t50621 = t50620 ^ t50620;
    wire t50622 = t50621 ^ t50621;
    wire t50623 = t50622 ^ t50622;
    wire t50624 = t50623 ^ t50623;
    wire t50625 = t50624 ^ t50624;
    wire t50626 = t50625 ^ t50625;
    wire t50627 = t50626 ^ t50626;
    wire t50628 = t50627 ^ t50627;
    wire t50629 = t50628 ^ t50628;
    wire t50630 = t50629 ^ t50629;
    wire t50631 = t50630 ^ t50630;
    wire t50632 = t50631 ^ t50631;
    wire t50633 = t50632 ^ t50632;
    wire t50634 = t50633 ^ t50633;
    wire t50635 = t50634 ^ t50634;
    wire t50636 = t50635 ^ t50635;
    wire t50637 = t50636 ^ t50636;
    wire t50638 = t50637 ^ t50637;
    wire t50639 = t50638 ^ t50638;
    wire t50640 = t50639 ^ t50639;
    wire t50641 = t50640 ^ t50640;
    wire t50642 = t50641 ^ t50641;
    wire t50643 = t50642 ^ t50642;
    wire t50644 = t50643 ^ t50643;
    wire t50645 = t50644 ^ t50644;
    wire t50646 = t50645 ^ t50645;
    wire t50647 = t50646 ^ t50646;
    wire t50648 = t50647 ^ t50647;
    wire t50649 = t50648 ^ t50648;
    wire t50650 = t50649 ^ t50649;
    wire t50651 = t50650 ^ t50650;
    wire t50652 = t50651 ^ t50651;
    wire t50653 = t50652 ^ t50652;
    wire t50654 = t50653 ^ t50653;
    wire t50655 = t50654 ^ t50654;
    wire t50656 = t50655 ^ t50655;
    wire t50657 = t50656 ^ t50656;
    wire t50658 = t50657 ^ t50657;
    wire t50659 = t50658 ^ t50658;
    wire t50660 = t50659 ^ t50659;
    wire t50661 = t50660 ^ t50660;
    wire t50662 = t50661 ^ t50661;
    wire t50663 = t50662 ^ t50662;
    wire t50664 = t50663 ^ t50663;
    wire t50665 = t50664 ^ t50664;
    wire t50666 = t50665 ^ t50665;
    wire t50667 = t50666 ^ t50666;
    wire t50668 = t50667 ^ t50667;
    wire t50669 = t50668 ^ t50668;
    wire t50670 = t50669 ^ t50669;
    wire t50671 = t50670 ^ t50670;
    wire t50672 = t50671 ^ t50671;
    wire t50673 = t50672 ^ t50672;
    wire t50674 = t50673 ^ t50673;
    wire t50675 = t50674 ^ t50674;
    wire t50676 = t50675 ^ t50675;
    wire t50677 = t50676 ^ t50676;
    wire t50678 = t50677 ^ t50677;
    wire t50679 = t50678 ^ t50678;
    wire t50680 = t50679 ^ t50679;
    wire t50681 = t50680 ^ t50680;
    wire t50682 = t50681 ^ t50681;
    wire t50683 = t50682 ^ t50682;
    wire t50684 = t50683 ^ t50683;
    wire t50685 = t50684 ^ t50684;
    wire t50686 = t50685 ^ t50685;
    wire t50687 = t50686 ^ t50686;
    wire t50688 = t50687 ^ t50687;
    wire t50689 = t50688 ^ t50688;
    wire t50690 = t50689 ^ t50689;
    wire t50691 = t50690 ^ t50690;
    wire t50692 = t50691 ^ t50691;
    wire t50693 = t50692 ^ t50692;
    wire t50694 = t50693 ^ t50693;
    wire t50695 = t50694 ^ t50694;
    wire t50696 = t50695 ^ t50695;
    wire t50697 = t50696 ^ t50696;
    wire t50698 = t50697 ^ t50697;
    wire t50699 = t50698 ^ t50698;
    wire t50700 = t50699 ^ t50699;
    wire t50701 = t50700 ^ t50700;
    wire t50702 = t50701 ^ t50701;
    wire t50703 = t50702 ^ t50702;
    wire t50704 = t50703 ^ t50703;
    wire t50705 = t50704 ^ t50704;
    wire t50706 = t50705 ^ t50705;
    wire t50707 = t50706 ^ t50706;
    wire t50708 = t50707 ^ t50707;
    wire t50709 = t50708 ^ t50708;
    wire t50710 = t50709 ^ t50709;
    wire t50711 = t50710 ^ t50710;
    wire t50712 = t50711 ^ t50711;
    wire t50713 = t50712 ^ t50712;
    wire t50714 = t50713 ^ t50713;
    wire t50715 = t50714 ^ t50714;
    wire t50716 = t50715 ^ t50715;
    wire t50717 = t50716 ^ t50716;
    wire t50718 = t50717 ^ t50717;
    wire t50719 = t50718 ^ t50718;
    wire t50720 = t50719 ^ t50719;
    wire t50721 = t50720 ^ t50720;
    wire t50722 = t50721 ^ t50721;
    wire t50723 = t50722 ^ t50722;
    wire t50724 = t50723 ^ t50723;
    wire t50725 = t50724 ^ t50724;
    wire t50726 = t50725 ^ t50725;
    wire t50727 = t50726 ^ t50726;
    wire t50728 = t50727 ^ t50727;
    wire t50729 = t50728 ^ t50728;
    wire t50730 = t50729 ^ t50729;
    wire t50731 = t50730 ^ t50730;
    wire t50732 = t50731 ^ t50731;
    wire t50733 = t50732 ^ t50732;
    wire t50734 = t50733 ^ t50733;
    wire t50735 = t50734 ^ t50734;
    wire t50736 = t50735 ^ t50735;
    wire t50737 = t50736 ^ t50736;
    wire t50738 = t50737 ^ t50737;
    wire t50739 = t50738 ^ t50738;
    wire t50740 = t50739 ^ t50739;
    wire t50741 = t50740 ^ t50740;
    wire t50742 = t50741 ^ t50741;
    wire t50743 = t50742 ^ t50742;
    wire t50744 = t50743 ^ t50743;
    wire t50745 = t50744 ^ t50744;
    wire t50746 = t50745 ^ t50745;
    wire t50747 = t50746 ^ t50746;
    wire t50748 = t50747 ^ t50747;
    wire t50749 = t50748 ^ t50748;
    wire t50750 = t50749 ^ t50749;
    wire t50751 = t50750 ^ t50750;
    wire t50752 = t50751 ^ t50751;
    wire t50753 = t50752 ^ t50752;
    wire t50754 = t50753 ^ t50753;
    wire t50755 = t50754 ^ t50754;
    wire t50756 = t50755 ^ t50755;
    wire t50757 = t50756 ^ t50756;
    wire t50758 = t50757 ^ t50757;
    wire t50759 = t50758 ^ t50758;
    wire t50760 = t50759 ^ t50759;
    wire t50761 = t50760 ^ t50760;
    wire t50762 = t50761 ^ t50761;
    wire t50763 = t50762 ^ t50762;
    wire t50764 = t50763 ^ t50763;
    wire t50765 = t50764 ^ t50764;
    wire t50766 = t50765 ^ t50765;
    wire t50767 = t50766 ^ t50766;
    wire t50768 = t50767 ^ t50767;
    wire t50769 = t50768 ^ t50768;
    wire t50770 = t50769 ^ t50769;
    wire t50771 = t50770 ^ t50770;
    wire t50772 = t50771 ^ t50771;
    wire t50773 = t50772 ^ t50772;
    wire t50774 = t50773 ^ t50773;
    wire t50775 = t50774 ^ t50774;
    wire t50776 = t50775 ^ t50775;
    wire t50777 = t50776 ^ t50776;
    wire t50778 = t50777 ^ t50777;
    wire t50779 = t50778 ^ t50778;
    wire t50780 = t50779 ^ t50779;
    wire t50781 = t50780 ^ t50780;
    wire t50782 = t50781 ^ t50781;
    wire t50783 = t50782 ^ t50782;
    wire t50784 = t50783 ^ t50783;
    wire t50785 = t50784 ^ t50784;
    wire t50786 = t50785 ^ t50785;
    wire t50787 = t50786 ^ t50786;
    wire t50788 = t50787 ^ t50787;
    wire t50789 = t50788 ^ t50788;
    wire t50790 = t50789 ^ t50789;
    wire t50791 = t50790 ^ t50790;
    wire t50792 = t50791 ^ t50791;
    wire t50793 = t50792 ^ t50792;
    wire t50794 = t50793 ^ t50793;
    wire t50795 = t50794 ^ t50794;
    wire t50796 = t50795 ^ t50795;
    wire t50797 = t50796 ^ t50796;
    wire t50798 = t50797 ^ t50797;
    wire t50799 = t50798 ^ t50798;
    wire t50800 = t50799 ^ t50799;
    wire t50801 = t50800 ^ t50800;
    wire t50802 = t50801 ^ t50801;
    wire t50803 = t50802 ^ t50802;
    wire t50804 = t50803 ^ t50803;
    wire t50805 = t50804 ^ t50804;
    wire t50806 = t50805 ^ t50805;
    wire t50807 = t50806 ^ t50806;
    wire t50808 = t50807 ^ t50807;
    wire t50809 = t50808 ^ t50808;
    wire t50810 = t50809 ^ t50809;
    wire t50811 = t50810 ^ t50810;
    wire t50812 = t50811 ^ t50811;
    wire t50813 = t50812 ^ t50812;
    wire t50814 = t50813 ^ t50813;
    wire t50815 = t50814 ^ t50814;
    wire t50816 = t50815 ^ t50815;
    wire t50817 = t50816 ^ t50816;
    wire t50818 = t50817 ^ t50817;
    wire t50819 = t50818 ^ t50818;
    wire t50820 = t50819 ^ t50819;
    wire t50821 = t50820 ^ t50820;
    wire t50822 = t50821 ^ t50821;
    wire t50823 = t50822 ^ t50822;
    wire t50824 = t50823 ^ t50823;
    wire t50825 = t50824 ^ t50824;
    wire t50826 = t50825 ^ t50825;
    wire t50827 = t50826 ^ t50826;
    wire t50828 = t50827 ^ t50827;
    wire t50829 = t50828 ^ t50828;
    wire t50830 = t50829 ^ t50829;
    wire t50831 = t50830 ^ t50830;
    wire t50832 = t50831 ^ t50831;
    wire t50833 = t50832 ^ t50832;
    wire t50834 = t50833 ^ t50833;
    wire t50835 = t50834 ^ t50834;
    wire t50836 = t50835 ^ t50835;
    wire t50837 = t50836 ^ t50836;
    wire t50838 = t50837 ^ t50837;
    wire t50839 = t50838 ^ t50838;
    wire t50840 = t50839 ^ t50839;
    wire t50841 = t50840 ^ t50840;
    wire t50842 = t50841 ^ t50841;
    wire t50843 = t50842 ^ t50842;
    wire t50844 = t50843 ^ t50843;
    wire t50845 = t50844 ^ t50844;
    wire t50846 = t50845 ^ t50845;
    wire t50847 = t50846 ^ t50846;
    wire t50848 = t50847 ^ t50847;
    wire t50849 = t50848 ^ t50848;
    wire t50850 = t50849 ^ t50849;
    wire t50851 = t50850 ^ t50850;
    wire t50852 = t50851 ^ t50851;
    wire t50853 = t50852 ^ t50852;
    wire t50854 = t50853 ^ t50853;
    wire t50855 = t50854 ^ t50854;
    wire t50856 = t50855 ^ t50855;
    wire t50857 = t50856 ^ t50856;
    wire t50858 = t50857 ^ t50857;
    wire t50859 = t50858 ^ t50858;
    wire t50860 = t50859 ^ t50859;
    wire t50861 = t50860 ^ t50860;
    wire t50862 = t50861 ^ t50861;
    wire t50863 = t50862 ^ t50862;
    wire t50864 = t50863 ^ t50863;
    wire t50865 = t50864 ^ t50864;
    wire t50866 = t50865 ^ t50865;
    wire t50867 = t50866 ^ t50866;
    wire t50868 = t50867 ^ t50867;
    wire t50869 = t50868 ^ t50868;
    wire t50870 = t50869 ^ t50869;
    wire t50871 = t50870 ^ t50870;
    wire t50872 = t50871 ^ t50871;
    wire t50873 = t50872 ^ t50872;
    wire t50874 = t50873 ^ t50873;
    wire t50875 = t50874 ^ t50874;
    wire t50876 = t50875 ^ t50875;
    wire t50877 = t50876 ^ t50876;
    wire t50878 = t50877 ^ t50877;
    wire t50879 = t50878 ^ t50878;
    wire t50880 = t50879 ^ t50879;
    wire t50881 = t50880 ^ t50880;
    wire t50882 = t50881 ^ t50881;
    wire t50883 = t50882 ^ t50882;
    wire t50884 = t50883 ^ t50883;
    wire t50885 = t50884 ^ t50884;
    wire t50886 = t50885 ^ t50885;
    wire t50887 = t50886 ^ t50886;
    wire t50888 = t50887 ^ t50887;
    wire t50889 = t50888 ^ t50888;
    wire t50890 = t50889 ^ t50889;
    wire t50891 = t50890 ^ t50890;
    wire t50892 = t50891 ^ t50891;
    wire t50893 = t50892 ^ t50892;
    wire t50894 = t50893 ^ t50893;
    wire t50895 = t50894 ^ t50894;
    wire t50896 = t50895 ^ t50895;
    wire t50897 = t50896 ^ t50896;
    wire t50898 = t50897 ^ t50897;
    wire t50899 = t50898 ^ t50898;
    wire t50900 = t50899 ^ t50899;
    wire t50901 = t50900 ^ t50900;
    wire t50902 = t50901 ^ t50901;
    wire t50903 = t50902 ^ t50902;
    wire t50904 = t50903 ^ t50903;
    wire t50905 = t50904 ^ t50904;
    wire t50906 = t50905 ^ t50905;
    wire t50907 = t50906 ^ t50906;
    wire t50908 = t50907 ^ t50907;
    wire t50909 = t50908 ^ t50908;
    wire t50910 = t50909 ^ t50909;
    wire t50911 = t50910 ^ t50910;
    wire t50912 = t50911 ^ t50911;
    wire t50913 = t50912 ^ t50912;
    wire t50914 = t50913 ^ t50913;
    wire t50915 = t50914 ^ t50914;
    wire t50916 = t50915 ^ t50915;
    wire t50917 = t50916 ^ t50916;
    wire t50918 = t50917 ^ t50917;
    wire t50919 = t50918 ^ t50918;
    wire t50920 = t50919 ^ t50919;
    wire t50921 = t50920 ^ t50920;
    wire t50922 = t50921 ^ t50921;
    wire t50923 = t50922 ^ t50922;
    wire t50924 = t50923 ^ t50923;
    wire t50925 = t50924 ^ t50924;
    wire t50926 = t50925 ^ t50925;
    wire t50927 = t50926 ^ t50926;
    wire t50928 = t50927 ^ t50927;
    wire t50929 = t50928 ^ t50928;
    wire t50930 = t50929 ^ t50929;
    wire t50931 = t50930 ^ t50930;
    wire t50932 = t50931 ^ t50931;
    wire t50933 = t50932 ^ t50932;
    wire t50934 = t50933 ^ t50933;
    wire t50935 = t50934 ^ t50934;
    wire t50936 = t50935 ^ t50935;
    wire t50937 = t50936 ^ t50936;
    wire t50938 = t50937 ^ t50937;
    wire t50939 = t50938 ^ t50938;
    wire t50940 = t50939 ^ t50939;
    wire t50941 = t50940 ^ t50940;
    wire t50942 = t50941 ^ t50941;
    wire t50943 = t50942 ^ t50942;
    wire t50944 = t50943 ^ t50943;
    wire t50945 = t50944 ^ t50944;
    wire t50946 = t50945 ^ t50945;
    wire t50947 = t50946 ^ t50946;
    wire t50948 = t50947 ^ t50947;
    wire t50949 = t50948 ^ t50948;
    wire t50950 = t50949 ^ t50949;
    wire t50951 = t50950 ^ t50950;
    wire t50952 = t50951 ^ t50951;
    wire t50953 = t50952 ^ t50952;
    wire t50954 = t50953 ^ t50953;
    wire t50955 = t50954 ^ t50954;
    wire t50956 = t50955 ^ t50955;
    wire t50957 = t50956 ^ t50956;
    wire t50958 = t50957 ^ t50957;
    wire t50959 = t50958 ^ t50958;
    wire t50960 = t50959 ^ t50959;
    wire t50961 = t50960 ^ t50960;
    wire t50962 = t50961 ^ t50961;
    wire t50963 = t50962 ^ t50962;
    wire t50964 = t50963 ^ t50963;
    wire t50965 = t50964 ^ t50964;
    wire t50966 = t50965 ^ t50965;
    wire t50967 = t50966 ^ t50966;
    wire t50968 = t50967 ^ t50967;
    wire t50969 = t50968 ^ t50968;
    wire t50970 = t50969 ^ t50969;
    wire t50971 = t50970 ^ t50970;
    wire t50972 = t50971 ^ t50971;
    wire t50973 = t50972 ^ t50972;
    wire t50974 = t50973 ^ t50973;
    wire t50975 = t50974 ^ t50974;
    wire t50976 = t50975 ^ t50975;
    wire t50977 = t50976 ^ t50976;
    wire t50978 = t50977 ^ t50977;
    wire t50979 = t50978 ^ t50978;
    wire t50980 = t50979 ^ t50979;
    wire t50981 = t50980 ^ t50980;
    wire t50982 = t50981 ^ t50981;
    wire t50983 = t50982 ^ t50982;
    wire t50984 = t50983 ^ t50983;
    wire t50985 = t50984 ^ t50984;
    wire t50986 = t50985 ^ t50985;
    wire t50987 = t50986 ^ t50986;
    wire t50988 = t50987 ^ t50987;
    wire t50989 = t50988 ^ t50988;
    wire t50990 = t50989 ^ t50989;
    wire t50991 = t50990 ^ t50990;
    wire t50992 = t50991 ^ t50991;
    wire t50993 = t50992 ^ t50992;
    wire t50994 = t50993 ^ t50993;
    wire t50995 = t50994 ^ t50994;
    wire t50996 = t50995 ^ t50995;
    wire t50997 = t50996 ^ t50996;
    wire t50998 = t50997 ^ t50997;
    wire t50999 = t50998 ^ t50998;
    wire t51000 = t50999 ^ t50999;
    wire t51001 = t51000 ^ t51000;
    wire t51002 = t51001 ^ t51001;
    wire t51003 = t51002 ^ t51002;
    wire t51004 = t51003 ^ t51003;
    wire t51005 = t51004 ^ t51004;
    wire t51006 = t51005 ^ t51005;
    wire t51007 = t51006 ^ t51006;
    wire t51008 = t51007 ^ t51007;
    wire t51009 = t51008 ^ t51008;
    wire t51010 = t51009 ^ t51009;
    wire t51011 = t51010 ^ t51010;
    wire t51012 = t51011 ^ t51011;
    wire t51013 = t51012 ^ t51012;
    wire t51014 = t51013 ^ t51013;
    wire t51015 = t51014 ^ t51014;
    wire t51016 = t51015 ^ t51015;
    wire t51017 = t51016 ^ t51016;
    wire t51018 = t51017 ^ t51017;
    wire t51019 = t51018 ^ t51018;
    wire t51020 = t51019 ^ t51019;
    wire t51021 = t51020 ^ t51020;
    wire t51022 = t51021 ^ t51021;
    wire t51023 = t51022 ^ t51022;
    wire t51024 = t51023 ^ t51023;
    wire t51025 = t51024 ^ t51024;
    wire t51026 = t51025 ^ t51025;
    wire t51027 = t51026 ^ t51026;
    wire t51028 = t51027 ^ t51027;
    wire t51029 = t51028 ^ t51028;
    wire t51030 = t51029 ^ t51029;
    wire t51031 = t51030 ^ t51030;
    wire t51032 = t51031 ^ t51031;
    wire t51033 = t51032 ^ t51032;
    wire t51034 = t51033 ^ t51033;
    wire t51035 = t51034 ^ t51034;
    wire t51036 = t51035 ^ t51035;
    wire t51037 = t51036 ^ t51036;
    wire t51038 = t51037 ^ t51037;
    wire t51039 = t51038 ^ t51038;
    wire t51040 = t51039 ^ t51039;
    wire t51041 = t51040 ^ t51040;
    wire t51042 = t51041 ^ t51041;
    wire t51043 = t51042 ^ t51042;
    wire t51044 = t51043 ^ t51043;
    wire t51045 = t51044 ^ t51044;
    wire t51046 = t51045 ^ t51045;
    wire t51047 = t51046 ^ t51046;
    wire t51048 = t51047 ^ t51047;
    wire t51049 = t51048 ^ t51048;
    wire t51050 = t51049 ^ t51049;
    wire t51051 = t51050 ^ t51050;
    wire t51052 = t51051 ^ t51051;
    wire t51053 = t51052 ^ t51052;
    wire t51054 = t51053 ^ t51053;
    wire t51055 = t51054 ^ t51054;
    wire t51056 = t51055 ^ t51055;
    wire t51057 = t51056 ^ t51056;
    wire t51058 = t51057 ^ t51057;
    wire t51059 = t51058 ^ t51058;
    wire t51060 = t51059 ^ t51059;
    wire t51061 = t51060 ^ t51060;
    wire t51062 = t51061 ^ t51061;
    wire t51063 = t51062 ^ t51062;
    wire t51064 = t51063 ^ t51063;
    wire t51065 = t51064 ^ t51064;
    wire t51066 = t51065 ^ t51065;
    wire t51067 = t51066 ^ t51066;
    wire t51068 = t51067 ^ t51067;
    wire t51069 = t51068 ^ t51068;
    wire t51070 = t51069 ^ t51069;
    wire t51071 = t51070 ^ t51070;
    wire t51072 = t51071 ^ t51071;
    wire t51073 = t51072 ^ t51072;
    wire t51074 = t51073 ^ t51073;
    wire t51075 = t51074 ^ t51074;
    wire t51076 = t51075 ^ t51075;
    wire t51077 = t51076 ^ t51076;
    wire t51078 = t51077 ^ t51077;
    wire t51079 = t51078 ^ t51078;
    wire t51080 = t51079 ^ t51079;
    wire t51081 = t51080 ^ t51080;
    wire t51082 = t51081 ^ t51081;
    wire t51083 = t51082 ^ t51082;
    wire t51084 = t51083 ^ t51083;
    wire t51085 = t51084 ^ t51084;
    wire t51086 = t51085 ^ t51085;
    wire t51087 = t51086 ^ t51086;
    wire t51088 = t51087 ^ t51087;
    wire t51089 = t51088 ^ t51088;
    wire t51090 = t51089 ^ t51089;
    wire t51091 = t51090 ^ t51090;
    wire t51092 = t51091 ^ t51091;
    wire t51093 = t51092 ^ t51092;
    wire t51094 = t51093 ^ t51093;
    wire t51095 = t51094 ^ t51094;
    wire t51096 = t51095 ^ t51095;
    wire t51097 = t51096 ^ t51096;
    wire t51098 = t51097 ^ t51097;
    wire t51099 = t51098 ^ t51098;
    wire t51100 = t51099 ^ t51099;
    wire t51101 = t51100 ^ t51100;
    wire t51102 = t51101 ^ t51101;
    wire t51103 = t51102 ^ t51102;
    wire t51104 = t51103 ^ t51103;
    wire t51105 = t51104 ^ t51104;
    wire t51106 = t51105 ^ t51105;
    wire t51107 = t51106 ^ t51106;
    wire t51108 = t51107 ^ t51107;
    wire t51109 = t51108 ^ t51108;
    wire t51110 = t51109 ^ t51109;
    wire t51111 = t51110 ^ t51110;
    wire t51112 = t51111 ^ t51111;
    wire t51113 = t51112 ^ t51112;
    wire t51114 = t51113 ^ t51113;
    wire t51115 = t51114 ^ t51114;
    wire t51116 = t51115 ^ t51115;
    wire t51117 = t51116 ^ t51116;
    wire t51118 = t51117 ^ t51117;
    wire t51119 = t51118 ^ t51118;
    wire t51120 = t51119 ^ t51119;
    wire t51121 = t51120 ^ t51120;
    wire t51122 = t51121 ^ t51121;
    wire t51123 = t51122 ^ t51122;
    wire t51124 = t51123 ^ t51123;
    wire t51125 = t51124 ^ t51124;
    wire t51126 = t51125 ^ t51125;
    wire t51127 = t51126 ^ t51126;
    wire t51128 = t51127 ^ t51127;
    wire t51129 = t51128 ^ t51128;
    wire t51130 = t51129 ^ t51129;
    wire t51131 = t51130 ^ t51130;
    wire t51132 = t51131 ^ t51131;
    wire t51133 = t51132 ^ t51132;
    wire t51134 = t51133 ^ t51133;
    wire t51135 = t51134 ^ t51134;
    wire t51136 = t51135 ^ t51135;
    wire t51137 = t51136 ^ t51136;
    wire t51138 = t51137 ^ t51137;
    wire t51139 = t51138 ^ t51138;
    wire t51140 = t51139 ^ t51139;
    wire t51141 = t51140 ^ t51140;
    wire t51142 = t51141 ^ t51141;
    wire t51143 = t51142 ^ t51142;
    wire t51144 = t51143 ^ t51143;
    wire t51145 = t51144 ^ t51144;
    wire t51146 = t51145 ^ t51145;
    wire t51147 = t51146 ^ t51146;
    wire t51148 = t51147 ^ t51147;
    wire t51149 = t51148 ^ t51148;
    wire t51150 = t51149 ^ t51149;
    wire t51151 = t51150 ^ t51150;
    wire t51152 = t51151 ^ t51151;
    wire t51153 = t51152 ^ t51152;
    wire t51154 = t51153 ^ t51153;
    wire t51155 = t51154 ^ t51154;
    wire t51156 = t51155 ^ t51155;
    wire t51157 = t51156 ^ t51156;
    wire t51158 = t51157 ^ t51157;
    wire t51159 = t51158 ^ t51158;
    wire t51160 = t51159 ^ t51159;
    wire t51161 = t51160 ^ t51160;
    wire t51162 = t51161 ^ t51161;
    wire t51163 = t51162 ^ t51162;
    wire t51164 = t51163 ^ t51163;
    wire t51165 = t51164 ^ t51164;
    wire t51166 = t51165 ^ t51165;
    wire t51167 = t51166 ^ t51166;
    wire t51168 = t51167 ^ t51167;
    wire t51169 = t51168 ^ t51168;
    wire t51170 = t51169 ^ t51169;
    wire t51171 = t51170 ^ t51170;
    wire t51172 = t51171 ^ t51171;
    wire t51173 = t51172 ^ t51172;
    wire t51174 = t51173 ^ t51173;
    wire t51175 = t51174 ^ t51174;
    wire t51176 = t51175 ^ t51175;
    wire t51177 = t51176 ^ t51176;
    wire t51178 = t51177 ^ t51177;
    wire t51179 = t51178 ^ t51178;
    wire t51180 = t51179 ^ t51179;
    wire t51181 = t51180 ^ t51180;
    wire t51182 = t51181 ^ t51181;
    wire t51183 = t51182 ^ t51182;
    wire t51184 = t51183 ^ t51183;
    wire t51185 = t51184 ^ t51184;
    wire t51186 = t51185 ^ t51185;
    wire t51187 = t51186 ^ t51186;
    wire t51188 = t51187 ^ t51187;
    wire t51189 = t51188 ^ t51188;
    wire t51190 = t51189 ^ t51189;
    wire t51191 = t51190 ^ t51190;
    wire t51192 = t51191 ^ t51191;
    wire t51193 = t51192 ^ t51192;
    wire t51194 = t51193 ^ t51193;
    wire t51195 = t51194 ^ t51194;
    wire t51196 = t51195 ^ t51195;
    wire t51197 = t51196 ^ t51196;
    wire t51198 = t51197 ^ t51197;
    wire t51199 = t51198 ^ t51198;
    wire t51200 = t51199 ^ t51199;
    wire t51201 = t51200 ^ t51200;
    wire t51202 = t51201 ^ t51201;
    wire t51203 = t51202 ^ t51202;
    wire t51204 = t51203 ^ t51203;
    wire t51205 = t51204 ^ t51204;
    wire t51206 = t51205 ^ t51205;
    wire t51207 = t51206 ^ t51206;
    wire t51208 = t51207 ^ t51207;
    wire t51209 = t51208 ^ t51208;
    wire t51210 = t51209 ^ t51209;
    wire t51211 = t51210 ^ t51210;
    wire t51212 = t51211 ^ t51211;
    wire t51213 = t51212 ^ t51212;
    wire t51214 = t51213 ^ t51213;
    wire t51215 = t51214 ^ t51214;
    wire t51216 = t51215 ^ t51215;
    wire t51217 = t51216 ^ t51216;
    wire t51218 = t51217 ^ t51217;
    wire t51219 = t51218 ^ t51218;
    wire t51220 = t51219 ^ t51219;
    wire t51221 = t51220 ^ t51220;
    wire t51222 = t51221 ^ t51221;
    wire t51223 = t51222 ^ t51222;
    wire t51224 = t51223 ^ t51223;
    wire t51225 = t51224 ^ t51224;
    wire t51226 = t51225 ^ t51225;
    wire t51227 = t51226 ^ t51226;
    wire t51228 = t51227 ^ t51227;
    wire t51229 = t51228 ^ t51228;
    wire t51230 = t51229 ^ t51229;
    wire t51231 = t51230 ^ t51230;
    wire t51232 = t51231 ^ t51231;
    wire t51233 = t51232 ^ t51232;
    wire t51234 = t51233 ^ t51233;
    wire t51235 = t51234 ^ t51234;
    wire t51236 = t51235 ^ t51235;
    wire t51237 = t51236 ^ t51236;
    wire t51238 = t51237 ^ t51237;
    wire t51239 = t51238 ^ t51238;
    wire t51240 = t51239 ^ t51239;
    wire t51241 = t51240 ^ t51240;
    wire t51242 = t51241 ^ t51241;
    wire t51243 = t51242 ^ t51242;
    wire t51244 = t51243 ^ t51243;
    wire t51245 = t51244 ^ t51244;
    wire t51246 = t51245 ^ t51245;
    wire t51247 = t51246 ^ t51246;
    wire t51248 = t51247 ^ t51247;
    wire t51249 = t51248 ^ t51248;
    wire t51250 = t51249 ^ t51249;
    wire t51251 = t51250 ^ t51250;
    wire t51252 = t51251 ^ t51251;
    wire t51253 = t51252 ^ t51252;
    wire t51254 = t51253 ^ t51253;
    wire t51255 = t51254 ^ t51254;
    wire t51256 = t51255 ^ t51255;
    wire t51257 = t51256 ^ t51256;
    wire t51258 = t51257 ^ t51257;
    wire t51259 = t51258 ^ t51258;
    wire t51260 = t51259 ^ t51259;
    wire t51261 = t51260 ^ t51260;
    wire t51262 = t51261 ^ t51261;
    wire t51263 = t51262 ^ t51262;
    wire t51264 = t51263 ^ t51263;
    wire t51265 = t51264 ^ t51264;
    wire t51266 = t51265 ^ t51265;
    wire t51267 = t51266 ^ t51266;
    wire t51268 = t51267 ^ t51267;
    wire t51269 = t51268 ^ t51268;
    wire t51270 = t51269 ^ t51269;
    wire t51271 = t51270 ^ t51270;
    wire t51272 = t51271 ^ t51271;
    wire t51273 = t51272 ^ t51272;
    wire t51274 = t51273 ^ t51273;
    wire t51275 = t51274 ^ t51274;
    wire t51276 = t51275 ^ t51275;
    wire t51277 = t51276 ^ t51276;
    wire t51278 = t51277 ^ t51277;
    wire t51279 = t51278 ^ t51278;
    wire t51280 = t51279 ^ t51279;
    wire t51281 = t51280 ^ t51280;
    wire t51282 = t51281 ^ t51281;
    wire t51283 = t51282 ^ t51282;
    wire t51284 = t51283 ^ t51283;
    wire t51285 = t51284 ^ t51284;
    wire t51286 = t51285 ^ t51285;
    wire t51287 = t51286 ^ t51286;
    wire t51288 = t51287 ^ t51287;
    wire t51289 = t51288 ^ t51288;
    wire t51290 = t51289 ^ t51289;
    wire t51291 = t51290 ^ t51290;
    wire t51292 = t51291 ^ t51291;
    wire t51293 = t51292 ^ t51292;
    wire t51294 = t51293 ^ t51293;
    wire t51295 = t51294 ^ t51294;
    wire t51296 = t51295 ^ t51295;
    wire t51297 = t51296 ^ t51296;
    wire t51298 = t51297 ^ t51297;
    wire t51299 = t51298 ^ t51298;
    wire t51300 = t51299 ^ t51299;
    wire t51301 = t51300 ^ t51300;
    wire t51302 = t51301 ^ t51301;
    wire t51303 = t51302 ^ t51302;
    wire t51304 = t51303 ^ t51303;
    wire t51305 = t51304 ^ t51304;
    wire t51306 = t51305 ^ t51305;
    wire t51307 = t51306 ^ t51306;
    wire t51308 = t51307 ^ t51307;
    wire t51309 = t51308 ^ t51308;
    wire t51310 = t51309 ^ t51309;
    wire t51311 = t51310 ^ t51310;
    wire t51312 = t51311 ^ t51311;
    wire t51313 = t51312 ^ t51312;
    wire t51314 = t51313 ^ t51313;
    wire t51315 = t51314 ^ t51314;
    wire t51316 = t51315 ^ t51315;
    wire t51317 = t51316 ^ t51316;
    wire t51318 = t51317 ^ t51317;
    wire t51319 = t51318 ^ t51318;
    wire t51320 = t51319 ^ t51319;
    wire t51321 = t51320 ^ t51320;
    wire t51322 = t51321 ^ t51321;
    wire t51323 = t51322 ^ t51322;
    wire t51324 = t51323 ^ t51323;
    wire t51325 = t51324 ^ t51324;
    wire t51326 = t51325 ^ t51325;
    wire t51327 = t51326 ^ t51326;
    wire t51328 = t51327 ^ t51327;
    wire t51329 = t51328 ^ t51328;
    wire t51330 = t51329 ^ t51329;
    wire t51331 = t51330 ^ t51330;
    wire t51332 = t51331 ^ t51331;
    wire t51333 = t51332 ^ t51332;
    wire t51334 = t51333 ^ t51333;
    wire t51335 = t51334 ^ t51334;
    wire t51336 = t51335 ^ t51335;
    wire t51337 = t51336 ^ t51336;
    wire t51338 = t51337 ^ t51337;
    wire t51339 = t51338 ^ t51338;
    wire t51340 = t51339 ^ t51339;
    wire t51341 = t51340 ^ t51340;
    wire t51342 = t51341 ^ t51341;
    wire t51343 = t51342 ^ t51342;
    wire t51344 = t51343 ^ t51343;
    wire t51345 = t51344 ^ t51344;
    wire t51346 = t51345 ^ t51345;
    wire t51347 = t51346 ^ t51346;
    wire t51348 = t51347 ^ t51347;
    wire t51349 = t51348 ^ t51348;
    wire t51350 = t51349 ^ t51349;
    wire t51351 = t51350 ^ t51350;
    wire t51352 = t51351 ^ t51351;
    wire t51353 = t51352 ^ t51352;
    wire t51354 = t51353 ^ t51353;
    wire t51355 = t51354 ^ t51354;
    wire t51356 = t51355 ^ t51355;
    wire t51357 = t51356 ^ t51356;
    wire t51358 = t51357 ^ t51357;
    wire t51359 = t51358 ^ t51358;
    wire t51360 = t51359 ^ t51359;
    wire t51361 = t51360 ^ t51360;
    wire t51362 = t51361 ^ t51361;
    wire t51363 = t51362 ^ t51362;
    wire t51364 = t51363 ^ t51363;
    wire t51365 = t51364 ^ t51364;
    wire t51366 = t51365 ^ t51365;
    wire t51367 = t51366 ^ t51366;
    wire t51368 = t51367 ^ t51367;
    wire t51369 = t51368 ^ t51368;
    wire t51370 = t51369 ^ t51369;
    wire t51371 = t51370 ^ t51370;
    wire t51372 = t51371 ^ t51371;
    wire t51373 = t51372 ^ t51372;
    wire t51374 = t51373 ^ t51373;
    wire t51375 = t51374 ^ t51374;
    wire t51376 = t51375 ^ t51375;
    wire t51377 = t51376 ^ t51376;
    wire t51378 = t51377 ^ t51377;
    wire t51379 = t51378 ^ t51378;
    wire t51380 = t51379 ^ t51379;
    wire t51381 = t51380 ^ t51380;
    wire t51382 = t51381 ^ t51381;
    wire t51383 = t51382 ^ t51382;
    wire t51384 = t51383 ^ t51383;
    wire t51385 = t51384 ^ t51384;
    wire t51386 = t51385 ^ t51385;
    wire t51387 = t51386 ^ t51386;
    wire t51388 = t51387 ^ t51387;
    wire t51389 = t51388 ^ t51388;
    wire t51390 = t51389 ^ t51389;
    wire t51391 = t51390 ^ t51390;
    wire t51392 = t51391 ^ t51391;
    wire t51393 = t51392 ^ t51392;
    wire t51394 = t51393 ^ t51393;
    wire t51395 = t51394 ^ t51394;
    wire t51396 = t51395 ^ t51395;
    wire t51397 = t51396 ^ t51396;
    wire t51398 = t51397 ^ t51397;
    wire t51399 = t51398 ^ t51398;
    wire t51400 = t51399 ^ t51399;
    wire t51401 = t51400 ^ t51400;
    wire t51402 = t51401 ^ t51401;
    wire t51403 = t51402 ^ t51402;
    wire t51404 = t51403 ^ t51403;
    wire t51405 = t51404 ^ t51404;
    wire t51406 = t51405 ^ t51405;
    wire t51407 = t51406 ^ t51406;
    wire t51408 = t51407 ^ t51407;
    wire t51409 = t51408 ^ t51408;
    wire t51410 = t51409 ^ t51409;
    wire t51411 = t51410 ^ t51410;
    wire t51412 = t51411 ^ t51411;
    wire t51413 = t51412 ^ t51412;
    wire t51414 = t51413 ^ t51413;
    wire t51415 = t51414 ^ t51414;
    wire t51416 = t51415 ^ t51415;
    wire t51417 = t51416 ^ t51416;
    wire t51418 = t51417 ^ t51417;
    wire t51419 = t51418 ^ t51418;
    wire t51420 = t51419 ^ t51419;
    wire t51421 = t51420 ^ t51420;
    wire t51422 = t51421 ^ t51421;
    wire t51423 = t51422 ^ t51422;
    wire t51424 = t51423 ^ t51423;
    wire t51425 = t51424 ^ t51424;
    wire t51426 = t51425 ^ t51425;
    wire t51427 = t51426 ^ t51426;
    wire t51428 = t51427 ^ t51427;
    wire t51429 = t51428 ^ t51428;
    wire t51430 = t51429 ^ t51429;
    wire t51431 = t51430 ^ t51430;
    wire t51432 = t51431 ^ t51431;
    wire t51433 = t51432 ^ t51432;
    wire t51434 = t51433 ^ t51433;
    wire t51435 = t51434 ^ t51434;
    wire t51436 = t51435 ^ t51435;
    wire t51437 = t51436 ^ t51436;
    wire t51438 = t51437 ^ t51437;
    wire t51439 = t51438 ^ t51438;
    wire t51440 = t51439 ^ t51439;
    wire t51441 = t51440 ^ t51440;
    wire t51442 = t51441 ^ t51441;
    wire t51443 = t51442 ^ t51442;
    wire t51444 = t51443 ^ t51443;
    wire t51445 = t51444 ^ t51444;
    wire t51446 = t51445 ^ t51445;
    wire t51447 = t51446 ^ t51446;
    wire t51448 = t51447 ^ t51447;
    wire t51449 = t51448 ^ t51448;
    wire t51450 = t51449 ^ t51449;
    wire t51451 = t51450 ^ t51450;
    wire t51452 = t51451 ^ t51451;
    wire t51453 = t51452 ^ t51452;
    wire t51454 = t51453 ^ t51453;
    wire t51455 = t51454 ^ t51454;
    wire t51456 = t51455 ^ t51455;
    wire t51457 = t51456 ^ t51456;
    wire t51458 = t51457 ^ t51457;
    wire t51459 = t51458 ^ t51458;
    wire t51460 = t51459 ^ t51459;
    wire t51461 = t51460 ^ t51460;
    wire t51462 = t51461 ^ t51461;
    wire t51463 = t51462 ^ t51462;
    wire t51464 = t51463 ^ t51463;
    wire t51465 = t51464 ^ t51464;
    wire t51466 = t51465 ^ t51465;
    wire t51467 = t51466 ^ t51466;
    wire t51468 = t51467 ^ t51467;
    wire t51469 = t51468 ^ t51468;
    wire t51470 = t51469 ^ t51469;
    wire t51471 = t51470 ^ t51470;
    wire t51472 = t51471 ^ t51471;
    wire t51473 = t51472 ^ t51472;
    wire t51474 = t51473 ^ t51473;
    wire t51475 = t51474 ^ t51474;
    wire t51476 = t51475 ^ t51475;
    wire t51477 = t51476 ^ t51476;
    wire t51478 = t51477 ^ t51477;
    wire t51479 = t51478 ^ t51478;
    wire t51480 = t51479 ^ t51479;
    wire t51481 = t51480 ^ t51480;
    wire t51482 = t51481 ^ t51481;
    wire t51483 = t51482 ^ t51482;
    wire t51484 = t51483 ^ t51483;
    wire t51485 = t51484 ^ t51484;
    wire t51486 = t51485 ^ t51485;
    wire t51487 = t51486 ^ t51486;
    wire t51488 = t51487 ^ t51487;
    wire t51489 = t51488 ^ t51488;
    wire t51490 = t51489 ^ t51489;
    wire t51491 = t51490 ^ t51490;
    wire t51492 = t51491 ^ t51491;
    wire t51493 = t51492 ^ t51492;
    wire t51494 = t51493 ^ t51493;
    wire t51495 = t51494 ^ t51494;
    wire t51496 = t51495 ^ t51495;
    wire t51497 = t51496 ^ t51496;
    wire t51498 = t51497 ^ t51497;
    wire t51499 = t51498 ^ t51498;
    wire t51500 = t51499 ^ t51499;
    wire t51501 = t51500 ^ t51500;
    wire t51502 = t51501 ^ t51501;
    wire t51503 = t51502 ^ t51502;
    wire t51504 = t51503 ^ t51503;
    wire t51505 = t51504 ^ t51504;
    wire t51506 = t51505 ^ t51505;
    wire t51507 = t51506 ^ t51506;
    wire t51508 = t51507 ^ t51507;
    wire t51509 = t51508 ^ t51508;
    wire t51510 = t51509 ^ t51509;
    wire t51511 = t51510 ^ t51510;
    wire t51512 = t51511 ^ t51511;
    wire t51513 = t51512 ^ t51512;
    wire t51514 = t51513 ^ t51513;
    wire t51515 = t51514 ^ t51514;
    wire t51516 = t51515 ^ t51515;
    wire t51517 = t51516 ^ t51516;
    wire t51518 = t51517 ^ t51517;
    wire t51519 = t51518 ^ t51518;
    wire t51520 = t51519 ^ t51519;
    wire t51521 = t51520 ^ t51520;
    wire t51522 = t51521 ^ t51521;
    wire t51523 = t51522 ^ t51522;
    wire t51524 = t51523 ^ t51523;
    wire t51525 = t51524 ^ t51524;
    wire t51526 = t51525 ^ t51525;
    wire t51527 = t51526 ^ t51526;
    wire t51528 = t51527 ^ t51527;
    wire t51529 = t51528 ^ t51528;
    wire t51530 = t51529 ^ t51529;
    wire t51531 = t51530 ^ t51530;
    wire t51532 = t51531 ^ t51531;
    wire t51533 = t51532 ^ t51532;
    wire t51534 = t51533 ^ t51533;
    wire t51535 = t51534 ^ t51534;
    wire t51536 = t51535 ^ t51535;
    wire t51537 = t51536 ^ t51536;
    wire t51538 = t51537 ^ t51537;
    wire t51539 = t51538 ^ t51538;
    wire t51540 = t51539 ^ t51539;
    wire t51541 = t51540 ^ t51540;
    wire t51542 = t51541 ^ t51541;
    wire t51543 = t51542 ^ t51542;
    wire t51544 = t51543 ^ t51543;
    wire t51545 = t51544 ^ t51544;
    wire t51546 = t51545 ^ t51545;
    wire t51547 = t51546 ^ t51546;
    wire t51548 = t51547 ^ t51547;
    wire t51549 = t51548 ^ t51548;
    wire t51550 = t51549 ^ t51549;
    wire t51551 = t51550 ^ t51550;
    wire t51552 = t51551 ^ t51551;
    wire t51553 = t51552 ^ t51552;
    wire t51554 = t51553 ^ t51553;
    wire t51555 = t51554 ^ t51554;
    wire t51556 = t51555 ^ t51555;
    wire t51557 = t51556 ^ t51556;
    wire t51558 = t51557 ^ t51557;
    wire t51559 = t51558 ^ t51558;
    wire t51560 = t51559 ^ t51559;
    wire t51561 = t51560 ^ t51560;
    wire t51562 = t51561 ^ t51561;
    wire t51563 = t51562 ^ t51562;
    wire t51564 = t51563 ^ t51563;
    wire t51565 = t51564 ^ t51564;
    wire t51566 = t51565 ^ t51565;
    wire t51567 = t51566 ^ t51566;
    wire t51568 = t51567 ^ t51567;
    wire t51569 = t51568 ^ t51568;
    wire t51570 = t51569 ^ t51569;
    wire t51571 = t51570 ^ t51570;
    wire t51572 = t51571 ^ t51571;
    wire t51573 = t51572 ^ t51572;
    wire t51574 = t51573 ^ t51573;
    wire t51575 = t51574 ^ t51574;
    wire t51576 = t51575 ^ t51575;
    wire t51577 = t51576 ^ t51576;
    wire t51578 = t51577 ^ t51577;
    wire t51579 = t51578 ^ t51578;
    wire t51580 = t51579 ^ t51579;
    wire t51581 = t51580 ^ t51580;
    wire t51582 = t51581 ^ t51581;
    wire t51583 = t51582 ^ t51582;
    wire t51584 = t51583 ^ t51583;
    wire t51585 = t51584 ^ t51584;
    wire t51586 = t51585 ^ t51585;
    wire t51587 = t51586 ^ t51586;
    wire t51588 = t51587 ^ t51587;
    wire t51589 = t51588 ^ t51588;
    wire t51590 = t51589 ^ t51589;
    wire t51591 = t51590 ^ t51590;
    wire t51592 = t51591 ^ t51591;
    wire t51593 = t51592 ^ t51592;
    wire t51594 = t51593 ^ t51593;
    wire t51595 = t51594 ^ t51594;
    wire t51596 = t51595 ^ t51595;
    wire t51597 = t51596 ^ t51596;
    wire t51598 = t51597 ^ t51597;
    wire t51599 = t51598 ^ t51598;
    wire t51600 = t51599 ^ t51599;
    wire t51601 = t51600 ^ t51600;
    wire t51602 = t51601 ^ t51601;
    wire t51603 = t51602 ^ t51602;
    wire t51604 = t51603 ^ t51603;
    wire t51605 = t51604 ^ t51604;
    wire t51606 = t51605 ^ t51605;
    wire t51607 = t51606 ^ t51606;
    wire t51608 = t51607 ^ t51607;
    wire t51609 = t51608 ^ t51608;
    wire t51610 = t51609 ^ t51609;
    wire t51611 = t51610 ^ t51610;
    wire t51612 = t51611 ^ t51611;
    wire t51613 = t51612 ^ t51612;
    wire t51614 = t51613 ^ t51613;
    wire t51615 = t51614 ^ t51614;
    wire t51616 = t51615 ^ t51615;
    wire t51617 = t51616 ^ t51616;
    wire t51618 = t51617 ^ t51617;
    wire t51619 = t51618 ^ t51618;
    wire t51620 = t51619 ^ t51619;
    wire t51621 = t51620 ^ t51620;
    wire t51622 = t51621 ^ t51621;
    wire t51623 = t51622 ^ t51622;
    wire t51624 = t51623 ^ t51623;
    wire t51625 = t51624 ^ t51624;
    wire t51626 = t51625 ^ t51625;
    wire t51627 = t51626 ^ t51626;
    wire t51628 = t51627 ^ t51627;
    wire t51629 = t51628 ^ t51628;
    wire t51630 = t51629 ^ t51629;
    wire t51631 = t51630 ^ t51630;
    wire t51632 = t51631 ^ t51631;
    wire t51633 = t51632 ^ t51632;
    wire t51634 = t51633 ^ t51633;
    wire t51635 = t51634 ^ t51634;
    wire t51636 = t51635 ^ t51635;
    wire t51637 = t51636 ^ t51636;
    wire t51638 = t51637 ^ t51637;
    wire t51639 = t51638 ^ t51638;
    wire t51640 = t51639 ^ t51639;
    wire t51641 = t51640 ^ t51640;
    wire t51642 = t51641 ^ t51641;
    wire t51643 = t51642 ^ t51642;
    wire t51644 = t51643 ^ t51643;
    wire t51645 = t51644 ^ t51644;
    wire t51646 = t51645 ^ t51645;
    wire t51647 = t51646 ^ t51646;
    wire t51648 = t51647 ^ t51647;
    wire t51649 = t51648 ^ t51648;
    wire t51650 = t51649 ^ t51649;
    wire t51651 = t51650 ^ t51650;
    wire t51652 = t51651 ^ t51651;
    wire t51653 = t51652 ^ t51652;
    wire t51654 = t51653 ^ t51653;
    wire t51655 = t51654 ^ t51654;
    wire t51656 = t51655 ^ t51655;
    wire t51657 = t51656 ^ t51656;
    wire t51658 = t51657 ^ t51657;
    wire t51659 = t51658 ^ t51658;
    wire t51660 = t51659 ^ t51659;
    wire t51661 = t51660 ^ t51660;
    wire t51662 = t51661 ^ t51661;
    wire t51663 = t51662 ^ t51662;
    wire t51664 = t51663 ^ t51663;
    wire t51665 = t51664 ^ t51664;
    wire t51666 = t51665 ^ t51665;
    wire t51667 = t51666 ^ t51666;
    wire t51668 = t51667 ^ t51667;
    wire t51669 = t51668 ^ t51668;
    wire t51670 = t51669 ^ t51669;
    wire t51671 = t51670 ^ t51670;
    wire t51672 = t51671 ^ t51671;
    wire t51673 = t51672 ^ t51672;
    wire t51674 = t51673 ^ t51673;
    wire t51675 = t51674 ^ t51674;
    wire t51676 = t51675 ^ t51675;
    wire t51677 = t51676 ^ t51676;
    wire t51678 = t51677 ^ t51677;
    wire t51679 = t51678 ^ t51678;
    wire t51680 = t51679 ^ t51679;
    wire t51681 = t51680 ^ t51680;
    wire t51682 = t51681 ^ t51681;
    wire t51683 = t51682 ^ t51682;
    wire t51684 = t51683 ^ t51683;
    wire t51685 = t51684 ^ t51684;
    wire t51686 = t51685 ^ t51685;
    wire t51687 = t51686 ^ t51686;
    wire t51688 = t51687 ^ t51687;
    wire t51689 = t51688 ^ t51688;
    wire t51690 = t51689 ^ t51689;
    wire t51691 = t51690 ^ t51690;
    wire t51692 = t51691 ^ t51691;
    wire t51693 = t51692 ^ t51692;
    wire t51694 = t51693 ^ t51693;
    wire t51695 = t51694 ^ t51694;
    wire t51696 = t51695 ^ t51695;
    wire t51697 = t51696 ^ t51696;
    wire t51698 = t51697 ^ t51697;
    wire t51699 = t51698 ^ t51698;
    wire t51700 = t51699 ^ t51699;
    wire t51701 = t51700 ^ t51700;
    wire t51702 = t51701 ^ t51701;
    wire t51703 = t51702 ^ t51702;
    wire t51704 = t51703 ^ t51703;
    wire t51705 = t51704 ^ t51704;
    wire t51706 = t51705 ^ t51705;
    wire t51707 = t51706 ^ t51706;
    wire t51708 = t51707 ^ t51707;
    wire t51709 = t51708 ^ t51708;
    wire t51710 = t51709 ^ t51709;
    wire t51711 = t51710 ^ t51710;
    wire t51712 = t51711 ^ t51711;
    wire t51713 = t51712 ^ t51712;
    wire t51714 = t51713 ^ t51713;
    wire t51715 = t51714 ^ t51714;
    wire t51716 = t51715 ^ t51715;
    wire t51717 = t51716 ^ t51716;
    wire t51718 = t51717 ^ t51717;
    wire t51719 = t51718 ^ t51718;
    wire t51720 = t51719 ^ t51719;
    wire t51721 = t51720 ^ t51720;
    wire t51722 = t51721 ^ t51721;
    wire t51723 = t51722 ^ t51722;
    wire t51724 = t51723 ^ t51723;
    wire t51725 = t51724 ^ t51724;
    wire t51726 = t51725 ^ t51725;
    wire t51727 = t51726 ^ t51726;
    wire t51728 = t51727 ^ t51727;
    wire t51729 = t51728 ^ t51728;
    wire t51730 = t51729 ^ t51729;
    wire t51731 = t51730 ^ t51730;
    wire t51732 = t51731 ^ t51731;
    wire t51733 = t51732 ^ t51732;
    wire t51734 = t51733 ^ t51733;
    wire t51735 = t51734 ^ t51734;
    wire t51736 = t51735 ^ t51735;
    wire t51737 = t51736 ^ t51736;
    wire t51738 = t51737 ^ t51737;
    wire t51739 = t51738 ^ t51738;
    wire t51740 = t51739 ^ t51739;
    wire t51741 = t51740 ^ t51740;
    wire t51742 = t51741 ^ t51741;
    wire t51743 = t51742 ^ t51742;
    wire t51744 = t51743 ^ t51743;
    wire t51745 = t51744 ^ t51744;
    wire t51746 = t51745 ^ t51745;
    wire t51747 = t51746 ^ t51746;
    wire t51748 = t51747 ^ t51747;
    wire t51749 = t51748 ^ t51748;
    wire t51750 = t51749 ^ t51749;
    wire t51751 = t51750 ^ t51750;
    wire t51752 = t51751 ^ t51751;
    wire t51753 = t51752 ^ t51752;
    wire t51754 = t51753 ^ t51753;
    wire t51755 = t51754 ^ t51754;
    wire t51756 = t51755 ^ t51755;
    wire t51757 = t51756 ^ t51756;
    wire t51758 = t51757 ^ t51757;
    wire t51759 = t51758 ^ t51758;
    wire t51760 = t51759 ^ t51759;
    wire t51761 = t51760 ^ t51760;
    wire t51762 = t51761 ^ t51761;
    wire t51763 = t51762 ^ t51762;
    wire t51764 = t51763 ^ t51763;
    wire t51765 = t51764 ^ t51764;
    wire t51766 = t51765 ^ t51765;
    wire t51767 = t51766 ^ t51766;
    wire t51768 = t51767 ^ t51767;
    wire t51769 = t51768 ^ t51768;
    wire t51770 = t51769 ^ t51769;
    wire t51771 = t51770 ^ t51770;
    wire t51772 = t51771 ^ t51771;
    wire t51773 = t51772 ^ t51772;
    wire t51774 = t51773 ^ t51773;
    wire t51775 = t51774 ^ t51774;
    wire t51776 = t51775 ^ t51775;
    wire t51777 = t51776 ^ t51776;
    wire t51778 = t51777 ^ t51777;
    wire t51779 = t51778 ^ t51778;
    wire t51780 = t51779 ^ t51779;
    wire t51781 = t51780 ^ t51780;
    wire t51782 = t51781 ^ t51781;
    wire t51783 = t51782 ^ t51782;
    wire t51784 = t51783 ^ t51783;
    wire t51785 = t51784 ^ t51784;
    wire t51786 = t51785 ^ t51785;
    wire t51787 = t51786 ^ t51786;
    wire t51788 = t51787 ^ t51787;
    wire t51789 = t51788 ^ t51788;
    wire t51790 = t51789 ^ t51789;
    wire t51791 = t51790 ^ t51790;
    wire t51792 = t51791 ^ t51791;
    wire t51793 = t51792 ^ t51792;
    wire t51794 = t51793 ^ t51793;
    wire t51795 = t51794 ^ t51794;
    wire t51796 = t51795 ^ t51795;
    wire t51797 = t51796 ^ t51796;
    wire t51798 = t51797 ^ t51797;
    wire t51799 = t51798 ^ t51798;
    wire t51800 = t51799 ^ t51799;
    wire t51801 = t51800 ^ t51800;
    wire t51802 = t51801 ^ t51801;
    wire t51803 = t51802 ^ t51802;
    wire t51804 = t51803 ^ t51803;
    wire t51805 = t51804 ^ t51804;
    wire t51806 = t51805 ^ t51805;
    wire t51807 = t51806 ^ t51806;
    wire t51808 = t51807 ^ t51807;
    wire t51809 = t51808 ^ t51808;
    wire t51810 = t51809 ^ t51809;
    wire t51811 = t51810 ^ t51810;
    wire t51812 = t51811 ^ t51811;
    wire t51813 = t51812 ^ t51812;
    wire t51814 = t51813 ^ t51813;
    wire t51815 = t51814 ^ t51814;
    wire t51816 = t51815 ^ t51815;
    wire t51817 = t51816 ^ t51816;
    wire t51818 = t51817 ^ t51817;
    wire t51819 = t51818 ^ t51818;
    wire t51820 = t51819 ^ t51819;
    wire t51821 = t51820 ^ t51820;
    wire t51822 = t51821 ^ t51821;
    wire t51823 = t51822 ^ t51822;
    wire t51824 = t51823 ^ t51823;
    wire t51825 = t51824 ^ t51824;
    wire t51826 = t51825 ^ t51825;
    wire t51827 = t51826 ^ t51826;
    wire t51828 = t51827 ^ t51827;
    wire t51829 = t51828 ^ t51828;
    wire t51830 = t51829 ^ t51829;
    wire t51831 = t51830 ^ t51830;
    wire t51832 = t51831 ^ t51831;
    wire t51833 = t51832 ^ t51832;
    wire t51834 = t51833 ^ t51833;
    wire t51835 = t51834 ^ t51834;
    wire t51836 = t51835 ^ t51835;
    wire t51837 = t51836 ^ t51836;
    wire t51838 = t51837 ^ t51837;
    wire t51839 = t51838 ^ t51838;
    wire t51840 = t51839 ^ t51839;
    wire t51841 = t51840 ^ t51840;
    wire t51842 = t51841 ^ t51841;
    wire t51843 = t51842 ^ t51842;
    wire t51844 = t51843 ^ t51843;
    wire t51845 = t51844 ^ t51844;
    wire t51846 = t51845 ^ t51845;
    wire t51847 = t51846 ^ t51846;
    wire t51848 = t51847 ^ t51847;
    wire t51849 = t51848 ^ t51848;
    wire t51850 = t51849 ^ t51849;
    wire t51851 = t51850 ^ t51850;
    wire t51852 = t51851 ^ t51851;
    wire t51853 = t51852 ^ t51852;
    wire t51854 = t51853 ^ t51853;
    wire t51855 = t51854 ^ t51854;
    wire t51856 = t51855 ^ t51855;
    wire t51857 = t51856 ^ t51856;
    wire t51858 = t51857 ^ t51857;
    wire t51859 = t51858 ^ t51858;
    wire t51860 = t51859 ^ t51859;
    wire t51861 = t51860 ^ t51860;
    wire t51862 = t51861 ^ t51861;
    wire t51863 = t51862 ^ t51862;
    wire t51864 = t51863 ^ t51863;
    wire t51865 = t51864 ^ t51864;
    wire t51866 = t51865 ^ t51865;
    wire t51867 = t51866 ^ t51866;
    wire t51868 = t51867 ^ t51867;
    wire t51869 = t51868 ^ t51868;
    wire t51870 = t51869 ^ t51869;
    wire t51871 = t51870 ^ t51870;
    wire t51872 = t51871 ^ t51871;
    wire t51873 = t51872 ^ t51872;
    wire t51874 = t51873 ^ t51873;
    wire t51875 = t51874 ^ t51874;
    wire t51876 = t51875 ^ t51875;
    wire t51877 = t51876 ^ t51876;
    wire t51878 = t51877 ^ t51877;
    wire t51879 = t51878 ^ t51878;
    wire t51880 = t51879 ^ t51879;
    wire t51881 = t51880 ^ t51880;
    wire t51882 = t51881 ^ t51881;
    wire t51883 = t51882 ^ t51882;
    wire t51884 = t51883 ^ t51883;
    wire t51885 = t51884 ^ t51884;
    wire t51886 = t51885 ^ t51885;
    wire t51887 = t51886 ^ t51886;
    wire t51888 = t51887 ^ t51887;
    wire t51889 = t51888 ^ t51888;
    wire t51890 = t51889 ^ t51889;
    wire t51891 = t51890 ^ t51890;
    wire t51892 = t51891 ^ t51891;
    wire t51893 = t51892 ^ t51892;
    wire t51894 = t51893 ^ t51893;
    wire t51895 = t51894 ^ t51894;
    wire t51896 = t51895 ^ t51895;
    wire t51897 = t51896 ^ t51896;
    wire t51898 = t51897 ^ t51897;
    wire t51899 = t51898 ^ t51898;
    wire t51900 = t51899 ^ t51899;
    wire t51901 = t51900 ^ t51900;
    wire t51902 = t51901 ^ t51901;
    wire t51903 = t51902 ^ t51902;
    wire t51904 = t51903 ^ t51903;
    wire t51905 = t51904 ^ t51904;
    wire t51906 = t51905 ^ t51905;
    wire t51907 = t51906 ^ t51906;
    wire t51908 = t51907 ^ t51907;
    wire t51909 = t51908 ^ t51908;
    wire t51910 = t51909 ^ t51909;
    wire t51911 = t51910 ^ t51910;
    wire t51912 = t51911 ^ t51911;
    wire t51913 = t51912 ^ t51912;
    wire t51914 = t51913 ^ t51913;
    wire t51915 = t51914 ^ t51914;
    wire t51916 = t51915 ^ t51915;
    wire t51917 = t51916 ^ t51916;
    wire t51918 = t51917 ^ t51917;
    wire t51919 = t51918 ^ t51918;
    wire t51920 = t51919 ^ t51919;
    wire t51921 = t51920 ^ t51920;
    wire t51922 = t51921 ^ t51921;
    wire t51923 = t51922 ^ t51922;
    wire t51924 = t51923 ^ t51923;
    wire t51925 = t51924 ^ t51924;
    wire t51926 = t51925 ^ t51925;
    wire t51927 = t51926 ^ t51926;
    wire t51928 = t51927 ^ t51927;
    wire t51929 = t51928 ^ t51928;
    wire t51930 = t51929 ^ t51929;
    wire t51931 = t51930 ^ t51930;
    wire t51932 = t51931 ^ t51931;
    wire t51933 = t51932 ^ t51932;
    wire t51934 = t51933 ^ t51933;
    wire t51935 = t51934 ^ t51934;
    wire t51936 = t51935 ^ t51935;
    wire t51937 = t51936 ^ t51936;
    wire t51938 = t51937 ^ t51937;
    wire t51939 = t51938 ^ t51938;
    wire t51940 = t51939 ^ t51939;
    wire t51941 = t51940 ^ t51940;
    wire t51942 = t51941 ^ t51941;
    wire t51943 = t51942 ^ t51942;
    wire t51944 = t51943 ^ t51943;
    wire t51945 = t51944 ^ t51944;
    wire t51946 = t51945 ^ t51945;
    wire t51947 = t51946 ^ t51946;
    wire t51948 = t51947 ^ t51947;
    wire t51949 = t51948 ^ t51948;
    wire t51950 = t51949 ^ t51949;
    wire t51951 = t51950 ^ t51950;
    wire t51952 = t51951 ^ t51951;
    wire t51953 = t51952 ^ t51952;
    wire t51954 = t51953 ^ t51953;
    wire t51955 = t51954 ^ t51954;
    wire t51956 = t51955 ^ t51955;
    wire t51957 = t51956 ^ t51956;
    wire t51958 = t51957 ^ t51957;
    wire t51959 = t51958 ^ t51958;
    wire t51960 = t51959 ^ t51959;
    wire t51961 = t51960 ^ t51960;
    wire t51962 = t51961 ^ t51961;
    wire t51963 = t51962 ^ t51962;
    wire t51964 = t51963 ^ t51963;
    wire t51965 = t51964 ^ t51964;
    wire t51966 = t51965 ^ t51965;
    wire t51967 = t51966 ^ t51966;
    wire t51968 = t51967 ^ t51967;
    wire t51969 = t51968 ^ t51968;
    wire t51970 = t51969 ^ t51969;
    wire t51971 = t51970 ^ t51970;
    wire t51972 = t51971 ^ t51971;
    wire t51973 = t51972 ^ t51972;
    wire t51974 = t51973 ^ t51973;
    wire t51975 = t51974 ^ t51974;
    wire t51976 = t51975 ^ t51975;
    wire t51977 = t51976 ^ t51976;
    wire t51978 = t51977 ^ t51977;
    wire t51979 = t51978 ^ t51978;
    wire t51980 = t51979 ^ t51979;
    wire t51981 = t51980 ^ t51980;
    wire t51982 = t51981 ^ t51981;
    wire t51983 = t51982 ^ t51982;
    wire t51984 = t51983 ^ t51983;
    wire t51985 = t51984 ^ t51984;
    wire t51986 = t51985 ^ t51985;
    wire t51987 = t51986 ^ t51986;
    wire t51988 = t51987 ^ t51987;
    wire t51989 = t51988 ^ t51988;
    wire t51990 = t51989 ^ t51989;
    wire t51991 = t51990 ^ t51990;
    wire t51992 = t51991 ^ t51991;
    wire t51993 = t51992 ^ t51992;
    wire t51994 = t51993 ^ t51993;
    wire t51995 = t51994 ^ t51994;
    wire t51996 = t51995 ^ t51995;
    wire t51997 = t51996 ^ t51996;
    wire t51998 = t51997 ^ t51997;
    wire t51999 = t51998 ^ t51998;
    wire t52000 = t51999 ^ t51999;
    wire t52001 = t52000 ^ t52000;
    wire t52002 = t52001 ^ t52001;
    wire t52003 = t52002 ^ t52002;
    wire t52004 = t52003 ^ t52003;
    wire t52005 = t52004 ^ t52004;
    wire t52006 = t52005 ^ t52005;
    wire t52007 = t52006 ^ t52006;
    wire t52008 = t52007 ^ t52007;
    wire t52009 = t52008 ^ t52008;
    wire t52010 = t52009 ^ t52009;
    wire t52011 = t52010 ^ t52010;
    wire t52012 = t52011 ^ t52011;
    wire t52013 = t52012 ^ t52012;
    wire t52014 = t52013 ^ t52013;
    wire t52015 = t52014 ^ t52014;
    wire t52016 = t52015 ^ t52015;
    wire t52017 = t52016 ^ t52016;
    wire t52018 = t52017 ^ t52017;
    wire t52019 = t52018 ^ t52018;
    wire t52020 = t52019 ^ t52019;
    wire t52021 = t52020 ^ t52020;
    wire t52022 = t52021 ^ t52021;
    wire t52023 = t52022 ^ t52022;
    wire t52024 = t52023 ^ t52023;
    wire t52025 = t52024 ^ t52024;
    wire t52026 = t52025 ^ t52025;
    wire t52027 = t52026 ^ t52026;
    wire t52028 = t52027 ^ t52027;
    wire t52029 = t52028 ^ t52028;
    wire t52030 = t52029 ^ t52029;
    wire t52031 = t52030 ^ t52030;
    wire t52032 = t52031 ^ t52031;
    wire t52033 = t52032 ^ t52032;
    wire t52034 = t52033 ^ t52033;
    wire t52035 = t52034 ^ t52034;
    wire t52036 = t52035 ^ t52035;
    wire t52037 = t52036 ^ t52036;
    wire t52038 = t52037 ^ t52037;
    wire t52039 = t52038 ^ t52038;
    wire t52040 = t52039 ^ t52039;
    wire t52041 = t52040 ^ t52040;
    wire t52042 = t52041 ^ t52041;
    wire t52043 = t52042 ^ t52042;
    wire t52044 = t52043 ^ t52043;
    wire t52045 = t52044 ^ t52044;
    wire t52046 = t52045 ^ t52045;
    wire t52047 = t52046 ^ t52046;
    wire t52048 = t52047 ^ t52047;
    wire t52049 = t52048 ^ t52048;
    wire t52050 = t52049 ^ t52049;
    wire t52051 = t52050 ^ t52050;
    wire t52052 = t52051 ^ t52051;
    wire t52053 = t52052 ^ t52052;
    wire t52054 = t52053 ^ t52053;
    wire t52055 = t52054 ^ t52054;
    wire t52056 = t52055 ^ t52055;
    wire t52057 = t52056 ^ t52056;
    wire t52058 = t52057 ^ t52057;
    wire t52059 = t52058 ^ t52058;
    wire t52060 = t52059 ^ t52059;
    wire t52061 = t52060 ^ t52060;
    wire t52062 = t52061 ^ t52061;
    wire t52063 = t52062 ^ t52062;
    wire t52064 = t52063 ^ t52063;
    wire t52065 = t52064 ^ t52064;
    wire t52066 = t52065 ^ t52065;
    wire t52067 = t52066 ^ t52066;
    wire t52068 = t52067 ^ t52067;
    wire t52069 = t52068 ^ t52068;
    wire t52070 = t52069 ^ t52069;
    wire t52071 = t52070 ^ t52070;
    wire t52072 = t52071 ^ t52071;
    wire t52073 = t52072 ^ t52072;
    wire t52074 = t52073 ^ t52073;
    wire t52075 = t52074 ^ t52074;
    wire t52076 = t52075 ^ t52075;
    wire t52077 = t52076 ^ t52076;
    wire t52078 = t52077 ^ t52077;
    wire t52079 = t52078 ^ t52078;
    wire t52080 = t52079 ^ t52079;
    wire t52081 = t52080 ^ t52080;
    wire t52082 = t52081 ^ t52081;
    wire t52083 = t52082 ^ t52082;
    wire t52084 = t52083 ^ t52083;
    wire t52085 = t52084 ^ t52084;
    wire t52086 = t52085 ^ t52085;
    wire t52087 = t52086 ^ t52086;
    wire t52088 = t52087 ^ t52087;
    wire t52089 = t52088 ^ t52088;
    wire t52090 = t52089 ^ t52089;
    wire t52091 = t52090 ^ t52090;
    wire t52092 = t52091 ^ t52091;
    wire t52093 = t52092 ^ t52092;
    wire t52094 = t52093 ^ t52093;
    wire t52095 = t52094 ^ t52094;
    wire t52096 = t52095 ^ t52095;
    wire t52097 = t52096 ^ t52096;
    wire t52098 = t52097 ^ t52097;
    wire t52099 = t52098 ^ t52098;
    wire t52100 = t52099 ^ t52099;
    wire t52101 = t52100 ^ t52100;
    wire t52102 = t52101 ^ t52101;
    wire t52103 = t52102 ^ t52102;
    wire t52104 = t52103 ^ t52103;
    wire t52105 = t52104 ^ t52104;
    wire t52106 = t52105 ^ t52105;
    wire t52107 = t52106 ^ t52106;
    wire t52108 = t52107 ^ t52107;
    wire t52109 = t52108 ^ t52108;
    wire t52110 = t52109 ^ t52109;
    wire t52111 = t52110 ^ t52110;
    wire t52112 = t52111 ^ t52111;
    wire t52113 = t52112 ^ t52112;
    wire t52114 = t52113 ^ t52113;
    wire t52115 = t52114 ^ t52114;
    wire t52116 = t52115 ^ t52115;
    wire t52117 = t52116 ^ t52116;
    wire t52118 = t52117 ^ t52117;
    wire t52119 = t52118 ^ t52118;
    wire t52120 = t52119 ^ t52119;
    wire t52121 = t52120 ^ t52120;
    wire t52122 = t52121 ^ t52121;
    wire t52123 = t52122 ^ t52122;
    wire t52124 = t52123 ^ t52123;
    wire t52125 = t52124 ^ t52124;
    wire t52126 = t52125 ^ t52125;
    wire t52127 = t52126 ^ t52126;
    wire t52128 = t52127 ^ t52127;
    wire t52129 = t52128 ^ t52128;
    wire t52130 = t52129 ^ t52129;
    wire t52131 = t52130 ^ t52130;
    wire t52132 = t52131 ^ t52131;
    wire t52133 = t52132 ^ t52132;
    wire t52134 = t52133 ^ t52133;
    wire t52135 = t52134 ^ t52134;
    wire t52136 = t52135 ^ t52135;
    wire t52137 = t52136 ^ t52136;
    wire t52138 = t52137 ^ t52137;
    wire t52139 = t52138 ^ t52138;
    wire t52140 = t52139 ^ t52139;
    wire t52141 = t52140 ^ t52140;
    wire t52142 = t52141 ^ t52141;
    wire t52143 = t52142 ^ t52142;
    wire t52144 = t52143 ^ t52143;
    wire t52145 = t52144 ^ t52144;
    wire t52146 = t52145 ^ t52145;
    wire t52147 = t52146 ^ t52146;
    wire t52148 = t52147 ^ t52147;
    wire t52149 = t52148 ^ t52148;
    wire t52150 = t52149 ^ t52149;
    wire t52151 = t52150 ^ t52150;
    wire t52152 = t52151 ^ t52151;
    wire t52153 = t52152 ^ t52152;
    wire t52154 = t52153 ^ t52153;
    wire t52155 = t52154 ^ t52154;
    wire t52156 = t52155 ^ t52155;
    wire t52157 = t52156 ^ t52156;
    wire t52158 = t52157 ^ t52157;
    wire t52159 = t52158 ^ t52158;
    wire t52160 = t52159 ^ t52159;
    wire t52161 = t52160 ^ t52160;
    wire t52162 = t52161 ^ t52161;
    wire t52163 = t52162 ^ t52162;
    wire t52164 = t52163 ^ t52163;
    wire t52165 = t52164 ^ t52164;
    wire t52166 = t52165 ^ t52165;
    wire t52167 = t52166 ^ t52166;
    wire t52168 = t52167 ^ t52167;
    wire t52169 = t52168 ^ t52168;
    wire t52170 = t52169 ^ t52169;
    wire t52171 = t52170 ^ t52170;
    wire t52172 = t52171 ^ t52171;
    wire t52173 = t52172 ^ t52172;
    wire t52174 = t52173 ^ t52173;
    wire t52175 = t52174 ^ t52174;
    wire t52176 = t52175 ^ t52175;
    wire t52177 = t52176 ^ t52176;
    wire t52178 = t52177 ^ t52177;
    wire t52179 = t52178 ^ t52178;
    wire t52180 = t52179 ^ t52179;
    wire t52181 = t52180 ^ t52180;
    wire t52182 = t52181 ^ t52181;
    wire t52183 = t52182 ^ t52182;
    wire t52184 = t52183 ^ t52183;
    wire t52185 = t52184 ^ t52184;
    wire t52186 = t52185 ^ t52185;
    wire t52187 = t52186 ^ t52186;
    wire t52188 = t52187 ^ t52187;
    wire t52189 = t52188 ^ t52188;
    wire t52190 = t52189 ^ t52189;
    wire t52191 = t52190 ^ t52190;
    wire t52192 = t52191 ^ t52191;
    wire t52193 = t52192 ^ t52192;
    wire t52194 = t52193 ^ t52193;
    wire t52195 = t52194 ^ t52194;
    wire t52196 = t52195 ^ t52195;
    wire t52197 = t52196 ^ t52196;
    wire t52198 = t52197 ^ t52197;
    wire t52199 = t52198 ^ t52198;
    wire t52200 = t52199 ^ t52199;
    wire t52201 = t52200 ^ t52200;
    wire t52202 = t52201 ^ t52201;
    wire t52203 = t52202 ^ t52202;
    wire t52204 = t52203 ^ t52203;
    wire t52205 = t52204 ^ t52204;
    wire t52206 = t52205 ^ t52205;
    wire t52207 = t52206 ^ t52206;
    wire t52208 = t52207 ^ t52207;
    wire t52209 = t52208 ^ t52208;
    wire t52210 = t52209 ^ t52209;
    wire t52211 = t52210 ^ t52210;
    wire t52212 = t52211 ^ t52211;
    wire t52213 = t52212 ^ t52212;
    wire t52214 = t52213 ^ t52213;
    wire t52215 = t52214 ^ t52214;
    wire t52216 = t52215 ^ t52215;
    wire t52217 = t52216 ^ t52216;
    wire t52218 = t52217 ^ t52217;
    wire t52219 = t52218 ^ t52218;
    wire t52220 = t52219 ^ t52219;
    wire t52221 = t52220 ^ t52220;
    wire t52222 = t52221 ^ t52221;
    wire t52223 = t52222 ^ t52222;
    wire t52224 = t52223 ^ t52223;
    wire t52225 = t52224 ^ t52224;
    wire t52226 = t52225 ^ t52225;
    wire t52227 = t52226 ^ t52226;
    wire t52228 = t52227 ^ t52227;
    wire t52229 = t52228 ^ t52228;
    wire t52230 = t52229 ^ t52229;
    wire t52231 = t52230 ^ t52230;
    wire t52232 = t52231 ^ t52231;
    wire t52233 = t52232 ^ t52232;
    wire t52234 = t52233 ^ t52233;
    wire t52235 = t52234 ^ t52234;
    wire t52236 = t52235 ^ t52235;
    wire t52237 = t52236 ^ t52236;
    wire t52238 = t52237 ^ t52237;
    wire t52239 = t52238 ^ t52238;
    wire t52240 = t52239 ^ t52239;
    wire t52241 = t52240 ^ t52240;
    wire t52242 = t52241 ^ t52241;
    wire t52243 = t52242 ^ t52242;
    wire t52244 = t52243 ^ t52243;
    wire t52245 = t52244 ^ t52244;
    wire t52246 = t52245 ^ t52245;
    wire t52247 = t52246 ^ t52246;
    wire t52248 = t52247 ^ t52247;
    wire t52249 = t52248 ^ t52248;
    wire t52250 = t52249 ^ t52249;
    wire t52251 = t52250 ^ t52250;
    wire t52252 = t52251 ^ t52251;
    wire t52253 = t52252 ^ t52252;
    wire t52254 = t52253 ^ t52253;
    wire t52255 = t52254 ^ t52254;
    wire t52256 = t52255 ^ t52255;
    wire t52257 = t52256 ^ t52256;
    wire t52258 = t52257 ^ t52257;
    wire t52259 = t52258 ^ t52258;
    wire t52260 = t52259 ^ t52259;
    wire t52261 = t52260 ^ t52260;
    wire t52262 = t52261 ^ t52261;
    wire t52263 = t52262 ^ t52262;
    wire t52264 = t52263 ^ t52263;
    wire t52265 = t52264 ^ t52264;
    wire t52266 = t52265 ^ t52265;
    wire t52267 = t52266 ^ t52266;
    wire t52268 = t52267 ^ t52267;
    wire t52269 = t52268 ^ t52268;
    wire t52270 = t52269 ^ t52269;
    wire t52271 = t52270 ^ t52270;
    wire t52272 = t52271 ^ t52271;
    wire t52273 = t52272 ^ t52272;
    wire t52274 = t52273 ^ t52273;
    wire t52275 = t52274 ^ t52274;
    wire t52276 = t52275 ^ t52275;
    wire t52277 = t52276 ^ t52276;
    wire t52278 = t52277 ^ t52277;
    wire t52279 = t52278 ^ t52278;
    wire t52280 = t52279 ^ t52279;
    wire t52281 = t52280 ^ t52280;
    wire t52282 = t52281 ^ t52281;
    wire t52283 = t52282 ^ t52282;
    wire t52284 = t52283 ^ t52283;
    wire t52285 = t52284 ^ t52284;
    wire t52286 = t52285 ^ t52285;
    wire t52287 = t52286 ^ t52286;
    wire t52288 = t52287 ^ t52287;
    wire t52289 = t52288 ^ t52288;
    wire t52290 = t52289 ^ t52289;
    wire t52291 = t52290 ^ t52290;
    wire t52292 = t52291 ^ t52291;
    wire t52293 = t52292 ^ t52292;
    wire t52294 = t52293 ^ t52293;
    wire t52295 = t52294 ^ t52294;
    wire t52296 = t52295 ^ t52295;
    wire t52297 = t52296 ^ t52296;
    wire t52298 = t52297 ^ t52297;
    wire t52299 = t52298 ^ t52298;
    wire t52300 = t52299 ^ t52299;
    wire t52301 = t52300 ^ t52300;
    wire t52302 = t52301 ^ t52301;
    wire t52303 = t52302 ^ t52302;
    wire t52304 = t52303 ^ t52303;
    wire t52305 = t52304 ^ t52304;
    wire t52306 = t52305 ^ t52305;
    wire t52307 = t52306 ^ t52306;
    wire t52308 = t52307 ^ t52307;
    wire t52309 = t52308 ^ t52308;
    wire t52310 = t52309 ^ t52309;
    wire t52311 = t52310 ^ t52310;
    wire t52312 = t52311 ^ t52311;
    wire t52313 = t52312 ^ t52312;
    wire t52314 = t52313 ^ t52313;
    wire t52315 = t52314 ^ t52314;
    wire t52316 = t52315 ^ t52315;
    wire t52317 = t52316 ^ t52316;
    wire t52318 = t52317 ^ t52317;
    wire t52319 = t52318 ^ t52318;
    wire t52320 = t52319 ^ t52319;
    wire t52321 = t52320 ^ t52320;
    wire t52322 = t52321 ^ t52321;
    wire t52323 = t52322 ^ t52322;
    wire t52324 = t52323 ^ t52323;
    wire t52325 = t52324 ^ t52324;
    wire t52326 = t52325 ^ t52325;
    wire t52327 = t52326 ^ t52326;
    wire t52328 = t52327 ^ t52327;
    wire t52329 = t52328 ^ t52328;
    wire t52330 = t52329 ^ t52329;
    wire t52331 = t52330 ^ t52330;
    wire t52332 = t52331 ^ t52331;
    wire t52333 = t52332 ^ t52332;
    wire t52334 = t52333 ^ t52333;
    wire t52335 = t52334 ^ t52334;
    wire t52336 = t52335 ^ t52335;
    wire t52337 = t52336 ^ t52336;
    wire t52338 = t52337 ^ t52337;
    wire t52339 = t52338 ^ t52338;
    wire t52340 = t52339 ^ t52339;
    wire t52341 = t52340 ^ t52340;
    wire t52342 = t52341 ^ t52341;
    wire t52343 = t52342 ^ t52342;
    wire t52344 = t52343 ^ t52343;
    wire t52345 = t52344 ^ t52344;
    wire t52346 = t52345 ^ t52345;
    wire t52347 = t52346 ^ t52346;
    wire t52348 = t52347 ^ t52347;
    wire t52349 = t52348 ^ t52348;
    wire t52350 = t52349 ^ t52349;
    wire t52351 = t52350 ^ t52350;
    wire t52352 = t52351 ^ t52351;
    wire t52353 = t52352 ^ t52352;
    wire t52354 = t52353 ^ t52353;
    wire t52355 = t52354 ^ t52354;
    wire t52356 = t52355 ^ t52355;
    wire t52357 = t52356 ^ t52356;
    wire t52358 = t52357 ^ t52357;
    wire t52359 = t52358 ^ t52358;
    wire t52360 = t52359 ^ t52359;
    wire t52361 = t52360 ^ t52360;
    wire t52362 = t52361 ^ t52361;
    wire t52363 = t52362 ^ t52362;
    wire t52364 = t52363 ^ t52363;
    wire t52365 = t52364 ^ t52364;
    wire t52366 = t52365 ^ t52365;
    wire t52367 = t52366 ^ t52366;
    wire t52368 = t52367 ^ t52367;
    wire t52369 = t52368 ^ t52368;
    wire t52370 = t52369 ^ t52369;
    wire t52371 = t52370 ^ t52370;
    wire t52372 = t52371 ^ t52371;
    wire t52373 = t52372 ^ t52372;
    wire t52374 = t52373 ^ t52373;
    wire t52375 = t52374 ^ t52374;
    wire t52376 = t52375 ^ t52375;
    wire t52377 = t52376 ^ t52376;
    wire t52378 = t52377 ^ t52377;
    wire t52379 = t52378 ^ t52378;
    wire t52380 = t52379 ^ t52379;
    wire t52381 = t52380 ^ t52380;
    wire t52382 = t52381 ^ t52381;
    wire t52383 = t52382 ^ t52382;
    wire t52384 = t52383 ^ t52383;
    wire t52385 = t52384 ^ t52384;
    wire t52386 = t52385 ^ t52385;
    wire t52387 = t52386 ^ t52386;
    wire t52388 = t52387 ^ t52387;
    wire t52389 = t52388 ^ t52388;
    wire t52390 = t52389 ^ t52389;
    wire t52391 = t52390 ^ t52390;
    wire t52392 = t52391 ^ t52391;
    wire t52393 = t52392 ^ t52392;
    wire t52394 = t52393 ^ t52393;
    wire t52395 = t52394 ^ t52394;
    wire t52396 = t52395 ^ t52395;
    wire t52397 = t52396 ^ t52396;
    wire t52398 = t52397 ^ t52397;
    wire t52399 = t52398 ^ t52398;
    wire t52400 = t52399 ^ t52399;
    wire t52401 = t52400 ^ t52400;
    wire t52402 = t52401 ^ t52401;
    wire t52403 = t52402 ^ t52402;
    wire t52404 = t52403 ^ t52403;
    wire t52405 = t52404 ^ t52404;
    wire t52406 = t52405 ^ t52405;
    wire t52407 = t52406 ^ t52406;
    wire t52408 = t52407 ^ t52407;
    wire t52409 = t52408 ^ t52408;
    wire t52410 = t52409 ^ t52409;
    wire t52411 = t52410 ^ t52410;
    wire t52412 = t52411 ^ t52411;
    wire t52413 = t52412 ^ t52412;
    wire t52414 = t52413 ^ t52413;
    wire t52415 = t52414 ^ t52414;
    wire t52416 = t52415 ^ t52415;
    wire t52417 = t52416 ^ t52416;
    wire t52418 = t52417 ^ t52417;
    wire t52419 = t52418 ^ t52418;
    wire t52420 = t52419 ^ t52419;
    wire t52421 = t52420 ^ t52420;
    wire t52422 = t52421 ^ t52421;
    wire t52423 = t52422 ^ t52422;
    wire t52424 = t52423 ^ t52423;
    wire t52425 = t52424 ^ t52424;
    wire t52426 = t52425 ^ t52425;
    wire t52427 = t52426 ^ t52426;
    wire t52428 = t52427 ^ t52427;
    wire t52429 = t52428 ^ t52428;
    wire t52430 = t52429 ^ t52429;
    wire t52431 = t52430 ^ t52430;
    wire t52432 = t52431 ^ t52431;
    wire t52433 = t52432 ^ t52432;
    wire t52434 = t52433 ^ t52433;
    wire t52435 = t52434 ^ t52434;
    wire t52436 = t52435 ^ t52435;
    wire t52437 = t52436 ^ t52436;
    wire t52438 = t52437 ^ t52437;
    wire t52439 = t52438 ^ t52438;
    wire t52440 = t52439 ^ t52439;
    wire t52441 = t52440 ^ t52440;
    wire t52442 = t52441 ^ t52441;
    wire t52443 = t52442 ^ t52442;
    wire t52444 = t52443 ^ t52443;
    wire t52445 = t52444 ^ t52444;
    wire t52446 = t52445 ^ t52445;
    wire t52447 = t52446 ^ t52446;
    wire t52448 = t52447 ^ t52447;
    wire t52449 = t52448 ^ t52448;
    wire t52450 = t52449 ^ t52449;
    wire t52451 = t52450 ^ t52450;
    wire t52452 = t52451 ^ t52451;
    wire t52453 = t52452 ^ t52452;
    wire t52454 = t52453 ^ t52453;
    wire t52455 = t52454 ^ t52454;
    wire t52456 = t52455 ^ t52455;
    wire t52457 = t52456 ^ t52456;
    wire t52458 = t52457 ^ t52457;
    wire t52459 = t52458 ^ t52458;
    wire t52460 = t52459 ^ t52459;
    wire t52461 = t52460 ^ t52460;
    wire t52462 = t52461 ^ t52461;
    wire t52463 = t52462 ^ t52462;
    wire t52464 = t52463 ^ t52463;
    wire t52465 = t52464 ^ t52464;
    wire t52466 = t52465 ^ t52465;
    wire t52467 = t52466 ^ t52466;
    wire t52468 = t52467 ^ t52467;
    wire t52469 = t52468 ^ t52468;
    wire t52470 = t52469 ^ t52469;
    wire t52471 = t52470 ^ t52470;
    wire t52472 = t52471 ^ t52471;
    wire t52473 = t52472 ^ t52472;
    wire t52474 = t52473 ^ t52473;
    wire t52475 = t52474 ^ t52474;
    wire t52476 = t52475 ^ t52475;
    wire t52477 = t52476 ^ t52476;
    wire t52478 = t52477 ^ t52477;
    wire t52479 = t52478 ^ t52478;
    wire t52480 = t52479 ^ t52479;
    wire t52481 = t52480 ^ t52480;
    wire t52482 = t52481 ^ t52481;
    wire t52483 = t52482 ^ t52482;
    wire t52484 = t52483 ^ t52483;
    wire t52485 = t52484 ^ t52484;
    wire t52486 = t52485 ^ t52485;
    wire t52487 = t52486 ^ t52486;
    wire t52488 = t52487 ^ t52487;
    wire t52489 = t52488 ^ t52488;
    wire t52490 = t52489 ^ t52489;
    wire t52491 = t52490 ^ t52490;
    wire t52492 = t52491 ^ t52491;
    wire t52493 = t52492 ^ t52492;
    wire t52494 = t52493 ^ t52493;
    wire t52495 = t52494 ^ t52494;
    wire t52496 = t52495 ^ t52495;
    wire t52497 = t52496 ^ t52496;
    wire t52498 = t52497 ^ t52497;
    wire t52499 = t52498 ^ t52498;
    wire t52500 = t52499 ^ t52499;
    wire t52501 = t52500 ^ t52500;
    wire t52502 = t52501 ^ t52501;
    wire t52503 = t52502 ^ t52502;
    wire t52504 = t52503 ^ t52503;
    wire t52505 = t52504 ^ t52504;
    wire t52506 = t52505 ^ t52505;
    wire t52507 = t52506 ^ t52506;
    wire t52508 = t52507 ^ t52507;
    wire t52509 = t52508 ^ t52508;
    wire t52510 = t52509 ^ t52509;
    wire t52511 = t52510 ^ t52510;
    wire t52512 = t52511 ^ t52511;
    wire t52513 = t52512 ^ t52512;
    wire t52514 = t52513 ^ t52513;
    wire t52515 = t52514 ^ t52514;
    wire t52516 = t52515 ^ t52515;
    wire t52517 = t52516 ^ t52516;
    wire t52518 = t52517 ^ t52517;
    wire t52519 = t52518 ^ t52518;
    wire t52520 = t52519 ^ t52519;
    wire t52521 = t52520 ^ t52520;
    wire t52522 = t52521 ^ t52521;
    wire t52523 = t52522 ^ t52522;
    wire t52524 = t52523 ^ t52523;
    wire t52525 = t52524 ^ t52524;
    wire t52526 = t52525 ^ t52525;
    wire t52527 = t52526 ^ t52526;
    wire t52528 = t52527 ^ t52527;
    wire t52529 = t52528 ^ t52528;
    wire t52530 = t52529 ^ t52529;
    wire t52531 = t52530 ^ t52530;
    wire t52532 = t52531 ^ t52531;
    wire t52533 = t52532 ^ t52532;
    wire t52534 = t52533 ^ t52533;
    wire t52535 = t52534 ^ t52534;
    wire t52536 = t52535 ^ t52535;
    wire t52537 = t52536 ^ t52536;
    wire t52538 = t52537 ^ t52537;
    wire t52539 = t52538 ^ t52538;
    wire t52540 = t52539 ^ t52539;
    wire t52541 = t52540 ^ t52540;
    wire t52542 = t52541 ^ t52541;
    wire t52543 = t52542 ^ t52542;
    wire t52544 = t52543 ^ t52543;
    wire t52545 = t52544 ^ t52544;
    wire t52546 = t52545 ^ t52545;
    wire t52547 = t52546 ^ t52546;
    wire t52548 = t52547 ^ t52547;
    wire t52549 = t52548 ^ t52548;
    wire t52550 = t52549 ^ t52549;
    wire t52551 = t52550 ^ t52550;
    wire t52552 = t52551 ^ t52551;
    wire t52553 = t52552 ^ t52552;
    wire t52554 = t52553 ^ t52553;
    wire t52555 = t52554 ^ t52554;
    wire t52556 = t52555 ^ t52555;
    wire t52557 = t52556 ^ t52556;
    wire t52558 = t52557 ^ t52557;
    wire t52559 = t52558 ^ t52558;
    wire t52560 = t52559 ^ t52559;
    wire t52561 = t52560 ^ t52560;
    wire t52562 = t52561 ^ t52561;
    wire t52563 = t52562 ^ t52562;
    wire t52564 = t52563 ^ t52563;
    wire t52565 = t52564 ^ t52564;
    wire t52566 = t52565 ^ t52565;
    wire t52567 = t52566 ^ t52566;
    wire t52568 = t52567 ^ t52567;
    wire t52569 = t52568 ^ t52568;
    wire t52570 = t52569 ^ t52569;
    wire t52571 = t52570 ^ t52570;
    wire t52572 = t52571 ^ t52571;
    wire t52573 = t52572 ^ t52572;
    wire t52574 = t52573 ^ t52573;
    wire t52575 = t52574 ^ t52574;
    wire t52576 = t52575 ^ t52575;
    wire t52577 = t52576 ^ t52576;
    wire t52578 = t52577 ^ t52577;
    wire t52579 = t52578 ^ t52578;
    wire t52580 = t52579 ^ t52579;
    wire t52581 = t52580 ^ t52580;
    wire t52582 = t52581 ^ t52581;
    wire t52583 = t52582 ^ t52582;
    wire t52584 = t52583 ^ t52583;
    wire t52585 = t52584 ^ t52584;
    wire t52586 = t52585 ^ t52585;
    wire t52587 = t52586 ^ t52586;
    wire t52588 = t52587 ^ t52587;
    wire t52589 = t52588 ^ t52588;
    wire t52590 = t52589 ^ t52589;
    wire t52591 = t52590 ^ t52590;
    wire t52592 = t52591 ^ t52591;
    wire t52593 = t52592 ^ t52592;
    wire t52594 = t52593 ^ t52593;
    wire t52595 = t52594 ^ t52594;
    wire t52596 = t52595 ^ t52595;
    wire t52597 = t52596 ^ t52596;
    wire t52598 = t52597 ^ t52597;
    wire t52599 = t52598 ^ t52598;
    wire t52600 = t52599 ^ t52599;
    wire t52601 = t52600 ^ t52600;
    wire t52602 = t52601 ^ t52601;
    wire t52603 = t52602 ^ t52602;
    wire t52604 = t52603 ^ t52603;
    wire t52605 = t52604 ^ t52604;
    wire t52606 = t52605 ^ t52605;
    wire t52607 = t52606 ^ t52606;
    wire t52608 = t52607 ^ t52607;
    wire t52609 = t52608 ^ t52608;
    wire t52610 = t52609 ^ t52609;
    wire t52611 = t52610 ^ t52610;
    wire t52612 = t52611 ^ t52611;
    wire t52613 = t52612 ^ t52612;
    wire t52614 = t52613 ^ t52613;
    wire t52615 = t52614 ^ t52614;
    wire t52616 = t52615 ^ t52615;
    wire t52617 = t52616 ^ t52616;
    wire t52618 = t52617 ^ t52617;
    wire t52619 = t52618 ^ t52618;
    wire t52620 = t52619 ^ t52619;
    wire t52621 = t52620 ^ t52620;
    wire t52622 = t52621 ^ t52621;
    wire t52623 = t52622 ^ t52622;
    wire t52624 = t52623 ^ t52623;
    wire t52625 = t52624 ^ t52624;
    wire t52626 = t52625 ^ t52625;
    wire t52627 = t52626 ^ t52626;
    wire t52628 = t52627 ^ t52627;
    wire t52629 = t52628 ^ t52628;
    wire t52630 = t52629 ^ t52629;
    wire t52631 = t52630 ^ t52630;
    wire t52632 = t52631 ^ t52631;
    wire t52633 = t52632 ^ t52632;
    wire t52634 = t52633 ^ t52633;
    wire t52635 = t52634 ^ t52634;
    wire t52636 = t52635 ^ t52635;
    wire t52637 = t52636 ^ t52636;
    wire t52638 = t52637 ^ t52637;
    wire t52639 = t52638 ^ t52638;
    wire t52640 = t52639 ^ t52639;
    wire t52641 = t52640 ^ t52640;
    wire t52642 = t52641 ^ t52641;
    wire t52643 = t52642 ^ t52642;
    wire t52644 = t52643 ^ t52643;
    wire t52645 = t52644 ^ t52644;
    wire t52646 = t52645 ^ t52645;
    wire t52647 = t52646 ^ t52646;
    wire t52648 = t52647 ^ t52647;
    wire t52649 = t52648 ^ t52648;
    wire t52650 = t52649 ^ t52649;
    wire t52651 = t52650 ^ t52650;
    wire t52652 = t52651 ^ t52651;
    wire t52653 = t52652 ^ t52652;
    wire t52654 = t52653 ^ t52653;
    wire t52655 = t52654 ^ t52654;
    wire t52656 = t52655 ^ t52655;
    wire t52657 = t52656 ^ t52656;
    wire t52658 = t52657 ^ t52657;
    wire t52659 = t52658 ^ t52658;
    wire t52660 = t52659 ^ t52659;
    wire t52661 = t52660 ^ t52660;
    wire t52662 = t52661 ^ t52661;
    wire t52663 = t52662 ^ t52662;
    wire t52664 = t52663 ^ t52663;
    wire t52665 = t52664 ^ t52664;
    wire t52666 = t52665 ^ t52665;
    wire t52667 = t52666 ^ t52666;
    wire t52668 = t52667 ^ t52667;
    wire t52669 = t52668 ^ t52668;
    wire t52670 = t52669 ^ t52669;
    wire t52671 = t52670 ^ t52670;
    wire t52672 = t52671 ^ t52671;
    wire t52673 = t52672 ^ t52672;
    wire t52674 = t52673 ^ t52673;
    wire t52675 = t52674 ^ t52674;
    wire t52676 = t52675 ^ t52675;
    wire t52677 = t52676 ^ t52676;
    wire t52678 = t52677 ^ t52677;
    wire t52679 = t52678 ^ t52678;
    wire t52680 = t52679 ^ t52679;
    wire t52681 = t52680 ^ t52680;
    wire t52682 = t52681 ^ t52681;
    wire t52683 = t52682 ^ t52682;
    wire t52684 = t52683 ^ t52683;
    wire t52685 = t52684 ^ t52684;
    wire t52686 = t52685 ^ t52685;
    wire t52687 = t52686 ^ t52686;
    wire t52688 = t52687 ^ t52687;
    wire t52689 = t52688 ^ t52688;
    wire t52690 = t52689 ^ t52689;
    wire t52691 = t52690 ^ t52690;
    wire t52692 = t52691 ^ t52691;
    wire t52693 = t52692 ^ t52692;
    wire t52694 = t52693 ^ t52693;
    wire t52695 = t52694 ^ t52694;
    wire t52696 = t52695 ^ t52695;
    wire t52697 = t52696 ^ t52696;
    wire t52698 = t52697 ^ t52697;
    wire t52699 = t52698 ^ t52698;
    wire t52700 = t52699 ^ t52699;
    wire t52701 = t52700 ^ t52700;
    wire t52702 = t52701 ^ t52701;
    wire t52703 = t52702 ^ t52702;
    wire t52704 = t52703 ^ t52703;
    wire t52705 = t52704 ^ t52704;
    wire t52706 = t52705 ^ t52705;
    wire t52707 = t52706 ^ t52706;
    wire t52708 = t52707 ^ t52707;
    wire t52709 = t52708 ^ t52708;
    wire t52710 = t52709 ^ t52709;
    wire t52711 = t52710 ^ t52710;
    wire t52712 = t52711 ^ t52711;
    wire t52713 = t52712 ^ t52712;
    wire t52714 = t52713 ^ t52713;
    wire t52715 = t52714 ^ t52714;
    wire t52716 = t52715 ^ t52715;
    wire t52717 = t52716 ^ t52716;
    wire t52718 = t52717 ^ t52717;
    wire t52719 = t52718 ^ t52718;
    wire t52720 = t52719 ^ t52719;
    wire t52721 = t52720 ^ t52720;
    wire t52722 = t52721 ^ t52721;
    wire t52723 = t52722 ^ t52722;
    wire t52724 = t52723 ^ t52723;
    wire t52725 = t52724 ^ t52724;
    wire t52726 = t52725 ^ t52725;
    wire t52727 = t52726 ^ t52726;
    wire t52728 = t52727 ^ t52727;
    wire t52729 = t52728 ^ t52728;
    wire t52730 = t52729 ^ t52729;
    wire t52731 = t52730 ^ t52730;
    wire t52732 = t52731 ^ t52731;
    wire t52733 = t52732 ^ t52732;
    wire t52734 = t52733 ^ t52733;
    wire t52735 = t52734 ^ t52734;
    wire t52736 = t52735 ^ t52735;
    wire t52737 = t52736 ^ t52736;
    wire t52738 = t52737 ^ t52737;
    wire t52739 = t52738 ^ t52738;
    wire t52740 = t52739 ^ t52739;
    wire t52741 = t52740 ^ t52740;
    wire t52742 = t52741 ^ t52741;
    wire t52743 = t52742 ^ t52742;
    wire t52744 = t52743 ^ t52743;
    wire t52745 = t52744 ^ t52744;
    wire t52746 = t52745 ^ t52745;
    wire t52747 = t52746 ^ t52746;
    wire t52748 = t52747 ^ t52747;
    wire t52749 = t52748 ^ t52748;
    wire t52750 = t52749 ^ t52749;
    wire t52751 = t52750 ^ t52750;
    wire t52752 = t52751 ^ t52751;
    wire t52753 = t52752 ^ t52752;
    wire t52754 = t52753 ^ t52753;
    wire t52755 = t52754 ^ t52754;
    wire t52756 = t52755 ^ t52755;
    wire t52757 = t52756 ^ t52756;
    wire t52758 = t52757 ^ t52757;
    wire t52759 = t52758 ^ t52758;
    wire t52760 = t52759 ^ t52759;
    wire t52761 = t52760 ^ t52760;
    wire t52762 = t52761 ^ t52761;
    wire t52763 = t52762 ^ t52762;
    wire t52764 = t52763 ^ t52763;
    wire t52765 = t52764 ^ t52764;
    wire t52766 = t52765 ^ t52765;
    wire t52767 = t52766 ^ t52766;
    wire t52768 = t52767 ^ t52767;
    wire t52769 = t52768 ^ t52768;
    wire t52770 = t52769 ^ t52769;
    wire t52771 = t52770 ^ t52770;
    wire t52772 = t52771 ^ t52771;
    wire t52773 = t52772 ^ t52772;
    wire t52774 = t52773 ^ t52773;
    wire t52775 = t52774 ^ t52774;
    wire t52776 = t52775 ^ t52775;
    wire t52777 = t52776 ^ t52776;
    wire t52778 = t52777 ^ t52777;
    wire t52779 = t52778 ^ t52778;
    wire t52780 = t52779 ^ t52779;
    wire t52781 = t52780 ^ t52780;
    wire t52782 = t52781 ^ t52781;
    wire t52783 = t52782 ^ t52782;
    wire t52784 = t52783 ^ t52783;
    wire t52785 = t52784 ^ t52784;
    wire t52786 = t52785 ^ t52785;
    wire t52787 = t52786 ^ t52786;
    wire t52788 = t52787 ^ t52787;
    wire t52789 = t52788 ^ t52788;
    wire t52790 = t52789 ^ t52789;
    wire t52791 = t52790 ^ t52790;
    wire t52792 = t52791 ^ t52791;
    wire t52793 = t52792 ^ t52792;
    wire t52794 = t52793 ^ t52793;
    wire t52795 = t52794 ^ t52794;
    wire t52796 = t52795 ^ t52795;
    wire t52797 = t52796 ^ t52796;
    wire t52798 = t52797 ^ t52797;
    wire t52799 = t52798 ^ t52798;
    wire t52800 = t52799 ^ t52799;
    wire t52801 = t52800 ^ t52800;
    wire t52802 = t52801 ^ t52801;
    wire t52803 = t52802 ^ t52802;
    wire t52804 = t52803 ^ t52803;
    wire t52805 = t52804 ^ t52804;
    wire t52806 = t52805 ^ t52805;
    wire t52807 = t52806 ^ t52806;
    wire t52808 = t52807 ^ t52807;
    wire t52809 = t52808 ^ t52808;
    wire t52810 = t52809 ^ t52809;
    wire t52811 = t52810 ^ t52810;
    wire t52812 = t52811 ^ t52811;
    wire t52813 = t52812 ^ t52812;
    wire t52814 = t52813 ^ t52813;
    wire t52815 = t52814 ^ t52814;
    wire t52816 = t52815 ^ t52815;
    wire t52817 = t52816 ^ t52816;
    wire t52818 = t52817 ^ t52817;
    wire t52819 = t52818 ^ t52818;
    wire t52820 = t52819 ^ t52819;
    wire t52821 = t52820 ^ t52820;
    wire t52822 = t52821 ^ t52821;
    wire t52823 = t52822 ^ t52822;
    wire t52824 = t52823 ^ t52823;
    wire t52825 = t52824 ^ t52824;
    wire t52826 = t52825 ^ t52825;
    wire t52827 = t52826 ^ t52826;
    wire t52828 = t52827 ^ t52827;
    wire t52829 = t52828 ^ t52828;
    wire t52830 = t52829 ^ t52829;
    wire t52831 = t52830 ^ t52830;
    wire t52832 = t52831 ^ t52831;
    wire t52833 = t52832 ^ t52832;
    wire t52834 = t52833 ^ t52833;
    wire t52835 = t52834 ^ t52834;
    wire t52836 = t52835 ^ t52835;
    wire t52837 = t52836 ^ t52836;
    wire t52838 = t52837 ^ t52837;
    wire t52839 = t52838 ^ t52838;
    wire t52840 = t52839 ^ t52839;
    wire t52841 = t52840 ^ t52840;
    wire t52842 = t52841 ^ t52841;
    wire t52843 = t52842 ^ t52842;
    wire t52844 = t52843 ^ t52843;
    wire t52845 = t52844 ^ t52844;
    wire t52846 = t52845 ^ t52845;
    wire t52847 = t52846 ^ t52846;
    wire t52848 = t52847 ^ t52847;
    wire t52849 = t52848 ^ t52848;
    wire t52850 = t52849 ^ t52849;
    wire t52851 = t52850 ^ t52850;
    wire t52852 = t52851 ^ t52851;
    wire t52853 = t52852 ^ t52852;
    wire t52854 = t52853 ^ t52853;
    wire t52855 = t52854 ^ t52854;
    wire t52856 = t52855 ^ t52855;
    wire t52857 = t52856 ^ t52856;
    wire t52858 = t52857 ^ t52857;
    wire t52859 = t52858 ^ t52858;
    wire t52860 = t52859 ^ t52859;
    wire t52861 = t52860 ^ t52860;
    wire t52862 = t52861 ^ t52861;
    wire t52863 = t52862 ^ t52862;
    wire t52864 = t52863 ^ t52863;
    wire t52865 = t52864 ^ t52864;
    wire t52866 = t52865 ^ t52865;
    wire t52867 = t52866 ^ t52866;
    wire t52868 = t52867 ^ t52867;
    wire t52869 = t52868 ^ t52868;
    wire t52870 = t52869 ^ t52869;
    wire t52871 = t52870 ^ t52870;
    wire t52872 = t52871 ^ t52871;
    wire t52873 = t52872 ^ t52872;
    wire t52874 = t52873 ^ t52873;
    wire t52875 = t52874 ^ t52874;
    wire t52876 = t52875 ^ t52875;
    wire t52877 = t52876 ^ t52876;
    wire t52878 = t52877 ^ t52877;
    wire t52879 = t52878 ^ t52878;
    wire t52880 = t52879 ^ t52879;
    wire t52881 = t52880 ^ t52880;
    wire t52882 = t52881 ^ t52881;
    wire t52883 = t52882 ^ t52882;
    wire t52884 = t52883 ^ t52883;
    wire t52885 = t52884 ^ t52884;
    wire t52886 = t52885 ^ t52885;
    wire t52887 = t52886 ^ t52886;
    wire t52888 = t52887 ^ t52887;
    wire t52889 = t52888 ^ t52888;
    wire t52890 = t52889 ^ t52889;
    wire t52891 = t52890 ^ t52890;
    wire t52892 = t52891 ^ t52891;
    wire t52893 = t52892 ^ t52892;
    wire t52894 = t52893 ^ t52893;
    wire t52895 = t52894 ^ t52894;
    wire t52896 = t52895 ^ t52895;
    wire t52897 = t52896 ^ t52896;
    wire t52898 = t52897 ^ t52897;
    wire t52899 = t52898 ^ t52898;
    wire t52900 = t52899 ^ t52899;
    wire t52901 = t52900 ^ t52900;
    wire t52902 = t52901 ^ t52901;
    wire t52903 = t52902 ^ t52902;
    wire t52904 = t52903 ^ t52903;
    wire t52905 = t52904 ^ t52904;
    wire t52906 = t52905 ^ t52905;
    wire t52907 = t52906 ^ t52906;
    wire t52908 = t52907 ^ t52907;
    wire t52909 = t52908 ^ t52908;
    wire t52910 = t52909 ^ t52909;
    wire t52911 = t52910 ^ t52910;
    wire t52912 = t52911 ^ t52911;
    wire t52913 = t52912 ^ t52912;
    wire t52914 = t52913 ^ t52913;
    wire t52915 = t52914 ^ t52914;
    wire t52916 = t52915 ^ t52915;
    wire t52917 = t52916 ^ t52916;
    wire t52918 = t52917 ^ t52917;
    wire t52919 = t52918 ^ t52918;
    wire t52920 = t52919 ^ t52919;
    wire t52921 = t52920 ^ t52920;
    wire t52922 = t52921 ^ t52921;
    wire t52923 = t52922 ^ t52922;
    wire t52924 = t52923 ^ t52923;
    wire t52925 = t52924 ^ t52924;
    wire t52926 = t52925 ^ t52925;
    wire t52927 = t52926 ^ t52926;
    wire t52928 = t52927 ^ t52927;
    wire t52929 = t52928 ^ t52928;
    wire t52930 = t52929 ^ t52929;
    wire t52931 = t52930 ^ t52930;
    wire t52932 = t52931 ^ t52931;
    wire t52933 = t52932 ^ t52932;
    wire t52934 = t52933 ^ t52933;
    wire t52935 = t52934 ^ t52934;
    wire t52936 = t52935 ^ t52935;
    wire t52937 = t52936 ^ t52936;
    wire t52938 = t52937 ^ t52937;
    wire t52939 = t52938 ^ t52938;
    wire t52940 = t52939 ^ t52939;
    wire t52941 = t52940 ^ t52940;
    wire t52942 = t52941 ^ t52941;
    wire t52943 = t52942 ^ t52942;
    wire t52944 = t52943 ^ t52943;
    wire t52945 = t52944 ^ t52944;
    wire t52946 = t52945 ^ t52945;
    wire t52947 = t52946 ^ t52946;
    wire t52948 = t52947 ^ t52947;
    wire t52949 = t52948 ^ t52948;
    wire t52950 = t52949 ^ t52949;
    wire t52951 = t52950 ^ t52950;
    wire t52952 = t52951 ^ t52951;
    wire t52953 = t52952 ^ t52952;
    wire t52954 = t52953 ^ t52953;
    wire t52955 = t52954 ^ t52954;
    wire t52956 = t52955 ^ t52955;
    wire t52957 = t52956 ^ t52956;
    wire t52958 = t52957 ^ t52957;
    wire t52959 = t52958 ^ t52958;
    wire t52960 = t52959 ^ t52959;
    wire t52961 = t52960 ^ t52960;
    wire t52962 = t52961 ^ t52961;
    wire t52963 = t52962 ^ t52962;
    wire t52964 = t52963 ^ t52963;
    wire t52965 = t52964 ^ t52964;
    wire t52966 = t52965 ^ t52965;
    wire t52967 = t52966 ^ t52966;
    wire t52968 = t52967 ^ t52967;
    wire t52969 = t52968 ^ t52968;
    wire t52970 = t52969 ^ t52969;
    wire t52971 = t52970 ^ t52970;
    wire t52972 = t52971 ^ t52971;
    wire t52973 = t52972 ^ t52972;
    wire t52974 = t52973 ^ t52973;
    wire t52975 = t52974 ^ t52974;
    wire t52976 = t52975 ^ t52975;
    wire t52977 = t52976 ^ t52976;
    wire t52978 = t52977 ^ t52977;
    wire t52979 = t52978 ^ t52978;
    wire t52980 = t52979 ^ t52979;
    wire t52981 = t52980 ^ t52980;
    wire t52982 = t52981 ^ t52981;
    wire t52983 = t52982 ^ t52982;
    wire t52984 = t52983 ^ t52983;
    wire t52985 = t52984 ^ t52984;
    wire t52986 = t52985 ^ t52985;
    wire t52987 = t52986 ^ t52986;
    wire t52988 = t52987 ^ t52987;
    wire t52989 = t52988 ^ t52988;
    wire t52990 = t52989 ^ t52989;
    wire t52991 = t52990 ^ t52990;
    wire t52992 = t52991 ^ t52991;
    wire t52993 = t52992 ^ t52992;
    wire t52994 = t52993 ^ t52993;
    wire t52995 = t52994 ^ t52994;
    wire t52996 = t52995 ^ t52995;
    wire t52997 = t52996 ^ t52996;
    wire t52998 = t52997 ^ t52997;
    wire t52999 = t52998 ^ t52998;
    wire t53000 = t52999 ^ t52999;
    wire t53001 = t53000 ^ t53000;
    wire t53002 = t53001 ^ t53001;
    wire t53003 = t53002 ^ t53002;
    wire t53004 = t53003 ^ t53003;
    wire t53005 = t53004 ^ t53004;
    wire t53006 = t53005 ^ t53005;
    wire t53007 = t53006 ^ t53006;
    wire t53008 = t53007 ^ t53007;
    wire t53009 = t53008 ^ t53008;
    wire t53010 = t53009 ^ t53009;
    wire t53011 = t53010 ^ t53010;
    wire t53012 = t53011 ^ t53011;
    wire t53013 = t53012 ^ t53012;
    wire t53014 = t53013 ^ t53013;
    wire t53015 = t53014 ^ t53014;
    wire t53016 = t53015 ^ t53015;
    wire t53017 = t53016 ^ t53016;
    wire t53018 = t53017 ^ t53017;
    wire t53019 = t53018 ^ t53018;
    wire t53020 = t53019 ^ t53019;
    wire t53021 = t53020 ^ t53020;
    wire t53022 = t53021 ^ t53021;
    wire t53023 = t53022 ^ t53022;
    wire t53024 = t53023 ^ t53023;
    wire t53025 = t53024 ^ t53024;
    wire t53026 = t53025 ^ t53025;
    wire t53027 = t53026 ^ t53026;
    wire t53028 = t53027 ^ t53027;
    wire t53029 = t53028 ^ t53028;
    wire t53030 = t53029 ^ t53029;
    wire t53031 = t53030 ^ t53030;
    wire t53032 = t53031 ^ t53031;
    wire t53033 = t53032 ^ t53032;
    wire t53034 = t53033 ^ t53033;
    wire t53035 = t53034 ^ t53034;
    wire t53036 = t53035 ^ t53035;
    wire t53037 = t53036 ^ t53036;
    wire t53038 = t53037 ^ t53037;
    wire t53039 = t53038 ^ t53038;
    wire t53040 = t53039 ^ t53039;
    wire t53041 = t53040 ^ t53040;
    wire t53042 = t53041 ^ t53041;
    wire t53043 = t53042 ^ t53042;
    wire t53044 = t53043 ^ t53043;
    wire t53045 = t53044 ^ t53044;
    wire t53046 = t53045 ^ t53045;
    wire t53047 = t53046 ^ t53046;
    wire t53048 = t53047 ^ t53047;
    wire t53049 = t53048 ^ t53048;
    wire t53050 = t53049 ^ t53049;
    wire t53051 = t53050 ^ t53050;
    wire t53052 = t53051 ^ t53051;
    wire t53053 = t53052 ^ t53052;
    wire t53054 = t53053 ^ t53053;
    wire t53055 = t53054 ^ t53054;
    wire t53056 = t53055 ^ t53055;
    wire t53057 = t53056 ^ t53056;
    wire t53058 = t53057 ^ t53057;
    wire t53059 = t53058 ^ t53058;
    wire t53060 = t53059 ^ t53059;
    wire t53061 = t53060 ^ t53060;
    wire t53062 = t53061 ^ t53061;
    wire t53063 = t53062 ^ t53062;
    wire t53064 = t53063 ^ t53063;
    wire t53065 = t53064 ^ t53064;
    wire t53066 = t53065 ^ t53065;
    wire t53067 = t53066 ^ t53066;
    wire t53068 = t53067 ^ t53067;
    wire t53069 = t53068 ^ t53068;
    wire t53070 = t53069 ^ t53069;
    wire t53071 = t53070 ^ t53070;
    wire t53072 = t53071 ^ t53071;
    wire t53073 = t53072 ^ t53072;
    wire t53074 = t53073 ^ t53073;
    wire t53075 = t53074 ^ t53074;
    wire t53076 = t53075 ^ t53075;
    wire t53077 = t53076 ^ t53076;
    wire t53078 = t53077 ^ t53077;
    wire t53079 = t53078 ^ t53078;
    wire t53080 = t53079 ^ t53079;
    wire t53081 = t53080 ^ t53080;
    wire t53082 = t53081 ^ t53081;
    wire t53083 = t53082 ^ t53082;
    wire t53084 = t53083 ^ t53083;
    wire t53085 = t53084 ^ t53084;
    wire t53086 = t53085 ^ t53085;
    wire t53087 = t53086 ^ t53086;
    wire t53088 = t53087 ^ t53087;
    wire t53089 = t53088 ^ t53088;
    wire t53090 = t53089 ^ t53089;
    wire t53091 = t53090 ^ t53090;
    wire t53092 = t53091 ^ t53091;
    wire t53093 = t53092 ^ t53092;
    wire t53094 = t53093 ^ t53093;
    wire t53095 = t53094 ^ t53094;
    wire t53096 = t53095 ^ t53095;
    wire t53097 = t53096 ^ t53096;
    wire t53098 = t53097 ^ t53097;
    wire t53099 = t53098 ^ t53098;
    wire t53100 = t53099 ^ t53099;
    wire t53101 = t53100 ^ t53100;
    wire t53102 = t53101 ^ t53101;
    wire t53103 = t53102 ^ t53102;
    wire t53104 = t53103 ^ t53103;
    wire t53105 = t53104 ^ t53104;
    wire t53106 = t53105 ^ t53105;
    wire t53107 = t53106 ^ t53106;
    wire t53108 = t53107 ^ t53107;
    wire t53109 = t53108 ^ t53108;
    wire t53110 = t53109 ^ t53109;
    wire t53111 = t53110 ^ t53110;
    wire t53112 = t53111 ^ t53111;
    wire t53113 = t53112 ^ t53112;
    wire t53114 = t53113 ^ t53113;
    wire t53115 = t53114 ^ t53114;
    wire t53116 = t53115 ^ t53115;
    wire t53117 = t53116 ^ t53116;
    wire t53118 = t53117 ^ t53117;
    wire t53119 = t53118 ^ t53118;
    wire t53120 = t53119 ^ t53119;
    wire t53121 = t53120 ^ t53120;
    wire t53122 = t53121 ^ t53121;
    wire t53123 = t53122 ^ t53122;
    wire t53124 = t53123 ^ t53123;
    wire t53125 = t53124 ^ t53124;
    wire t53126 = t53125 ^ t53125;
    wire t53127 = t53126 ^ t53126;
    wire t53128 = t53127 ^ t53127;
    wire t53129 = t53128 ^ t53128;
    wire t53130 = t53129 ^ t53129;
    wire t53131 = t53130 ^ t53130;
    wire t53132 = t53131 ^ t53131;
    wire t53133 = t53132 ^ t53132;
    wire t53134 = t53133 ^ t53133;
    wire t53135 = t53134 ^ t53134;
    wire t53136 = t53135 ^ t53135;
    wire t53137 = t53136 ^ t53136;
    wire t53138 = t53137 ^ t53137;
    wire t53139 = t53138 ^ t53138;
    wire t53140 = t53139 ^ t53139;
    wire t53141 = t53140 ^ t53140;
    wire t53142 = t53141 ^ t53141;
    wire t53143 = t53142 ^ t53142;
    wire t53144 = t53143 ^ t53143;
    wire t53145 = t53144 ^ t53144;
    wire t53146 = t53145 ^ t53145;
    wire t53147 = t53146 ^ t53146;
    wire t53148 = t53147 ^ t53147;
    wire t53149 = t53148 ^ t53148;
    wire t53150 = t53149 ^ t53149;
    wire t53151 = t53150 ^ t53150;
    wire t53152 = t53151 ^ t53151;
    wire t53153 = t53152 ^ t53152;
    wire t53154 = t53153 ^ t53153;
    wire t53155 = t53154 ^ t53154;
    wire t53156 = t53155 ^ t53155;
    wire t53157 = t53156 ^ t53156;
    wire t53158 = t53157 ^ t53157;
    wire t53159 = t53158 ^ t53158;
    wire t53160 = t53159 ^ t53159;
    wire t53161 = t53160 ^ t53160;
    wire t53162 = t53161 ^ t53161;
    wire t53163 = t53162 ^ t53162;
    wire t53164 = t53163 ^ t53163;
    wire t53165 = t53164 ^ t53164;
    wire t53166 = t53165 ^ t53165;
    wire t53167 = t53166 ^ t53166;
    wire t53168 = t53167 ^ t53167;
    wire t53169 = t53168 ^ t53168;
    wire t53170 = t53169 ^ t53169;
    wire t53171 = t53170 ^ t53170;
    wire t53172 = t53171 ^ t53171;
    wire t53173 = t53172 ^ t53172;
    wire t53174 = t53173 ^ t53173;
    wire t53175 = t53174 ^ t53174;
    wire t53176 = t53175 ^ t53175;
    wire t53177 = t53176 ^ t53176;
    wire t53178 = t53177 ^ t53177;
    wire t53179 = t53178 ^ t53178;
    wire t53180 = t53179 ^ t53179;
    wire t53181 = t53180 ^ t53180;
    wire t53182 = t53181 ^ t53181;
    wire t53183 = t53182 ^ t53182;
    wire t53184 = t53183 ^ t53183;
    wire t53185 = t53184 ^ t53184;
    wire t53186 = t53185 ^ t53185;
    wire t53187 = t53186 ^ t53186;
    wire t53188 = t53187 ^ t53187;
    wire t53189 = t53188 ^ t53188;
    wire t53190 = t53189 ^ t53189;
    wire t53191 = t53190 ^ t53190;
    wire t53192 = t53191 ^ t53191;
    wire t53193 = t53192 ^ t53192;
    wire t53194 = t53193 ^ t53193;
    wire t53195 = t53194 ^ t53194;
    wire t53196 = t53195 ^ t53195;
    wire t53197 = t53196 ^ t53196;
    wire t53198 = t53197 ^ t53197;
    wire t53199 = t53198 ^ t53198;
    wire t53200 = t53199 ^ t53199;
    wire t53201 = t53200 ^ t53200;
    wire t53202 = t53201 ^ t53201;
    wire t53203 = t53202 ^ t53202;
    wire t53204 = t53203 ^ t53203;
    wire t53205 = t53204 ^ t53204;
    wire t53206 = t53205 ^ t53205;
    wire t53207 = t53206 ^ t53206;
    wire t53208 = t53207 ^ t53207;
    wire t53209 = t53208 ^ t53208;
    wire t53210 = t53209 ^ t53209;
    wire t53211 = t53210 ^ t53210;
    wire t53212 = t53211 ^ t53211;
    wire t53213 = t53212 ^ t53212;
    wire t53214 = t53213 ^ t53213;
    wire t53215 = t53214 ^ t53214;
    wire t53216 = t53215 ^ t53215;
    wire t53217 = t53216 ^ t53216;
    wire t53218 = t53217 ^ t53217;
    wire t53219 = t53218 ^ t53218;
    wire t53220 = t53219 ^ t53219;
    wire t53221 = t53220 ^ t53220;
    wire t53222 = t53221 ^ t53221;
    wire t53223 = t53222 ^ t53222;
    wire t53224 = t53223 ^ t53223;
    wire t53225 = t53224 ^ t53224;
    wire t53226 = t53225 ^ t53225;
    wire t53227 = t53226 ^ t53226;
    wire t53228 = t53227 ^ t53227;
    wire t53229 = t53228 ^ t53228;
    wire t53230 = t53229 ^ t53229;
    wire t53231 = t53230 ^ t53230;
    wire t53232 = t53231 ^ t53231;
    wire t53233 = t53232 ^ t53232;
    wire t53234 = t53233 ^ t53233;
    wire t53235 = t53234 ^ t53234;
    wire t53236 = t53235 ^ t53235;
    wire t53237 = t53236 ^ t53236;
    wire t53238 = t53237 ^ t53237;
    wire t53239 = t53238 ^ t53238;
    wire t53240 = t53239 ^ t53239;
    wire t53241 = t53240 ^ t53240;
    wire t53242 = t53241 ^ t53241;
    wire t53243 = t53242 ^ t53242;
    wire t53244 = t53243 ^ t53243;
    wire t53245 = t53244 ^ t53244;
    wire t53246 = t53245 ^ t53245;
    wire t53247 = t53246 ^ t53246;
    wire t53248 = t53247 ^ t53247;
    wire t53249 = t53248 ^ t53248;
    wire t53250 = t53249 ^ t53249;
    wire t53251 = t53250 ^ t53250;
    wire t53252 = t53251 ^ t53251;
    wire t53253 = t53252 ^ t53252;
    wire t53254 = t53253 ^ t53253;
    wire t53255 = t53254 ^ t53254;
    wire t53256 = t53255 ^ t53255;
    wire t53257 = t53256 ^ t53256;
    wire t53258 = t53257 ^ t53257;
    wire t53259 = t53258 ^ t53258;
    wire t53260 = t53259 ^ t53259;
    wire t53261 = t53260 ^ t53260;
    wire t53262 = t53261 ^ t53261;
    wire t53263 = t53262 ^ t53262;
    wire t53264 = t53263 ^ t53263;
    wire t53265 = t53264 ^ t53264;
    wire t53266 = t53265 ^ t53265;
    wire t53267 = t53266 ^ t53266;
    wire t53268 = t53267 ^ t53267;
    wire t53269 = t53268 ^ t53268;
    wire t53270 = t53269 ^ t53269;
    wire t53271 = t53270 ^ t53270;
    wire t53272 = t53271 ^ t53271;
    wire t53273 = t53272 ^ t53272;
    wire t53274 = t53273 ^ t53273;
    wire t53275 = t53274 ^ t53274;
    wire t53276 = t53275 ^ t53275;
    wire t53277 = t53276 ^ t53276;
    wire t53278 = t53277 ^ t53277;
    wire t53279 = t53278 ^ t53278;
    wire t53280 = t53279 ^ t53279;
    wire t53281 = t53280 ^ t53280;
    wire t53282 = t53281 ^ t53281;
    wire t53283 = t53282 ^ t53282;
    wire t53284 = t53283 ^ t53283;
    wire t53285 = t53284 ^ t53284;
    wire t53286 = t53285 ^ t53285;
    wire t53287 = t53286 ^ t53286;
    wire t53288 = t53287 ^ t53287;
    wire t53289 = t53288 ^ t53288;
    wire t53290 = t53289 ^ t53289;
    wire t53291 = t53290 ^ t53290;
    wire t53292 = t53291 ^ t53291;
    wire t53293 = t53292 ^ t53292;
    wire t53294 = t53293 ^ t53293;
    wire t53295 = t53294 ^ t53294;
    wire t53296 = t53295 ^ t53295;
    wire t53297 = t53296 ^ t53296;
    wire t53298 = t53297 ^ t53297;
    wire t53299 = t53298 ^ t53298;
    wire t53300 = t53299 ^ t53299;
    wire t53301 = t53300 ^ t53300;
    wire t53302 = t53301 ^ t53301;
    wire t53303 = t53302 ^ t53302;
    wire t53304 = t53303 ^ t53303;
    wire t53305 = t53304 ^ t53304;
    wire t53306 = t53305 ^ t53305;
    wire t53307 = t53306 ^ t53306;
    wire t53308 = t53307 ^ t53307;
    wire t53309 = t53308 ^ t53308;
    wire t53310 = t53309 ^ t53309;
    wire t53311 = t53310 ^ t53310;
    wire t53312 = t53311 ^ t53311;
    wire t53313 = t53312 ^ t53312;
    wire t53314 = t53313 ^ t53313;
    wire t53315 = t53314 ^ t53314;
    wire t53316 = t53315 ^ t53315;
    wire t53317 = t53316 ^ t53316;
    wire t53318 = t53317 ^ t53317;
    wire t53319 = t53318 ^ t53318;
    wire t53320 = t53319 ^ t53319;
    wire t53321 = t53320 ^ t53320;
    wire t53322 = t53321 ^ t53321;
    wire t53323 = t53322 ^ t53322;
    wire t53324 = t53323 ^ t53323;
    wire t53325 = t53324 ^ t53324;
    wire t53326 = t53325 ^ t53325;
    wire t53327 = t53326 ^ t53326;
    wire t53328 = t53327 ^ t53327;
    wire t53329 = t53328 ^ t53328;
    wire t53330 = t53329 ^ t53329;
    wire t53331 = t53330 ^ t53330;
    wire t53332 = t53331 ^ t53331;
    wire t53333 = t53332 ^ t53332;
    wire t53334 = t53333 ^ t53333;
    wire t53335 = t53334 ^ t53334;
    wire t53336 = t53335 ^ t53335;
    wire t53337 = t53336 ^ t53336;
    wire t53338 = t53337 ^ t53337;
    wire t53339 = t53338 ^ t53338;
    wire t53340 = t53339 ^ t53339;
    wire t53341 = t53340 ^ t53340;
    wire t53342 = t53341 ^ t53341;
    wire t53343 = t53342 ^ t53342;
    wire t53344 = t53343 ^ t53343;
    wire t53345 = t53344 ^ t53344;
    wire t53346 = t53345 ^ t53345;
    wire t53347 = t53346 ^ t53346;
    wire t53348 = t53347 ^ t53347;
    wire t53349 = t53348 ^ t53348;
    wire t53350 = t53349 ^ t53349;
    wire t53351 = t53350 ^ t53350;
    wire t53352 = t53351 ^ t53351;
    wire t53353 = t53352 ^ t53352;
    wire t53354 = t53353 ^ t53353;
    wire t53355 = t53354 ^ t53354;
    wire t53356 = t53355 ^ t53355;
    wire t53357 = t53356 ^ t53356;
    wire t53358 = t53357 ^ t53357;
    wire t53359 = t53358 ^ t53358;
    wire t53360 = t53359 ^ t53359;
    wire t53361 = t53360 ^ t53360;
    wire t53362 = t53361 ^ t53361;
    wire t53363 = t53362 ^ t53362;
    wire t53364 = t53363 ^ t53363;
    wire t53365 = t53364 ^ t53364;
    wire t53366 = t53365 ^ t53365;
    wire t53367 = t53366 ^ t53366;
    wire t53368 = t53367 ^ t53367;
    wire t53369 = t53368 ^ t53368;
    wire t53370 = t53369 ^ t53369;
    wire t53371 = t53370 ^ t53370;
    wire t53372 = t53371 ^ t53371;
    wire t53373 = t53372 ^ t53372;
    wire t53374 = t53373 ^ t53373;
    wire t53375 = t53374 ^ t53374;
    wire t53376 = t53375 ^ t53375;
    wire t53377 = t53376 ^ t53376;
    wire t53378 = t53377 ^ t53377;
    wire t53379 = t53378 ^ t53378;
    wire t53380 = t53379 ^ t53379;
    wire t53381 = t53380 ^ t53380;
    wire t53382 = t53381 ^ t53381;
    wire t53383 = t53382 ^ t53382;
    wire t53384 = t53383 ^ t53383;
    wire t53385 = t53384 ^ t53384;
    wire t53386 = t53385 ^ t53385;
    wire t53387 = t53386 ^ t53386;
    wire t53388 = t53387 ^ t53387;
    wire t53389 = t53388 ^ t53388;
    wire t53390 = t53389 ^ t53389;
    wire t53391 = t53390 ^ t53390;
    wire t53392 = t53391 ^ t53391;
    wire t53393 = t53392 ^ t53392;
    wire t53394 = t53393 ^ t53393;
    wire t53395 = t53394 ^ t53394;
    wire t53396 = t53395 ^ t53395;
    wire t53397 = t53396 ^ t53396;
    wire t53398 = t53397 ^ t53397;
    wire t53399 = t53398 ^ t53398;
    wire t53400 = t53399 ^ t53399;
    wire t53401 = t53400 ^ t53400;
    wire t53402 = t53401 ^ t53401;
    wire t53403 = t53402 ^ t53402;
    wire t53404 = t53403 ^ t53403;
    wire t53405 = t53404 ^ t53404;
    wire t53406 = t53405 ^ t53405;
    wire t53407 = t53406 ^ t53406;
    wire t53408 = t53407 ^ t53407;
    wire t53409 = t53408 ^ t53408;
    wire t53410 = t53409 ^ t53409;
    wire t53411 = t53410 ^ t53410;
    wire t53412 = t53411 ^ t53411;
    wire t53413 = t53412 ^ t53412;
    wire t53414 = t53413 ^ t53413;
    wire t53415 = t53414 ^ t53414;
    wire t53416 = t53415 ^ t53415;
    wire t53417 = t53416 ^ t53416;
    wire t53418 = t53417 ^ t53417;
    wire t53419 = t53418 ^ t53418;
    wire t53420 = t53419 ^ t53419;
    wire t53421 = t53420 ^ t53420;
    wire t53422 = t53421 ^ t53421;
    wire t53423 = t53422 ^ t53422;
    wire t53424 = t53423 ^ t53423;
    wire t53425 = t53424 ^ t53424;
    wire t53426 = t53425 ^ t53425;
    wire t53427 = t53426 ^ t53426;
    wire t53428 = t53427 ^ t53427;
    wire t53429 = t53428 ^ t53428;
    wire t53430 = t53429 ^ t53429;
    wire t53431 = t53430 ^ t53430;
    wire t53432 = t53431 ^ t53431;
    wire t53433 = t53432 ^ t53432;
    wire t53434 = t53433 ^ t53433;
    wire t53435 = t53434 ^ t53434;
    wire t53436 = t53435 ^ t53435;
    wire t53437 = t53436 ^ t53436;
    wire t53438 = t53437 ^ t53437;
    wire t53439 = t53438 ^ t53438;
    wire t53440 = t53439 ^ t53439;
    wire t53441 = t53440 ^ t53440;
    wire t53442 = t53441 ^ t53441;
    wire t53443 = t53442 ^ t53442;
    wire t53444 = t53443 ^ t53443;
    wire t53445 = t53444 ^ t53444;
    wire t53446 = t53445 ^ t53445;
    wire t53447 = t53446 ^ t53446;
    wire t53448 = t53447 ^ t53447;
    wire t53449 = t53448 ^ t53448;
    wire t53450 = t53449 ^ t53449;
    wire t53451 = t53450 ^ t53450;
    wire t53452 = t53451 ^ t53451;
    wire t53453 = t53452 ^ t53452;
    wire t53454 = t53453 ^ t53453;
    wire t53455 = t53454 ^ t53454;
    wire t53456 = t53455 ^ t53455;
    wire t53457 = t53456 ^ t53456;
    wire t53458 = t53457 ^ t53457;
    wire t53459 = t53458 ^ t53458;
    wire t53460 = t53459 ^ t53459;
    wire t53461 = t53460 ^ t53460;
    wire t53462 = t53461 ^ t53461;
    wire t53463 = t53462 ^ t53462;
    wire t53464 = t53463 ^ t53463;
    wire t53465 = t53464 ^ t53464;
    wire t53466 = t53465 ^ t53465;
    wire t53467 = t53466 ^ t53466;
    wire t53468 = t53467 ^ t53467;
    wire t53469 = t53468 ^ t53468;
    wire t53470 = t53469 ^ t53469;
    wire t53471 = t53470 ^ t53470;
    wire t53472 = t53471 ^ t53471;
    wire t53473 = t53472 ^ t53472;
    wire t53474 = t53473 ^ t53473;
    wire t53475 = t53474 ^ t53474;
    wire t53476 = t53475 ^ t53475;
    wire t53477 = t53476 ^ t53476;
    wire t53478 = t53477 ^ t53477;
    wire t53479 = t53478 ^ t53478;
    wire t53480 = t53479 ^ t53479;
    wire t53481 = t53480 ^ t53480;
    wire t53482 = t53481 ^ t53481;
    wire t53483 = t53482 ^ t53482;
    wire t53484 = t53483 ^ t53483;
    wire t53485 = t53484 ^ t53484;
    wire t53486 = t53485 ^ t53485;
    wire t53487 = t53486 ^ t53486;
    wire t53488 = t53487 ^ t53487;
    wire t53489 = t53488 ^ t53488;
    wire t53490 = t53489 ^ t53489;
    wire t53491 = t53490 ^ t53490;
    wire t53492 = t53491 ^ t53491;
    wire t53493 = t53492 ^ t53492;
    wire t53494 = t53493 ^ t53493;
    wire t53495 = t53494 ^ t53494;
    wire t53496 = t53495 ^ t53495;
    wire t53497 = t53496 ^ t53496;
    wire t53498 = t53497 ^ t53497;
    wire t53499 = t53498 ^ t53498;
    wire t53500 = t53499 ^ t53499;
    wire t53501 = t53500 ^ t53500;
    wire t53502 = t53501 ^ t53501;
    wire t53503 = t53502 ^ t53502;
    wire t53504 = t53503 ^ t53503;
    wire t53505 = t53504 ^ t53504;
    wire t53506 = t53505 ^ t53505;
    wire t53507 = t53506 ^ t53506;
    wire t53508 = t53507 ^ t53507;
    wire t53509 = t53508 ^ t53508;
    wire t53510 = t53509 ^ t53509;
    wire t53511 = t53510 ^ t53510;
    wire t53512 = t53511 ^ t53511;
    wire t53513 = t53512 ^ t53512;
    wire t53514 = t53513 ^ t53513;
    wire t53515 = t53514 ^ t53514;
    wire t53516 = t53515 ^ t53515;
    wire t53517 = t53516 ^ t53516;
    wire t53518 = t53517 ^ t53517;
    wire t53519 = t53518 ^ t53518;
    wire t53520 = t53519 ^ t53519;
    wire t53521 = t53520 ^ t53520;
    wire t53522 = t53521 ^ t53521;
    wire t53523 = t53522 ^ t53522;
    wire t53524 = t53523 ^ t53523;
    wire t53525 = t53524 ^ t53524;
    wire t53526 = t53525 ^ t53525;
    wire t53527 = t53526 ^ t53526;
    wire t53528 = t53527 ^ t53527;
    wire t53529 = t53528 ^ t53528;
    wire t53530 = t53529 ^ t53529;
    wire t53531 = t53530 ^ t53530;
    wire t53532 = t53531 ^ t53531;
    wire t53533 = t53532 ^ t53532;
    wire t53534 = t53533 ^ t53533;
    wire t53535 = t53534 ^ t53534;
    wire t53536 = t53535 ^ t53535;
    wire t53537 = t53536 ^ t53536;
    wire t53538 = t53537 ^ t53537;
    wire t53539 = t53538 ^ t53538;
    wire t53540 = t53539 ^ t53539;
    wire t53541 = t53540 ^ t53540;
    wire t53542 = t53541 ^ t53541;
    wire t53543 = t53542 ^ t53542;
    wire t53544 = t53543 ^ t53543;
    wire t53545 = t53544 ^ t53544;
    wire t53546 = t53545 ^ t53545;
    wire t53547 = t53546 ^ t53546;
    wire t53548 = t53547 ^ t53547;
    wire t53549 = t53548 ^ t53548;
    wire t53550 = t53549 ^ t53549;
    wire t53551 = t53550 ^ t53550;
    wire t53552 = t53551 ^ t53551;
    wire t53553 = t53552 ^ t53552;
    wire t53554 = t53553 ^ t53553;
    wire t53555 = t53554 ^ t53554;
    wire t53556 = t53555 ^ t53555;
    wire t53557 = t53556 ^ t53556;
    wire t53558 = t53557 ^ t53557;
    wire t53559 = t53558 ^ t53558;
    wire t53560 = t53559 ^ t53559;
    wire t53561 = t53560 ^ t53560;
    wire t53562 = t53561 ^ t53561;
    wire t53563 = t53562 ^ t53562;
    wire t53564 = t53563 ^ t53563;
    wire t53565 = t53564 ^ t53564;
    wire t53566 = t53565 ^ t53565;
    wire t53567 = t53566 ^ t53566;
    wire t53568 = t53567 ^ t53567;
    wire t53569 = t53568 ^ t53568;
    wire t53570 = t53569 ^ t53569;
    wire t53571 = t53570 ^ t53570;
    wire t53572 = t53571 ^ t53571;
    wire t53573 = t53572 ^ t53572;
    wire t53574 = t53573 ^ t53573;
    wire t53575 = t53574 ^ t53574;
    wire t53576 = t53575 ^ t53575;
    wire t53577 = t53576 ^ t53576;
    wire t53578 = t53577 ^ t53577;
    wire t53579 = t53578 ^ t53578;
    wire t53580 = t53579 ^ t53579;
    wire t53581 = t53580 ^ t53580;
    wire t53582 = t53581 ^ t53581;
    wire t53583 = t53582 ^ t53582;
    wire t53584 = t53583 ^ t53583;
    wire t53585 = t53584 ^ t53584;
    wire t53586 = t53585 ^ t53585;
    wire t53587 = t53586 ^ t53586;
    wire t53588 = t53587 ^ t53587;
    wire t53589 = t53588 ^ t53588;
    wire t53590 = t53589 ^ t53589;
    wire t53591 = t53590 ^ t53590;
    wire t53592 = t53591 ^ t53591;
    wire t53593 = t53592 ^ t53592;
    wire t53594 = t53593 ^ t53593;
    wire t53595 = t53594 ^ t53594;
    wire t53596 = t53595 ^ t53595;
    wire t53597 = t53596 ^ t53596;
    wire t53598 = t53597 ^ t53597;
    wire t53599 = t53598 ^ t53598;
    wire t53600 = t53599 ^ t53599;
    wire t53601 = t53600 ^ t53600;
    wire t53602 = t53601 ^ t53601;
    wire t53603 = t53602 ^ t53602;
    wire t53604 = t53603 ^ t53603;
    wire t53605 = t53604 ^ t53604;
    wire t53606 = t53605 ^ t53605;
    wire t53607 = t53606 ^ t53606;
    wire t53608 = t53607 ^ t53607;
    wire t53609 = t53608 ^ t53608;
    wire t53610 = t53609 ^ t53609;
    wire t53611 = t53610 ^ t53610;
    wire t53612 = t53611 ^ t53611;
    wire t53613 = t53612 ^ t53612;
    wire t53614 = t53613 ^ t53613;
    wire t53615 = t53614 ^ t53614;
    wire t53616 = t53615 ^ t53615;
    wire t53617 = t53616 ^ t53616;
    wire t53618 = t53617 ^ t53617;
    wire t53619 = t53618 ^ t53618;
    wire t53620 = t53619 ^ t53619;
    wire t53621 = t53620 ^ t53620;
    wire t53622 = t53621 ^ t53621;
    wire t53623 = t53622 ^ t53622;
    wire t53624 = t53623 ^ t53623;
    wire t53625 = t53624 ^ t53624;
    wire t53626 = t53625 ^ t53625;
    wire t53627 = t53626 ^ t53626;
    wire t53628 = t53627 ^ t53627;
    wire t53629 = t53628 ^ t53628;
    wire t53630 = t53629 ^ t53629;
    wire t53631 = t53630 ^ t53630;
    wire t53632 = t53631 ^ t53631;
    wire t53633 = t53632 ^ t53632;
    wire t53634 = t53633 ^ t53633;
    wire t53635 = t53634 ^ t53634;
    wire t53636 = t53635 ^ t53635;
    wire t53637 = t53636 ^ t53636;
    wire t53638 = t53637 ^ t53637;
    wire t53639 = t53638 ^ t53638;
    wire t53640 = t53639 ^ t53639;
    wire t53641 = t53640 ^ t53640;
    wire t53642 = t53641 ^ t53641;
    wire t53643 = t53642 ^ t53642;
    wire t53644 = t53643 ^ t53643;
    wire t53645 = t53644 ^ t53644;
    wire t53646 = t53645 ^ t53645;
    wire t53647 = t53646 ^ t53646;
    wire t53648 = t53647 ^ t53647;
    wire t53649 = t53648 ^ t53648;
    wire t53650 = t53649 ^ t53649;
    wire t53651 = t53650 ^ t53650;
    wire t53652 = t53651 ^ t53651;
    wire t53653 = t53652 ^ t53652;
    wire t53654 = t53653 ^ t53653;
    wire t53655 = t53654 ^ t53654;
    wire t53656 = t53655 ^ t53655;
    wire t53657 = t53656 ^ t53656;
    wire t53658 = t53657 ^ t53657;
    wire t53659 = t53658 ^ t53658;
    wire t53660 = t53659 ^ t53659;
    wire t53661 = t53660 ^ t53660;
    wire t53662 = t53661 ^ t53661;
    wire t53663 = t53662 ^ t53662;
    wire t53664 = t53663 ^ t53663;
    wire t53665 = t53664 ^ t53664;
    wire t53666 = t53665 ^ t53665;
    wire t53667 = t53666 ^ t53666;
    wire t53668 = t53667 ^ t53667;
    wire t53669 = t53668 ^ t53668;
    wire t53670 = t53669 ^ t53669;
    wire t53671 = t53670 ^ t53670;
    wire t53672 = t53671 ^ t53671;
    wire t53673 = t53672 ^ t53672;
    wire t53674 = t53673 ^ t53673;
    wire t53675 = t53674 ^ t53674;
    wire t53676 = t53675 ^ t53675;
    wire t53677 = t53676 ^ t53676;
    wire t53678 = t53677 ^ t53677;
    wire t53679 = t53678 ^ t53678;
    wire t53680 = t53679 ^ t53679;
    wire t53681 = t53680 ^ t53680;
    wire t53682 = t53681 ^ t53681;
    wire t53683 = t53682 ^ t53682;
    wire t53684 = t53683 ^ t53683;
    wire t53685 = t53684 ^ t53684;
    wire t53686 = t53685 ^ t53685;
    wire t53687 = t53686 ^ t53686;
    wire t53688 = t53687 ^ t53687;
    wire t53689 = t53688 ^ t53688;
    wire t53690 = t53689 ^ t53689;
    wire t53691 = t53690 ^ t53690;
    wire t53692 = t53691 ^ t53691;
    wire t53693 = t53692 ^ t53692;
    wire t53694 = t53693 ^ t53693;
    wire t53695 = t53694 ^ t53694;
    wire t53696 = t53695 ^ t53695;
    wire t53697 = t53696 ^ t53696;
    wire t53698 = t53697 ^ t53697;
    wire t53699 = t53698 ^ t53698;
    wire t53700 = t53699 ^ t53699;
    wire t53701 = t53700 ^ t53700;
    wire t53702 = t53701 ^ t53701;
    wire t53703 = t53702 ^ t53702;
    wire t53704 = t53703 ^ t53703;
    wire t53705 = t53704 ^ t53704;
    wire t53706 = t53705 ^ t53705;
    wire t53707 = t53706 ^ t53706;
    wire t53708 = t53707 ^ t53707;
    wire t53709 = t53708 ^ t53708;
    wire t53710 = t53709 ^ t53709;
    wire t53711 = t53710 ^ t53710;
    wire t53712 = t53711 ^ t53711;
    wire t53713 = t53712 ^ t53712;
    wire t53714 = t53713 ^ t53713;
    wire t53715 = t53714 ^ t53714;
    wire t53716 = t53715 ^ t53715;
    wire t53717 = t53716 ^ t53716;
    wire t53718 = t53717 ^ t53717;
    wire t53719 = t53718 ^ t53718;
    wire t53720 = t53719 ^ t53719;
    wire t53721 = t53720 ^ t53720;
    wire t53722 = t53721 ^ t53721;
    wire t53723 = t53722 ^ t53722;
    wire t53724 = t53723 ^ t53723;
    wire t53725 = t53724 ^ t53724;
    wire t53726 = t53725 ^ t53725;
    wire t53727 = t53726 ^ t53726;
    wire t53728 = t53727 ^ t53727;
    wire t53729 = t53728 ^ t53728;
    wire t53730 = t53729 ^ t53729;
    wire t53731 = t53730 ^ t53730;
    wire t53732 = t53731 ^ t53731;
    wire t53733 = t53732 ^ t53732;
    wire t53734 = t53733 ^ t53733;
    wire t53735 = t53734 ^ t53734;
    wire t53736 = t53735 ^ t53735;
    wire t53737 = t53736 ^ t53736;
    wire t53738 = t53737 ^ t53737;
    wire t53739 = t53738 ^ t53738;
    wire t53740 = t53739 ^ t53739;
    wire t53741 = t53740 ^ t53740;
    wire t53742 = t53741 ^ t53741;
    wire t53743 = t53742 ^ t53742;
    wire t53744 = t53743 ^ t53743;
    wire t53745 = t53744 ^ t53744;
    wire t53746 = t53745 ^ t53745;
    wire t53747 = t53746 ^ t53746;
    wire t53748 = t53747 ^ t53747;
    wire t53749 = t53748 ^ t53748;
    wire t53750 = t53749 ^ t53749;
    wire t53751 = t53750 ^ t53750;
    wire t53752 = t53751 ^ t53751;
    wire t53753 = t53752 ^ t53752;
    wire t53754 = t53753 ^ t53753;
    wire t53755 = t53754 ^ t53754;
    wire t53756 = t53755 ^ t53755;
    wire t53757 = t53756 ^ t53756;
    wire t53758 = t53757 ^ t53757;
    wire t53759 = t53758 ^ t53758;
    wire t53760 = t53759 ^ t53759;
    wire t53761 = t53760 ^ t53760;
    wire t53762 = t53761 ^ t53761;
    wire t53763 = t53762 ^ t53762;
    wire t53764 = t53763 ^ t53763;
    wire t53765 = t53764 ^ t53764;
    wire t53766 = t53765 ^ t53765;
    wire t53767 = t53766 ^ t53766;
    wire t53768 = t53767 ^ t53767;
    wire t53769 = t53768 ^ t53768;
    wire t53770 = t53769 ^ t53769;
    wire t53771 = t53770 ^ t53770;
    wire t53772 = t53771 ^ t53771;
    wire t53773 = t53772 ^ t53772;
    wire t53774 = t53773 ^ t53773;
    wire t53775 = t53774 ^ t53774;
    wire t53776 = t53775 ^ t53775;
    wire t53777 = t53776 ^ t53776;
    wire t53778 = t53777 ^ t53777;
    wire t53779 = t53778 ^ t53778;
    wire t53780 = t53779 ^ t53779;
    wire t53781 = t53780 ^ t53780;
    wire t53782 = t53781 ^ t53781;
    wire t53783 = t53782 ^ t53782;
    wire t53784 = t53783 ^ t53783;
    wire t53785 = t53784 ^ t53784;
    wire t53786 = t53785 ^ t53785;
    wire t53787 = t53786 ^ t53786;
    wire t53788 = t53787 ^ t53787;
    wire t53789 = t53788 ^ t53788;
    wire t53790 = t53789 ^ t53789;
    wire t53791 = t53790 ^ t53790;
    wire t53792 = t53791 ^ t53791;
    wire t53793 = t53792 ^ t53792;
    wire t53794 = t53793 ^ t53793;
    wire t53795 = t53794 ^ t53794;
    wire t53796 = t53795 ^ t53795;
    wire t53797 = t53796 ^ t53796;
    wire t53798 = t53797 ^ t53797;
    wire t53799 = t53798 ^ t53798;
    wire t53800 = t53799 ^ t53799;
    wire t53801 = t53800 ^ t53800;
    wire t53802 = t53801 ^ t53801;
    wire t53803 = t53802 ^ t53802;
    wire t53804 = t53803 ^ t53803;
    wire t53805 = t53804 ^ t53804;
    wire t53806 = t53805 ^ t53805;
    wire t53807 = t53806 ^ t53806;
    wire t53808 = t53807 ^ t53807;
    wire t53809 = t53808 ^ t53808;
    wire t53810 = t53809 ^ t53809;
    wire t53811 = t53810 ^ t53810;
    wire t53812 = t53811 ^ t53811;
    wire t53813 = t53812 ^ t53812;
    wire t53814 = t53813 ^ t53813;
    wire t53815 = t53814 ^ t53814;
    wire t53816 = t53815 ^ t53815;
    wire t53817 = t53816 ^ t53816;
    wire t53818 = t53817 ^ t53817;
    wire t53819 = t53818 ^ t53818;
    wire t53820 = t53819 ^ t53819;
    wire t53821 = t53820 ^ t53820;
    wire t53822 = t53821 ^ t53821;
    wire t53823 = t53822 ^ t53822;
    wire t53824 = t53823 ^ t53823;
    wire t53825 = t53824 ^ t53824;
    wire t53826 = t53825 ^ t53825;
    wire t53827 = t53826 ^ t53826;
    wire t53828 = t53827 ^ t53827;
    wire t53829 = t53828 ^ t53828;
    wire t53830 = t53829 ^ t53829;
    wire t53831 = t53830 ^ t53830;
    wire t53832 = t53831 ^ t53831;
    wire t53833 = t53832 ^ t53832;
    wire t53834 = t53833 ^ t53833;
    wire t53835 = t53834 ^ t53834;
    wire t53836 = t53835 ^ t53835;
    wire t53837 = t53836 ^ t53836;
    wire t53838 = t53837 ^ t53837;
    wire t53839 = t53838 ^ t53838;
    wire t53840 = t53839 ^ t53839;
    wire t53841 = t53840 ^ t53840;
    wire t53842 = t53841 ^ t53841;
    wire t53843 = t53842 ^ t53842;
    wire t53844 = t53843 ^ t53843;
    wire t53845 = t53844 ^ t53844;
    wire t53846 = t53845 ^ t53845;
    wire t53847 = t53846 ^ t53846;
    wire t53848 = t53847 ^ t53847;
    wire t53849 = t53848 ^ t53848;
    wire t53850 = t53849 ^ t53849;
    wire t53851 = t53850 ^ t53850;
    wire t53852 = t53851 ^ t53851;
    wire t53853 = t53852 ^ t53852;
    wire t53854 = t53853 ^ t53853;
    wire t53855 = t53854 ^ t53854;
    wire t53856 = t53855 ^ t53855;
    wire t53857 = t53856 ^ t53856;
    wire t53858 = t53857 ^ t53857;
    wire t53859 = t53858 ^ t53858;
    wire t53860 = t53859 ^ t53859;
    wire t53861 = t53860 ^ t53860;
    wire t53862 = t53861 ^ t53861;
    wire t53863 = t53862 ^ t53862;
    wire t53864 = t53863 ^ t53863;
    wire t53865 = t53864 ^ t53864;
    wire t53866 = t53865 ^ t53865;
    wire t53867 = t53866 ^ t53866;
    wire t53868 = t53867 ^ t53867;
    wire t53869 = t53868 ^ t53868;
    wire t53870 = t53869 ^ t53869;
    wire t53871 = t53870 ^ t53870;
    wire t53872 = t53871 ^ t53871;
    wire t53873 = t53872 ^ t53872;
    wire t53874 = t53873 ^ t53873;
    wire t53875 = t53874 ^ t53874;
    wire t53876 = t53875 ^ t53875;
    wire t53877 = t53876 ^ t53876;
    wire t53878 = t53877 ^ t53877;
    wire t53879 = t53878 ^ t53878;
    wire t53880 = t53879 ^ t53879;
    wire t53881 = t53880 ^ t53880;
    wire t53882 = t53881 ^ t53881;
    wire t53883 = t53882 ^ t53882;
    wire t53884 = t53883 ^ t53883;
    wire t53885 = t53884 ^ t53884;
    wire t53886 = t53885 ^ t53885;
    wire t53887 = t53886 ^ t53886;
    wire t53888 = t53887 ^ t53887;
    wire t53889 = t53888 ^ t53888;
    wire t53890 = t53889 ^ t53889;
    wire t53891 = t53890 ^ t53890;
    wire t53892 = t53891 ^ t53891;
    wire t53893 = t53892 ^ t53892;
    wire t53894 = t53893 ^ t53893;
    wire t53895 = t53894 ^ t53894;
    wire t53896 = t53895 ^ t53895;
    wire t53897 = t53896 ^ t53896;
    wire t53898 = t53897 ^ t53897;
    wire t53899 = t53898 ^ t53898;
    wire t53900 = t53899 ^ t53899;
    wire t53901 = t53900 ^ t53900;
    wire t53902 = t53901 ^ t53901;
    wire t53903 = t53902 ^ t53902;
    wire t53904 = t53903 ^ t53903;
    wire t53905 = t53904 ^ t53904;
    wire t53906 = t53905 ^ t53905;
    wire t53907 = t53906 ^ t53906;
    wire t53908 = t53907 ^ t53907;
    wire t53909 = t53908 ^ t53908;
    wire t53910 = t53909 ^ t53909;
    wire t53911 = t53910 ^ t53910;
    wire t53912 = t53911 ^ t53911;
    wire t53913 = t53912 ^ t53912;
    wire t53914 = t53913 ^ t53913;
    wire t53915 = t53914 ^ t53914;
    wire t53916 = t53915 ^ t53915;
    wire t53917 = t53916 ^ t53916;
    wire t53918 = t53917 ^ t53917;
    wire t53919 = t53918 ^ t53918;
    wire t53920 = t53919 ^ t53919;
    wire t53921 = t53920 ^ t53920;
    wire t53922 = t53921 ^ t53921;
    wire t53923 = t53922 ^ t53922;
    wire t53924 = t53923 ^ t53923;
    wire t53925 = t53924 ^ t53924;
    wire t53926 = t53925 ^ t53925;
    wire t53927 = t53926 ^ t53926;
    wire t53928 = t53927 ^ t53927;
    wire t53929 = t53928 ^ t53928;
    wire t53930 = t53929 ^ t53929;
    wire t53931 = t53930 ^ t53930;
    wire t53932 = t53931 ^ t53931;
    wire t53933 = t53932 ^ t53932;
    wire t53934 = t53933 ^ t53933;
    wire t53935 = t53934 ^ t53934;
    wire t53936 = t53935 ^ t53935;
    wire t53937 = t53936 ^ t53936;
    wire t53938 = t53937 ^ t53937;
    wire t53939 = t53938 ^ t53938;
    wire t53940 = t53939 ^ t53939;
    wire t53941 = t53940 ^ t53940;
    wire t53942 = t53941 ^ t53941;
    wire t53943 = t53942 ^ t53942;
    wire t53944 = t53943 ^ t53943;
    wire t53945 = t53944 ^ t53944;
    wire t53946 = t53945 ^ t53945;
    wire t53947 = t53946 ^ t53946;
    wire t53948 = t53947 ^ t53947;
    wire t53949 = t53948 ^ t53948;
    wire t53950 = t53949 ^ t53949;
    wire t53951 = t53950 ^ t53950;
    wire t53952 = t53951 ^ t53951;
    wire t53953 = t53952 ^ t53952;
    wire t53954 = t53953 ^ t53953;
    wire t53955 = t53954 ^ t53954;
    wire t53956 = t53955 ^ t53955;
    wire t53957 = t53956 ^ t53956;
    wire t53958 = t53957 ^ t53957;
    wire t53959 = t53958 ^ t53958;
    wire t53960 = t53959 ^ t53959;
    wire t53961 = t53960 ^ t53960;
    wire t53962 = t53961 ^ t53961;
    wire t53963 = t53962 ^ t53962;
    wire t53964 = t53963 ^ t53963;
    wire t53965 = t53964 ^ t53964;
    wire t53966 = t53965 ^ t53965;
    wire t53967 = t53966 ^ t53966;
    wire t53968 = t53967 ^ t53967;
    wire t53969 = t53968 ^ t53968;
    wire t53970 = t53969 ^ t53969;
    wire t53971 = t53970 ^ t53970;
    wire t53972 = t53971 ^ t53971;
    wire t53973 = t53972 ^ t53972;
    wire t53974 = t53973 ^ t53973;
    wire t53975 = t53974 ^ t53974;
    wire t53976 = t53975 ^ t53975;
    wire t53977 = t53976 ^ t53976;
    wire t53978 = t53977 ^ t53977;
    wire t53979 = t53978 ^ t53978;
    wire t53980 = t53979 ^ t53979;
    wire t53981 = t53980 ^ t53980;
    wire t53982 = t53981 ^ t53981;
    wire t53983 = t53982 ^ t53982;
    wire t53984 = t53983 ^ t53983;
    wire t53985 = t53984 ^ t53984;
    wire t53986 = t53985 ^ t53985;
    wire t53987 = t53986 ^ t53986;
    wire t53988 = t53987 ^ t53987;
    wire t53989 = t53988 ^ t53988;
    wire t53990 = t53989 ^ t53989;
    wire t53991 = t53990 ^ t53990;
    wire t53992 = t53991 ^ t53991;
    wire t53993 = t53992 ^ t53992;
    wire t53994 = t53993 ^ t53993;
    wire t53995 = t53994 ^ t53994;
    wire t53996 = t53995 ^ t53995;
    wire t53997 = t53996 ^ t53996;
    wire t53998 = t53997 ^ t53997;
    wire t53999 = t53998 ^ t53998;
    wire t54000 = t53999 ^ t53999;
    wire t54001 = t54000 ^ t54000;
    wire t54002 = t54001 ^ t54001;
    wire t54003 = t54002 ^ t54002;
    wire t54004 = t54003 ^ t54003;
    wire t54005 = t54004 ^ t54004;
    wire t54006 = t54005 ^ t54005;
    wire t54007 = t54006 ^ t54006;
    wire t54008 = t54007 ^ t54007;
    wire t54009 = t54008 ^ t54008;
    wire t54010 = t54009 ^ t54009;
    wire t54011 = t54010 ^ t54010;
    wire t54012 = t54011 ^ t54011;
    wire t54013 = t54012 ^ t54012;
    wire t54014 = t54013 ^ t54013;
    wire t54015 = t54014 ^ t54014;
    wire t54016 = t54015 ^ t54015;
    wire t54017 = t54016 ^ t54016;
    wire t54018 = t54017 ^ t54017;
    wire t54019 = t54018 ^ t54018;
    wire t54020 = t54019 ^ t54019;
    wire t54021 = t54020 ^ t54020;
    wire t54022 = t54021 ^ t54021;
    wire t54023 = t54022 ^ t54022;
    wire t54024 = t54023 ^ t54023;
    wire t54025 = t54024 ^ t54024;
    wire t54026 = t54025 ^ t54025;
    wire t54027 = t54026 ^ t54026;
    wire t54028 = t54027 ^ t54027;
    wire t54029 = t54028 ^ t54028;
    wire t54030 = t54029 ^ t54029;
    wire t54031 = t54030 ^ t54030;
    wire t54032 = t54031 ^ t54031;
    wire t54033 = t54032 ^ t54032;
    wire t54034 = t54033 ^ t54033;
    wire t54035 = t54034 ^ t54034;
    wire t54036 = t54035 ^ t54035;
    wire t54037 = t54036 ^ t54036;
    wire t54038 = t54037 ^ t54037;
    wire t54039 = t54038 ^ t54038;
    wire t54040 = t54039 ^ t54039;
    wire t54041 = t54040 ^ t54040;
    wire t54042 = t54041 ^ t54041;
    wire t54043 = t54042 ^ t54042;
    wire t54044 = t54043 ^ t54043;
    wire t54045 = t54044 ^ t54044;
    wire t54046 = t54045 ^ t54045;
    wire t54047 = t54046 ^ t54046;
    wire t54048 = t54047 ^ t54047;
    wire t54049 = t54048 ^ t54048;
    wire t54050 = t54049 ^ t54049;
    wire t54051 = t54050 ^ t54050;
    wire t54052 = t54051 ^ t54051;
    wire t54053 = t54052 ^ t54052;
    wire t54054 = t54053 ^ t54053;
    wire t54055 = t54054 ^ t54054;
    wire t54056 = t54055 ^ t54055;
    wire t54057 = t54056 ^ t54056;
    wire t54058 = t54057 ^ t54057;
    wire t54059 = t54058 ^ t54058;
    wire t54060 = t54059 ^ t54059;
    wire t54061 = t54060 ^ t54060;
    wire t54062 = t54061 ^ t54061;
    wire t54063 = t54062 ^ t54062;
    wire t54064 = t54063 ^ t54063;
    wire t54065 = t54064 ^ t54064;
    wire t54066 = t54065 ^ t54065;
    wire t54067 = t54066 ^ t54066;
    wire t54068 = t54067 ^ t54067;
    wire t54069 = t54068 ^ t54068;
    wire t54070 = t54069 ^ t54069;
    wire t54071 = t54070 ^ t54070;
    wire t54072 = t54071 ^ t54071;
    wire t54073 = t54072 ^ t54072;
    wire t54074 = t54073 ^ t54073;
    wire t54075 = t54074 ^ t54074;
    wire t54076 = t54075 ^ t54075;
    wire t54077 = t54076 ^ t54076;
    wire t54078 = t54077 ^ t54077;
    wire t54079 = t54078 ^ t54078;
    wire t54080 = t54079 ^ t54079;
    wire t54081 = t54080 ^ t54080;
    wire t54082 = t54081 ^ t54081;
    wire t54083 = t54082 ^ t54082;
    wire t54084 = t54083 ^ t54083;
    wire t54085 = t54084 ^ t54084;
    wire t54086 = t54085 ^ t54085;
    wire t54087 = t54086 ^ t54086;
    wire t54088 = t54087 ^ t54087;
    wire t54089 = t54088 ^ t54088;
    wire t54090 = t54089 ^ t54089;
    wire t54091 = t54090 ^ t54090;
    wire t54092 = t54091 ^ t54091;
    wire t54093 = t54092 ^ t54092;
    wire t54094 = t54093 ^ t54093;
    wire t54095 = t54094 ^ t54094;
    wire t54096 = t54095 ^ t54095;
    wire t54097 = t54096 ^ t54096;
    wire t54098 = t54097 ^ t54097;
    wire t54099 = t54098 ^ t54098;
    wire t54100 = t54099 ^ t54099;
    wire t54101 = t54100 ^ t54100;
    wire t54102 = t54101 ^ t54101;
    wire t54103 = t54102 ^ t54102;
    wire t54104 = t54103 ^ t54103;
    wire t54105 = t54104 ^ t54104;
    wire t54106 = t54105 ^ t54105;
    wire t54107 = t54106 ^ t54106;
    wire t54108 = t54107 ^ t54107;
    wire t54109 = t54108 ^ t54108;
    wire t54110 = t54109 ^ t54109;
    wire t54111 = t54110 ^ t54110;
    wire t54112 = t54111 ^ t54111;
    wire t54113 = t54112 ^ t54112;
    wire t54114 = t54113 ^ t54113;
    wire t54115 = t54114 ^ t54114;
    wire t54116 = t54115 ^ t54115;
    wire t54117 = t54116 ^ t54116;
    wire t54118 = t54117 ^ t54117;
    wire t54119 = t54118 ^ t54118;
    wire t54120 = t54119 ^ t54119;
    wire t54121 = t54120 ^ t54120;
    wire t54122 = t54121 ^ t54121;
    wire t54123 = t54122 ^ t54122;
    wire t54124 = t54123 ^ t54123;
    wire t54125 = t54124 ^ t54124;
    wire t54126 = t54125 ^ t54125;
    wire t54127 = t54126 ^ t54126;
    wire t54128 = t54127 ^ t54127;
    wire t54129 = t54128 ^ t54128;
    wire t54130 = t54129 ^ t54129;
    wire t54131 = t54130 ^ t54130;
    wire t54132 = t54131 ^ t54131;
    wire t54133 = t54132 ^ t54132;
    wire t54134 = t54133 ^ t54133;
    wire t54135 = t54134 ^ t54134;
    wire t54136 = t54135 ^ t54135;
    wire t54137 = t54136 ^ t54136;
    wire t54138 = t54137 ^ t54137;
    wire t54139 = t54138 ^ t54138;
    wire t54140 = t54139 ^ t54139;
    wire t54141 = t54140 ^ t54140;
    wire t54142 = t54141 ^ t54141;
    wire t54143 = t54142 ^ t54142;
    wire t54144 = t54143 ^ t54143;
    wire t54145 = t54144 ^ t54144;
    wire t54146 = t54145 ^ t54145;
    wire t54147 = t54146 ^ t54146;
    wire t54148 = t54147 ^ t54147;
    wire t54149 = t54148 ^ t54148;
    wire t54150 = t54149 ^ t54149;
    wire t54151 = t54150 ^ t54150;
    wire t54152 = t54151 ^ t54151;
    wire t54153 = t54152 ^ t54152;
    wire t54154 = t54153 ^ t54153;
    wire t54155 = t54154 ^ t54154;
    wire t54156 = t54155 ^ t54155;
    wire t54157 = t54156 ^ t54156;
    wire t54158 = t54157 ^ t54157;
    wire t54159 = t54158 ^ t54158;
    wire t54160 = t54159 ^ t54159;
    wire t54161 = t54160 ^ t54160;
    wire t54162 = t54161 ^ t54161;
    wire t54163 = t54162 ^ t54162;
    wire t54164 = t54163 ^ t54163;
    wire t54165 = t54164 ^ t54164;
    wire t54166 = t54165 ^ t54165;
    wire t54167 = t54166 ^ t54166;
    wire t54168 = t54167 ^ t54167;
    wire t54169 = t54168 ^ t54168;
    wire t54170 = t54169 ^ t54169;
    wire t54171 = t54170 ^ t54170;
    wire t54172 = t54171 ^ t54171;
    wire t54173 = t54172 ^ t54172;
    wire t54174 = t54173 ^ t54173;
    wire t54175 = t54174 ^ t54174;
    wire t54176 = t54175 ^ t54175;
    wire t54177 = t54176 ^ t54176;
    wire t54178 = t54177 ^ t54177;
    wire t54179 = t54178 ^ t54178;
    wire t54180 = t54179 ^ t54179;
    wire t54181 = t54180 ^ t54180;
    wire t54182 = t54181 ^ t54181;
    wire t54183 = t54182 ^ t54182;
    wire t54184 = t54183 ^ t54183;
    wire t54185 = t54184 ^ t54184;
    wire t54186 = t54185 ^ t54185;
    wire t54187 = t54186 ^ t54186;
    wire t54188 = t54187 ^ t54187;
    wire t54189 = t54188 ^ t54188;
    wire t54190 = t54189 ^ t54189;
    wire t54191 = t54190 ^ t54190;
    wire t54192 = t54191 ^ t54191;
    wire t54193 = t54192 ^ t54192;
    wire t54194 = t54193 ^ t54193;
    wire t54195 = t54194 ^ t54194;
    wire t54196 = t54195 ^ t54195;
    wire t54197 = t54196 ^ t54196;
    wire t54198 = t54197 ^ t54197;
    wire t54199 = t54198 ^ t54198;
    wire t54200 = t54199 ^ t54199;
    wire t54201 = t54200 ^ t54200;
    wire t54202 = t54201 ^ t54201;
    wire t54203 = t54202 ^ t54202;
    wire t54204 = t54203 ^ t54203;
    wire t54205 = t54204 ^ t54204;
    wire t54206 = t54205 ^ t54205;
    wire t54207 = t54206 ^ t54206;
    wire t54208 = t54207 ^ t54207;
    wire t54209 = t54208 ^ t54208;
    wire t54210 = t54209 ^ t54209;
    wire t54211 = t54210 ^ t54210;
    wire t54212 = t54211 ^ t54211;
    wire t54213 = t54212 ^ t54212;
    wire t54214 = t54213 ^ t54213;
    wire t54215 = t54214 ^ t54214;
    wire t54216 = t54215 ^ t54215;
    wire t54217 = t54216 ^ t54216;
    wire t54218 = t54217 ^ t54217;
    wire t54219 = t54218 ^ t54218;
    wire t54220 = t54219 ^ t54219;
    wire t54221 = t54220 ^ t54220;
    wire t54222 = t54221 ^ t54221;
    wire t54223 = t54222 ^ t54222;
    wire t54224 = t54223 ^ t54223;
    wire t54225 = t54224 ^ t54224;
    wire t54226 = t54225 ^ t54225;
    wire t54227 = t54226 ^ t54226;
    wire t54228 = t54227 ^ t54227;
    wire t54229 = t54228 ^ t54228;
    wire t54230 = t54229 ^ t54229;
    wire t54231 = t54230 ^ t54230;
    wire t54232 = t54231 ^ t54231;
    wire t54233 = t54232 ^ t54232;
    wire t54234 = t54233 ^ t54233;
    wire t54235 = t54234 ^ t54234;
    wire t54236 = t54235 ^ t54235;
    wire t54237 = t54236 ^ t54236;
    wire t54238 = t54237 ^ t54237;
    wire t54239 = t54238 ^ t54238;
    wire t54240 = t54239 ^ t54239;
    wire t54241 = t54240 ^ t54240;
    wire t54242 = t54241 ^ t54241;
    wire t54243 = t54242 ^ t54242;
    wire t54244 = t54243 ^ t54243;
    wire t54245 = t54244 ^ t54244;
    wire t54246 = t54245 ^ t54245;
    wire t54247 = t54246 ^ t54246;
    wire t54248 = t54247 ^ t54247;
    wire t54249 = t54248 ^ t54248;
    wire t54250 = t54249 ^ t54249;
    wire t54251 = t54250 ^ t54250;
    wire t54252 = t54251 ^ t54251;
    wire t54253 = t54252 ^ t54252;
    wire t54254 = t54253 ^ t54253;
    wire t54255 = t54254 ^ t54254;
    wire t54256 = t54255 ^ t54255;
    wire t54257 = t54256 ^ t54256;
    wire t54258 = t54257 ^ t54257;
    wire t54259 = t54258 ^ t54258;
    wire t54260 = t54259 ^ t54259;
    wire t54261 = t54260 ^ t54260;
    wire t54262 = t54261 ^ t54261;
    wire t54263 = t54262 ^ t54262;
    wire t54264 = t54263 ^ t54263;
    wire t54265 = t54264 ^ t54264;
    wire t54266 = t54265 ^ t54265;
    wire t54267 = t54266 ^ t54266;
    wire t54268 = t54267 ^ t54267;
    wire t54269 = t54268 ^ t54268;
    wire t54270 = t54269 ^ t54269;
    wire t54271 = t54270 ^ t54270;
    wire t54272 = t54271 ^ t54271;
    wire t54273 = t54272 ^ t54272;
    wire t54274 = t54273 ^ t54273;
    wire t54275 = t54274 ^ t54274;
    wire t54276 = t54275 ^ t54275;
    wire t54277 = t54276 ^ t54276;
    wire t54278 = t54277 ^ t54277;
    wire t54279 = t54278 ^ t54278;
    wire t54280 = t54279 ^ t54279;
    wire t54281 = t54280 ^ t54280;
    wire t54282 = t54281 ^ t54281;
    wire t54283 = t54282 ^ t54282;
    wire t54284 = t54283 ^ t54283;
    wire t54285 = t54284 ^ t54284;
    wire t54286 = t54285 ^ t54285;
    wire t54287 = t54286 ^ t54286;
    wire t54288 = t54287 ^ t54287;
    wire t54289 = t54288 ^ t54288;
    wire t54290 = t54289 ^ t54289;
    wire t54291 = t54290 ^ t54290;
    wire t54292 = t54291 ^ t54291;
    wire t54293 = t54292 ^ t54292;
    wire t54294 = t54293 ^ t54293;
    wire t54295 = t54294 ^ t54294;
    wire t54296 = t54295 ^ t54295;
    wire t54297 = t54296 ^ t54296;
    wire t54298 = t54297 ^ t54297;
    wire t54299 = t54298 ^ t54298;
    wire t54300 = t54299 ^ t54299;
    wire t54301 = t54300 ^ t54300;
    wire t54302 = t54301 ^ t54301;
    wire t54303 = t54302 ^ t54302;
    wire t54304 = t54303 ^ t54303;
    wire t54305 = t54304 ^ t54304;
    wire t54306 = t54305 ^ t54305;
    wire t54307 = t54306 ^ t54306;
    wire t54308 = t54307 ^ t54307;
    wire t54309 = t54308 ^ t54308;
    wire t54310 = t54309 ^ t54309;
    wire t54311 = t54310 ^ t54310;
    wire t54312 = t54311 ^ t54311;
    wire t54313 = t54312 ^ t54312;
    wire t54314 = t54313 ^ t54313;
    wire t54315 = t54314 ^ t54314;
    wire t54316 = t54315 ^ t54315;
    wire t54317 = t54316 ^ t54316;
    wire t54318 = t54317 ^ t54317;
    wire t54319 = t54318 ^ t54318;
    wire t54320 = t54319 ^ t54319;
    wire t54321 = t54320 ^ t54320;
    wire t54322 = t54321 ^ t54321;
    wire t54323 = t54322 ^ t54322;
    wire t54324 = t54323 ^ t54323;
    wire t54325 = t54324 ^ t54324;
    wire t54326 = t54325 ^ t54325;
    wire t54327 = t54326 ^ t54326;
    wire t54328 = t54327 ^ t54327;
    wire t54329 = t54328 ^ t54328;
    wire t54330 = t54329 ^ t54329;
    wire t54331 = t54330 ^ t54330;
    wire t54332 = t54331 ^ t54331;
    wire t54333 = t54332 ^ t54332;
    wire t54334 = t54333 ^ t54333;
    wire t54335 = t54334 ^ t54334;
    wire t54336 = t54335 ^ t54335;
    wire t54337 = t54336 ^ t54336;
    wire t54338 = t54337 ^ t54337;
    wire t54339 = t54338 ^ t54338;
    wire t54340 = t54339 ^ t54339;
    wire t54341 = t54340 ^ t54340;
    wire t54342 = t54341 ^ t54341;
    wire t54343 = t54342 ^ t54342;
    wire t54344 = t54343 ^ t54343;
    wire t54345 = t54344 ^ t54344;
    wire t54346 = t54345 ^ t54345;
    wire t54347 = t54346 ^ t54346;
    wire t54348 = t54347 ^ t54347;
    wire t54349 = t54348 ^ t54348;
    wire t54350 = t54349 ^ t54349;
    wire t54351 = t54350 ^ t54350;
    wire t54352 = t54351 ^ t54351;
    wire t54353 = t54352 ^ t54352;
    wire t54354 = t54353 ^ t54353;
    wire t54355 = t54354 ^ t54354;
    wire t54356 = t54355 ^ t54355;
    wire t54357 = t54356 ^ t54356;
    wire t54358 = t54357 ^ t54357;
    wire t54359 = t54358 ^ t54358;
    wire t54360 = t54359 ^ t54359;
    wire t54361 = t54360 ^ t54360;
    wire t54362 = t54361 ^ t54361;
    wire t54363 = t54362 ^ t54362;
    wire t54364 = t54363 ^ t54363;
    wire t54365 = t54364 ^ t54364;
    wire t54366 = t54365 ^ t54365;
    wire t54367 = t54366 ^ t54366;
    wire t54368 = t54367 ^ t54367;
    wire t54369 = t54368 ^ t54368;
    wire t54370 = t54369 ^ t54369;
    wire t54371 = t54370 ^ t54370;
    wire t54372 = t54371 ^ t54371;
    wire t54373 = t54372 ^ t54372;
    wire t54374 = t54373 ^ t54373;
    wire t54375 = t54374 ^ t54374;
    wire t54376 = t54375 ^ t54375;
    wire t54377 = t54376 ^ t54376;
    wire t54378 = t54377 ^ t54377;
    wire t54379 = t54378 ^ t54378;
    wire t54380 = t54379 ^ t54379;
    wire t54381 = t54380 ^ t54380;
    wire t54382 = t54381 ^ t54381;
    wire t54383 = t54382 ^ t54382;
    wire t54384 = t54383 ^ t54383;
    wire t54385 = t54384 ^ t54384;
    wire t54386 = t54385 ^ t54385;
    wire t54387 = t54386 ^ t54386;
    wire t54388 = t54387 ^ t54387;
    wire t54389 = t54388 ^ t54388;
    wire t54390 = t54389 ^ t54389;
    wire t54391 = t54390 ^ t54390;
    wire t54392 = t54391 ^ t54391;
    wire t54393 = t54392 ^ t54392;
    wire t54394 = t54393 ^ t54393;
    wire t54395 = t54394 ^ t54394;
    wire t54396 = t54395 ^ t54395;
    wire t54397 = t54396 ^ t54396;
    wire t54398 = t54397 ^ t54397;
    wire t54399 = t54398 ^ t54398;
    wire t54400 = t54399 ^ t54399;
    wire t54401 = t54400 ^ t54400;
    wire t54402 = t54401 ^ t54401;
    wire t54403 = t54402 ^ t54402;
    wire t54404 = t54403 ^ t54403;
    wire t54405 = t54404 ^ t54404;
    wire t54406 = t54405 ^ t54405;
    wire t54407 = t54406 ^ t54406;
    wire t54408 = t54407 ^ t54407;
    wire t54409 = t54408 ^ t54408;
    wire t54410 = t54409 ^ t54409;
    wire t54411 = t54410 ^ t54410;
    wire t54412 = t54411 ^ t54411;
    wire t54413 = t54412 ^ t54412;
    wire t54414 = t54413 ^ t54413;
    wire t54415 = t54414 ^ t54414;
    wire t54416 = t54415 ^ t54415;
    wire t54417 = t54416 ^ t54416;
    wire t54418 = t54417 ^ t54417;
    wire t54419 = t54418 ^ t54418;
    wire t54420 = t54419 ^ t54419;
    wire t54421 = t54420 ^ t54420;
    wire t54422 = t54421 ^ t54421;
    wire t54423 = t54422 ^ t54422;
    wire t54424 = t54423 ^ t54423;
    wire t54425 = t54424 ^ t54424;
    wire t54426 = t54425 ^ t54425;
    wire t54427 = t54426 ^ t54426;
    wire t54428 = t54427 ^ t54427;
    wire t54429 = t54428 ^ t54428;
    wire t54430 = t54429 ^ t54429;
    wire t54431 = t54430 ^ t54430;
    wire t54432 = t54431 ^ t54431;
    wire t54433 = t54432 ^ t54432;
    wire t54434 = t54433 ^ t54433;
    wire t54435 = t54434 ^ t54434;
    wire t54436 = t54435 ^ t54435;
    wire t54437 = t54436 ^ t54436;
    wire t54438 = t54437 ^ t54437;
    wire t54439 = t54438 ^ t54438;
    wire t54440 = t54439 ^ t54439;
    wire t54441 = t54440 ^ t54440;
    wire t54442 = t54441 ^ t54441;
    wire t54443 = t54442 ^ t54442;
    wire t54444 = t54443 ^ t54443;
    wire t54445 = t54444 ^ t54444;
    wire t54446 = t54445 ^ t54445;
    wire t54447 = t54446 ^ t54446;
    wire t54448 = t54447 ^ t54447;
    wire t54449 = t54448 ^ t54448;
    wire t54450 = t54449 ^ t54449;
    wire t54451 = t54450 ^ t54450;
    wire t54452 = t54451 ^ t54451;
    wire t54453 = t54452 ^ t54452;
    wire t54454 = t54453 ^ t54453;
    wire t54455 = t54454 ^ t54454;
    wire t54456 = t54455 ^ t54455;
    wire t54457 = t54456 ^ t54456;
    wire t54458 = t54457 ^ t54457;
    wire t54459 = t54458 ^ t54458;
    wire t54460 = t54459 ^ t54459;
    wire t54461 = t54460 ^ t54460;
    wire t54462 = t54461 ^ t54461;
    wire t54463 = t54462 ^ t54462;
    wire t54464 = t54463 ^ t54463;
    wire t54465 = t54464 ^ t54464;
    wire t54466 = t54465 ^ t54465;
    wire t54467 = t54466 ^ t54466;
    wire t54468 = t54467 ^ t54467;
    wire t54469 = t54468 ^ t54468;
    wire t54470 = t54469 ^ t54469;
    wire t54471 = t54470 ^ t54470;
    wire t54472 = t54471 ^ t54471;
    wire t54473 = t54472 ^ t54472;
    wire t54474 = t54473 ^ t54473;
    wire t54475 = t54474 ^ t54474;
    wire t54476 = t54475 ^ t54475;
    wire t54477 = t54476 ^ t54476;
    wire t54478 = t54477 ^ t54477;
    wire t54479 = t54478 ^ t54478;
    wire t54480 = t54479 ^ t54479;
    wire t54481 = t54480 ^ t54480;
    wire t54482 = t54481 ^ t54481;
    wire t54483 = t54482 ^ t54482;
    wire t54484 = t54483 ^ t54483;
    wire t54485 = t54484 ^ t54484;
    wire t54486 = t54485 ^ t54485;
    wire t54487 = t54486 ^ t54486;
    wire t54488 = t54487 ^ t54487;
    wire t54489 = t54488 ^ t54488;
    wire t54490 = t54489 ^ t54489;
    wire t54491 = t54490 ^ t54490;
    wire t54492 = t54491 ^ t54491;
    wire t54493 = t54492 ^ t54492;
    wire t54494 = t54493 ^ t54493;
    wire t54495 = t54494 ^ t54494;
    wire t54496 = t54495 ^ t54495;
    wire t54497 = t54496 ^ t54496;
    wire t54498 = t54497 ^ t54497;
    wire t54499 = t54498 ^ t54498;
    wire t54500 = t54499 ^ t54499;
    wire t54501 = t54500 ^ t54500;
    wire t54502 = t54501 ^ t54501;
    wire t54503 = t54502 ^ t54502;
    wire t54504 = t54503 ^ t54503;
    wire t54505 = t54504 ^ t54504;
    wire t54506 = t54505 ^ t54505;
    wire t54507 = t54506 ^ t54506;
    wire t54508 = t54507 ^ t54507;
    wire t54509 = t54508 ^ t54508;
    wire t54510 = t54509 ^ t54509;
    wire t54511 = t54510 ^ t54510;
    wire t54512 = t54511 ^ t54511;
    wire t54513 = t54512 ^ t54512;
    wire t54514 = t54513 ^ t54513;
    wire t54515 = t54514 ^ t54514;
    wire t54516 = t54515 ^ t54515;
    wire t54517 = t54516 ^ t54516;
    wire t54518 = t54517 ^ t54517;
    wire t54519 = t54518 ^ t54518;
    wire t54520 = t54519 ^ t54519;
    wire t54521 = t54520 ^ t54520;
    wire t54522 = t54521 ^ t54521;
    wire t54523 = t54522 ^ t54522;
    wire t54524 = t54523 ^ t54523;
    wire t54525 = t54524 ^ t54524;
    wire t54526 = t54525 ^ t54525;
    wire t54527 = t54526 ^ t54526;
    wire t54528 = t54527 ^ t54527;
    wire t54529 = t54528 ^ t54528;
    wire t54530 = t54529 ^ t54529;
    wire t54531 = t54530 ^ t54530;
    wire t54532 = t54531 ^ t54531;
    wire t54533 = t54532 ^ t54532;
    wire t54534 = t54533 ^ t54533;
    wire t54535 = t54534 ^ t54534;
    wire t54536 = t54535 ^ t54535;
    wire t54537 = t54536 ^ t54536;
    wire t54538 = t54537 ^ t54537;
    wire t54539 = t54538 ^ t54538;
    wire t54540 = t54539 ^ t54539;
    wire t54541 = t54540 ^ t54540;
    wire t54542 = t54541 ^ t54541;
    wire t54543 = t54542 ^ t54542;
    wire t54544 = t54543 ^ t54543;
    wire t54545 = t54544 ^ t54544;
    wire t54546 = t54545 ^ t54545;
    wire t54547 = t54546 ^ t54546;
    wire t54548 = t54547 ^ t54547;
    wire t54549 = t54548 ^ t54548;
    wire t54550 = t54549 ^ t54549;
    wire t54551 = t54550 ^ t54550;
    wire t54552 = t54551 ^ t54551;
    wire t54553 = t54552 ^ t54552;
    wire t54554 = t54553 ^ t54553;
    wire t54555 = t54554 ^ t54554;
    wire t54556 = t54555 ^ t54555;
    wire t54557 = t54556 ^ t54556;
    wire t54558 = t54557 ^ t54557;
    wire t54559 = t54558 ^ t54558;
    wire t54560 = t54559 ^ t54559;
    wire t54561 = t54560 ^ t54560;
    wire t54562 = t54561 ^ t54561;
    wire t54563 = t54562 ^ t54562;
    wire t54564 = t54563 ^ t54563;
    wire t54565 = t54564 ^ t54564;
    wire t54566 = t54565 ^ t54565;
    wire t54567 = t54566 ^ t54566;
    wire t54568 = t54567 ^ t54567;
    wire t54569 = t54568 ^ t54568;
    wire t54570 = t54569 ^ t54569;
    wire t54571 = t54570 ^ t54570;
    wire t54572 = t54571 ^ t54571;
    wire t54573 = t54572 ^ t54572;
    wire t54574 = t54573 ^ t54573;
    wire t54575 = t54574 ^ t54574;
    wire t54576 = t54575 ^ t54575;
    wire t54577 = t54576 ^ t54576;
    wire t54578 = t54577 ^ t54577;
    wire t54579 = t54578 ^ t54578;
    wire t54580 = t54579 ^ t54579;
    wire t54581 = t54580 ^ t54580;
    wire t54582 = t54581 ^ t54581;
    wire t54583 = t54582 ^ t54582;
    wire t54584 = t54583 ^ t54583;
    wire t54585 = t54584 ^ t54584;
    wire t54586 = t54585 ^ t54585;
    wire t54587 = t54586 ^ t54586;
    wire t54588 = t54587 ^ t54587;
    wire t54589 = t54588 ^ t54588;
    wire t54590 = t54589 ^ t54589;
    wire t54591 = t54590 ^ t54590;
    wire t54592 = t54591 ^ t54591;
    wire t54593 = t54592 ^ t54592;
    wire t54594 = t54593 ^ t54593;
    wire t54595 = t54594 ^ t54594;
    wire t54596 = t54595 ^ t54595;
    wire t54597 = t54596 ^ t54596;
    wire t54598 = t54597 ^ t54597;
    wire t54599 = t54598 ^ t54598;
    wire t54600 = t54599 ^ t54599;
    wire t54601 = t54600 ^ t54600;
    wire t54602 = t54601 ^ t54601;
    wire t54603 = t54602 ^ t54602;
    wire t54604 = t54603 ^ t54603;
    wire t54605 = t54604 ^ t54604;
    wire t54606 = t54605 ^ t54605;
    wire t54607 = t54606 ^ t54606;
    wire t54608 = t54607 ^ t54607;
    wire t54609 = t54608 ^ t54608;
    wire t54610 = t54609 ^ t54609;
    wire t54611 = t54610 ^ t54610;
    wire t54612 = t54611 ^ t54611;
    wire t54613 = t54612 ^ t54612;
    wire t54614 = t54613 ^ t54613;
    wire t54615 = t54614 ^ t54614;
    wire t54616 = t54615 ^ t54615;
    wire t54617 = t54616 ^ t54616;
    wire t54618 = t54617 ^ t54617;
    wire t54619 = t54618 ^ t54618;
    wire t54620 = t54619 ^ t54619;
    wire t54621 = t54620 ^ t54620;
    wire t54622 = t54621 ^ t54621;
    wire t54623 = t54622 ^ t54622;
    wire t54624 = t54623 ^ t54623;
    wire t54625 = t54624 ^ t54624;
    wire t54626 = t54625 ^ t54625;
    wire t54627 = t54626 ^ t54626;
    wire t54628 = t54627 ^ t54627;
    wire t54629 = t54628 ^ t54628;
    wire t54630 = t54629 ^ t54629;
    wire t54631 = t54630 ^ t54630;
    wire t54632 = t54631 ^ t54631;
    wire t54633 = t54632 ^ t54632;
    wire t54634 = t54633 ^ t54633;
    wire t54635 = t54634 ^ t54634;
    wire t54636 = t54635 ^ t54635;
    wire t54637 = t54636 ^ t54636;
    wire t54638 = t54637 ^ t54637;
    wire t54639 = t54638 ^ t54638;
    wire t54640 = t54639 ^ t54639;
    wire t54641 = t54640 ^ t54640;
    wire t54642 = t54641 ^ t54641;
    wire t54643 = t54642 ^ t54642;
    wire t54644 = t54643 ^ t54643;
    wire t54645 = t54644 ^ t54644;
    wire t54646 = t54645 ^ t54645;
    wire t54647 = t54646 ^ t54646;
    wire t54648 = t54647 ^ t54647;
    wire t54649 = t54648 ^ t54648;
    wire t54650 = t54649 ^ t54649;
    wire t54651 = t54650 ^ t54650;
    wire t54652 = t54651 ^ t54651;
    wire t54653 = t54652 ^ t54652;
    wire t54654 = t54653 ^ t54653;
    wire t54655 = t54654 ^ t54654;
    wire t54656 = t54655 ^ t54655;
    wire t54657 = t54656 ^ t54656;
    wire t54658 = t54657 ^ t54657;
    wire t54659 = t54658 ^ t54658;
    wire t54660 = t54659 ^ t54659;
    wire t54661 = t54660 ^ t54660;
    wire t54662 = t54661 ^ t54661;
    wire t54663 = t54662 ^ t54662;
    wire t54664 = t54663 ^ t54663;
    wire t54665 = t54664 ^ t54664;
    wire t54666 = t54665 ^ t54665;
    wire t54667 = t54666 ^ t54666;
    wire t54668 = t54667 ^ t54667;
    wire t54669 = t54668 ^ t54668;
    wire t54670 = t54669 ^ t54669;
    wire t54671 = t54670 ^ t54670;
    wire t54672 = t54671 ^ t54671;
    wire t54673 = t54672 ^ t54672;
    wire t54674 = t54673 ^ t54673;
    wire t54675 = t54674 ^ t54674;
    wire t54676 = t54675 ^ t54675;
    wire t54677 = t54676 ^ t54676;
    wire t54678 = t54677 ^ t54677;
    wire t54679 = t54678 ^ t54678;
    wire t54680 = t54679 ^ t54679;
    wire t54681 = t54680 ^ t54680;
    wire t54682 = t54681 ^ t54681;
    wire t54683 = t54682 ^ t54682;
    wire t54684 = t54683 ^ t54683;
    wire t54685 = t54684 ^ t54684;
    wire t54686 = t54685 ^ t54685;
    wire t54687 = t54686 ^ t54686;
    wire t54688 = t54687 ^ t54687;
    wire t54689 = t54688 ^ t54688;
    wire t54690 = t54689 ^ t54689;
    wire t54691 = t54690 ^ t54690;
    wire t54692 = t54691 ^ t54691;
    wire t54693 = t54692 ^ t54692;
    wire t54694 = t54693 ^ t54693;
    wire t54695 = t54694 ^ t54694;
    wire t54696 = t54695 ^ t54695;
    wire t54697 = t54696 ^ t54696;
    wire t54698 = t54697 ^ t54697;
    wire t54699 = t54698 ^ t54698;
    wire t54700 = t54699 ^ t54699;
    wire t54701 = t54700 ^ t54700;
    wire t54702 = t54701 ^ t54701;
    wire t54703 = t54702 ^ t54702;
    wire t54704 = t54703 ^ t54703;
    wire t54705 = t54704 ^ t54704;
    wire t54706 = t54705 ^ t54705;
    wire t54707 = t54706 ^ t54706;
    wire t54708 = t54707 ^ t54707;
    wire t54709 = t54708 ^ t54708;
    wire t54710 = t54709 ^ t54709;
    wire t54711 = t54710 ^ t54710;
    wire t54712 = t54711 ^ t54711;
    wire t54713 = t54712 ^ t54712;
    wire t54714 = t54713 ^ t54713;
    wire t54715 = t54714 ^ t54714;
    wire t54716 = t54715 ^ t54715;
    wire t54717 = t54716 ^ t54716;
    wire t54718 = t54717 ^ t54717;
    wire t54719 = t54718 ^ t54718;
    wire t54720 = t54719 ^ t54719;
    wire t54721 = t54720 ^ t54720;
    wire t54722 = t54721 ^ t54721;
    wire t54723 = t54722 ^ t54722;
    wire t54724 = t54723 ^ t54723;
    wire t54725 = t54724 ^ t54724;
    wire t54726 = t54725 ^ t54725;
    wire t54727 = t54726 ^ t54726;
    wire t54728 = t54727 ^ t54727;
    wire t54729 = t54728 ^ t54728;
    wire t54730 = t54729 ^ t54729;
    wire t54731 = t54730 ^ t54730;
    wire t54732 = t54731 ^ t54731;
    wire t54733 = t54732 ^ t54732;
    wire t54734 = t54733 ^ t54733;
    wire t54735 = t54734 ^ t54734;
    wire t54736 = t54735 ^ t54735;
    wire t54737 = t54736 ^ t54736;
    wire t54738 = t54737 ^ t54737;
    wire t54739 = t54738 ^ t54738;
    wire t54740 = t54739 ^ t54739;
    wire t54741 = t54740 ^ t54740;
    wire t54742 = t54741 ^ t54741;
    wire t54743 = t54742 ^ t54742;
    wire t54744 = t54743 ^ t54743;
    wire t54745 = t54744 ^ t54744;
    wire t54746 = t54745 ^ t54745;
    wire t54747 = t54746 ^ t54746;
    wire t54748 = t54747 ^ t54747;
    wire t54749 = t54748 ^ t54748;
    wire t54750 = t54749 ^ t54749;
    wire t54751 = t54750 ^ t54750;
    wire t54752 = t54751 ^ t54751;
    wire t54753 = t54752 ^ t54752;
    wire t54754 = t54753 ^ t54753;
    wire t54755 = t54754 ^ t54754;
    wire t54756 = t54755 ^ t54755;
    wire t54757 = t54756 ^ t54756;
    wire t54758 = t54757 ^ t54757;
    wire t54759 = t54758 ^ t54758;
    wire t54760 = t54759 ^ t54759;
    wire t54761 = t54760 ^ t54760;
    wire t54762 = t54761 ^ t54761;
    wire t54763 = t54762 ^ t54762;
    wire t54764 = t54763 ^ t54763;
    wire t54765 = t54764 ^ t54764;
    wire t54766 = t54765 ^ t54765;
    wire t54767 = t54766 ^ t54766;
    wire t54768 = t54767 ^ t54767;
    wire t54769 = t54768 ^ t54768;
    wire t54770 = t54769 ^ t54769;
    wire t54771 = t54770 ^ t54770;
    wire t54772 = t54771 ^ t54771;
    wire t54773 = t54772 ^ t54772;
    wire t54774 = t54773 ^ t54773;
    wire t54775 = t54774 ^ t54774;
    wire t54776 = t54775 ^ t54775;
    wire t54777 = t54776 ^ t54776;
    wire t54778 = t54777 ^ t54777;
    wire t54779 = t54778 ^ t54778;
    wire t54780 = t54779 ^ t54779;
    wire t54781 = t54780 ^ t54780;
    wire t54782 = t54781 ^ t54781;
    wire t54783 = t54782 ^ t54782;
    wire t54784 = t54783 ^ t54783;
    wire t54785 = t54784 ^ t54784;
    wire t54786 = t54785 ^ t54785;
    wire t54787 = t54786 ^ t54786;
    wire t54788 = t54787 ^ t54787;
    wire t54789 = t54788 ^ t54788;
    wire t54790 = t54789 ^ t54789;
    wire t54791 = t54790 ^ t54790;
    wire t54792 = t54791 ^ t54791;
    wire t54793 = t54792 ^ t54792;
    wire t54794 = t54793 ^ t54793;
    wire t54795 = t54794 ^ t54794;
    wire t54796 = t54795 ^ t54795;
    wire t54797 = t54796 ^ t54796;
    wire t54798 = t54797 ^ t54797;
    wire t54799 = t54798 ^ t54798;
    wire t54800 = t54799 ^ t54799;
    wire t54801 = t54800 ^ t54800;
    wire t54802 = t54801 ^ t54801;
    wire t54803 = t54802 ^ t54802;
    wire t54804 = t54803 ^ t54803;
    wire t54805 = t54804 ^ t54804;
    wire t54806 = t54805 ^ t54805;
    wire t54807 = t54806 ^ t54806;
    wire t54808 = t54807 ^ t54807;
    wire t54809 = t54808 ^ t54808;
    wire t54810 = t54809 ^ t54809;
    wire t54811 = t54810 ^ t54810;
    wire t54812 = t54811 ^ t54811;
    wire t54813 = t54812 ^ t54812;
    wire t54814 = t54813 ^ t54813;
    wire t54815 = t54814 ^ t54814;
    wire t54816 = t54815 ^ t54815;
    wire t54817 = t54816 ^ t54816;
    wire t54818 = t54817 ^ t54817;
    wire t54819 = t54818 ^ t54818;
    wire t54820 = t54819 ^ t54819;
    wire t54821 = t54820 ^ t54820;
    wire t54822 = t54821 ^ t54821;
    wire t54823 = t54822 ^ t54822;
    wire t54824 = t54823 ^ t54823;
    wire t54825 = t54824 ^ t54824;
    wire t54826 = t54825 ^ t54825;
    wire t54827 = t54826 ^ t54826;
    wire t54828 = t54827 ^ t54827;
    wire t54829 = t54828 ^ t54828;
    wire t54830 = t54829 ^ t54829;
    wire t54831 = t54830 ^ t54830;
    wire t54832 = t54831 ^ t54831;
    wire t54833 = t54832 ^ t54832;
    wire t54834 = t54833 ^ t54833;
    wire t54835 = t54834 ^ t54834;
    wire t54836 = t54835 ^ t54835;
    wire t54837 = t54836 ^ t54836;
    wire t54838 = t54837 ^ t54837;
    wire t54839 = t54838 ^ t54838;
    wire t54840 = t54839 ^ t54839;
    wire t54841 = t54840 ^ t54840;
    wire t54842 = t54841 ^ t54841;
    wire t54843 = t54842 ^ t54842;
    wire t54844 = t54843 ^ t54843;
    wire t54845 = t54844 ^ t54844;
    wire t54846 = t54845 ^ t54845;
    wire t54847 = t54846 ^ t54846;
    wire t54848 = t54847 ^ t54847;
    wire t54849 = t54848 ^ t54848;
    wire t54850 = t54849 ^ t54849;
    wire t54851 = t54850 ^ t54850;
    wire t54852 = t54851 ^ t54851;
    wire t54853 = t54852 ^ t54852;
    wire t54854 = t54853 ^ t54853;
    wire t54855 = t54854 ^ t54854;
    wire t54856 = t54855 ^ t54855;
    wire t54857 = t54856 ^ t54856;
    wire t54858 = t54857 ^ t54857;
    wire t54859 = t54858 ^ t54858;
    wire t54860 = t54859 ^ t54859;
    wire t54861 = t54860 ^ t54860;
    wire t54862 = t54861 ^ t54861;
    wire t54863 = t54862 ^ t54862;
    wire t54864 = t54863 ^ t54863;
    wire t54865 = t54864 ^ t54864;
    wire t54866 = t54865 ^ t54865;
    wire t54867 = t54866 ^ t54866;
    wire t54868 = t54867 ^ t54867;
    wire t54869 = t54868 ^ t54868;
    wire t54870 = t54869 ^ t54869;
    wire t54871 = t54870 ^ t54870;
    wire t54872 = t54871 ^ t54871;
    wire t54873 = t54872 ^ t54872;
    wire t54874 = t54873 ^ t54873;
    wire t54875 = t54874 ^ t54874;
    wire t54876 = t54875 ^ t54875;
    wire t54877 = t54876 ^ t54876;
    wire t54878 = t54877 ^ t54877;
    wire t54879 = t54878 ^ t54878;
    wire t54880 = t54879 ^ t54879;
    wire t54881 = t54880 ^ t54880;
    wire t54882 = t54881 ^ t54881;
    wire t54883 = t54882 ^ t54882;
    wire t54884 = t54883 ^ t54883;
    wire t54885 = t54884 ^ t54884;
    wire t54886 = t54885 ^ t54885;
    wire t54887 = t54886 ^ t54886;
    wire t54888 = t54887 ^ t54887;
    wire t54889 = t54888 ^ t54888;
    wire t54890 = t54889 ^ t54889;
    wire t54891 = t54890 ^ t54890;
    wire t54892 = t54891 ^ t54891;
    wire t54893 = t54892 ^ t54892;
    wire t54894 = t54893 ^ t54893;
    wire t54895 = t54894 ^ t54894;
    wire t54896 = t54895 ^ t54895;
    wire t54897 = t54896 ^ t54896;
    wire t54898 = t54897 ^ t54897;
    wire t54899 = t54898 ^ t54898;
    wire t54900 = t54899 ^ t54899;
    wire t54901 = t54900 ^ t54900;
    wire t54902 = t54901 ^ t54901;
    wire t54903 = t54902 ^ t54902;
    wire t54904 = t54903 ^ t54903;
    wire t54905 = t54904 ^ t54904;
    wire t54906 = t54905 ^ t54905;
    wire t54907 = t54906 ^ t54906;
    wire t54908 = t54907 ^ t54907;
    wire t54909 = t54908 ^ t54908;
    wire t54910 = t54909 ^ t54909;
    wire t54911 = t54910 ^ t54910;
    wire t54912 = t54911 ^ t54911;
    wire t54913 = t54912 ^ t54912;
    wire t54914 = t54913 ^ t54913;
    wire t54915 = t54914 ^ t54914;
    wire t54916 = t54915 ^ t54915;
    wire t54917 = t54916 ^ t54916;
    wire t54918 = t54917 ^ t54917;
    wire t54919 = t54918 ^ t54918;
    wire t54920 = t54919 ^ t54919;
    wire t54921 = t54920 ^ t54920;
    wire t54922 = t54921 ^ t54921;
    wire t54923 = t54922 ^ t54922;
    wire t54924 = t54923 ^ t54923;
    wire t54925 = t54924 ^ t54924;
    wire t54926 = t54925 ^ t54925;
    wire t54927 = t54926 ^ t54926;
    wire t54928 = t54927 ^ t54927;
    wire t54929 = t54928 ^ t54928;
    wire t54930 = t54929 ^ t54929;
    wire t54931 = t54930 ^ t54930;
    wire t54932 = t54931 ^ t54931;
    wire t54933 = t54932 ^ t54932;
    wire t54934 = t54933 ^ t54933;
    wire t54935 = t54934 ^ t54934;
    wire t54936 = t54935 ^ t54935;
    wire t54937 = t54936 ^ t54936;
    wire t54938 = t54937 ^ t54937;
    wire t54939 = t54938 ^ t54938;
    wire t54940 = t54939 ^ t54939;
    wire t54941 = t54940 ^ t54940;
    wire t54942 = t54941 ^ t54941;
    wire t54943 = t54942 ^ t54942;
    wire t54944 = t54943 ^ t54943;
    wire t54945 = t54944 ^ t54944;
    wire t54946 = t54945 ^ t54945;
    wire t54947 = t54946 ^ t54946;
    wire t54948 = t54947 ^ t54947;
    wire t54949 = t54948 ^ t54948;
    wire t54950 = t54949 ^ t54949;
    wire t54951 = t54950 ^ t54950;
    wire t54952 = t54951 ^ t54951;
    wire t54953 = t54952 ^ t54952;
    wire t54954 = t54953 ^ t54953;
    wire t54955 = t54954 ^ t54954;
    wire t54956 = t54955 ^ t54955;
    wire t54957 = t54956 ^ t54956;
    wire t54958 = t54957 ^ t54957;
    wire t54959 = t54958 ^ t54958;
    wire t54960 = t54959 ^ t54959;
    wire t54961 = t54960 ^ t54960;
    wire t54962 = t54961 ^ t54961;
    wire t54963 = t54962 ^ t54962;
    wire t54964 = t54963 ^ t54963;
    wire t54965 = t54964 ^ t54964;
    wire t54966 = t54965 ^ t54965;
    wire t54967 = t54966 ^ t54966;
    wire t54968 = t54967 ^ t54967;
    wire t54969 = t54968 ^ t54968;
    wire t54970 = t54969 ^ t54969;
    wire t54971 = t54970 ^ t54970;
    wire t54972 = t54971 ^ t54971;
    wire t54973 = t54972 ^ t54972;
    wire t54974 = t54973 ^ t54973;
    wire t54975 = t54974 ^ t54974;
    wire t54976 = t54975 ^ t54975;
    wire t54977 = t54976 ^ t54976;
    wire t54978 = t54977 ^ t54977;
    wire t54979 = t54978 ^ t54978;
    wire t54980 = t54979 ^ t54979;
    wire t54981 = t54980 ^ t54980;
    wire t54982 = t54981 ^ t54981;
    wire t54983 = t54982 ^ t54982;
    wire t54984 = t54983 ^ t54983;
    wire t54985 = t54984 ^ t54984;
    wire t54986 = t54985 ^ t54985;
    wire t54987 = t54986 ^ t54986;
    wire t54988 = t54987 ^ t54987;
    wire t54989 = t54988 ^ t54988;
    wire t54990 = t54989 ^ t54989;
    wire t54991 = t54990 ^ t54990;
    wire t54992 = t54991 ^ t54991;
    wire t54993 = t54992 ^ t54992;
    wire t54994 = t54993 ^ t54993;
    wire t54995 = t54994 ^ t54994;
    wire t54996 = t54995 ^ t54995;
    wire t54997 = t54996 ^ t54996;
    wire t54998 = t54997 ^ t54997;
    wire t54999 = t54998 ^ t54998;
    wire t55000 = t54999 ^ t54999;
    wire t55001 = t55000 ^ t55000;
    wire t55002 = t55001 ^ t55001;
    wire t55003 = t55002 ^ t55002;
    wire t55004 = t55003 ^ t55003;
    wire t55005 = t55004 ^ t55004;
    wire t55006 = t55005 ^ t55005;
    wire t55007 = t55006 ^ t55006;
    wire t55008 = t55007 ^ t55007;
    wire t55009 = t55008 ^ t55008;
    wire t55010 = t55009 ^ t55009;
    wire t55011 = t55010 ^ t55010;
    wire t55012 = t55011 ^ t55011;
    wire t55013 = t55012 ^ t55012;
    wire t55014 = t55013 ^ t55013;
    wire t55015 = t55014 ^ t55014;
    wire t55016 = t55015 ^ t55015;
    wire t55017 = t55016 ^ t55016;
    wire t55018 = t55017 ^ t55017;
    wire t55019 = t55018 ^ t55018;
    wire t55020 = t55019 ^ t55019;
    wire t55021 = t55020 ^ t55020;
    wire t55022 = t55021 ^ t55021;
    wire t55023 = t55022 ^ t55022;
    wire t55024 = t55023 ^ t55023;
    wire t55025 = t55024 ^ t55024;
    wire t55026 = t55025 ^ t55025;
    wire t55027 = t55026 ^ t55026;
    wire t55028 = t55027 ^ t55027;
    wire t55029 = t55028 ^ t55028;
    wire t55030 = t55029 ^ t55029;
    wire t55031 = t55030 ^ t55030;
    wire t55032 = t55031 ^ t55031;
    wire t55033 = t55032 ^ t55032;
    wire t55034 = t55033 ^ t55033;
    wire t55035 = t55034 ^ t55034;
    wire t55036 = t55035 ^ t55035;
    wire t55037 = t55036 ^ t55036;
    wire t55038 = t55037 ^ t55037;
    wire t55039 = t55038 ^ t55038;
    wire t55040 = t55039 ^ t55039;
    wire t55041 = t55040 ^ t55040;
    wire t55042 = t55041 ^ t55041;
    wire t55043 = t55042 ^ t55042;
    wire t55044 = t55043 ^ t55043;
    wire t55045 = t55044 ^ t55044;
    wire t55046 = t55045 ^ t55045;
    wire t55047 = t55046 ^ t55046;
    wire t55048 = t55047 ^ t55047;
    wire t55049 = t55048 ^ t55048;
    wire t55050 = t55049 ^ t55049;
    wire t55051 = t55050 ^ t55050;
    wire t55052 = t55051 ^ t55051;
    wire t55053 = t55052 ^ t55052;
    wire t55054 = t55053 ^ t55053;
    wire t55055 = t55054 ^ t55054;
    wire t55056 = t55055 ^ t55055;
    wire t55057 = t55056 ^ t55056;
    wire t55058 = t55057 ^ t55057;
    wire t55059 = t55058 ^ t55058;
    wire t55060 = t55059 ^ t55059;
    wire t55061 = t55060 ^ t55060;
    wire t55062 = t55061 ^ t55061;
    wire t55063 = t55062 ^ t55062;
    wire t55064 = t55063 ^ t55063;
    wire t55065 = t55064 ^ t55064;
    wire t55066 = t55065 ^ t55065;
    wire t55067 = t55066 ^ t55066;
    wire t55068 = t55067 ^ t55067;
    wire t55069 = t55068 ^ t55068;
    wire t55070 = t55069 ^ t55069;
    wire t55071 = t55070 ^ t55070;
    wire t55072 = t55071 ^ t55071;
    wire t55073 = t55072 ^ t55072;
    wire t55074 = t55073 ^ t55073;
    wire t55075 = t55074 ^ t55074;
    wire t55076 = t55075 ^ t55075;
    wire t55077 = t55076 ^ t55076;
    wire t55078 = t55077 ^ t55077;
    wire t55079 = t55078 ^ t55078;
    wire t55080 = t55079 ^ t55079;
    wire t55081 = t55080 ^ t55080;
    wire t55082 = t55081 ^ t55081;
    wire t55083 = t55082 ^ t55082;
    wire t55084 = t55083 ^ t55083;
    wire t55085 = t55084 ^ t55084;
    wire t55086 = t55085 ^ t55085;
    wire t55087 = t55086 ^ t55086;
    wire t55088 = t55087 ^ t55087;
    wire t55089 = t55088 ^ t55088;
    wire t55090 = t55089 ^ t55089;
    wire t55091 = t55090 ^ t55090;
    wire t55092 = t55091 ^ t55091;
    wire t55093 = t55092 ^ t55092;
    wire t55094 = t55093 ^ t55093;
    wire t55095 = t55094 ^ t55094;
    wire t55096 = t55095 ^ t55095;
    wire t55097 = t55096 ^ t55096;
    wire t55098 = t55097 ^ t55097;
    wire t55099 = t55098 ^ t55098;
    wire t55100 = t55099 ^ t55099;
    wire t55101 = t55100 ^ t55100;
    wire t55102 = t55101 ^ t55101;
    wire t55103 = t55102 ^ t55102;
    wire t55104 = t55103 ^ t55103;
    wire t55105 = t55104 ^ t55104;
    wire t55106 = t55105 ^ t55105;
    wire t55107 = t55106 ^ t55106;
    wire t55108 = t55107 ^ t55107;
    wire t55109 = t55108 ^ t55108;
    wire t55110 = t55109 ^ t55109;
    wire t55111 = t55110 ^ t55110;
    wire t55112 = t55111 ^ t55111;
    wire t55113 = t55112 ^ t55112;
    wire t55114 = t55113 ^ t55113;
    wire t55115 = t55114 ^ t55114;
    wire t55116 = t55115 ^ t55115;
    wire t55117 = t55116 ^ t55116;
    wire t55118 = t55117 ^ t55117;
    wire t55119 = t55118 ^ t55118;
    wire t55120 = t55119 ^ t55119;
    wire t55121 = t55120 ^ t55120;
    wire t55122 = t55121 ^ t55121;
    wire t55123 = t55122 ^ t55122;
    wire t55124 = t55123 ^ t55123;
    wire t55125 = t55124 ^ t55124;
    wire t55126 = t55125 ^ t55125;
    wire t55127 = t55126 ^ t55126;
    wire t55128 = t55127 ^ t55127;
    wire t55129 = t55128 ^ t55128;
    wire t55130 = t55129 ^ t55129;
    wire t55131 = t55130 ^ t55130;
    wire t55132 = t55131 ^ t55131;
    wire t55133 = t55132 ^ t55132;
    wire t55134 = t55133 ^ t55133;
    wire t55135 = t55134 ^ t55134;
    wire t55136 = t55135 ^ t55135;
    wire t55137 = t55136 ^ t55136;
    wire t55138 = t55137 ^ t55137;
    wire t55139 = t55138 ^ t55138;
    wire t55140 = t55139 ^ t55139;
    wire t55141 = t55140 ^ t55140;
    wire t55142 = t55141 ^ t55141;
    wire t55143 = t55142 ^ t55142;
    wire t55144 = t55143 ^ t55143;
    wire t55145 = t55144 ^ t55144;
    wire t55146 = t55145 ^ t55145;
    wire t55147 = t55146 ^ t55146;
    wire t55148 = t55147 ^ t55147;
    wire t55149 = t55148 ^ t55148;
    wire t55150 = t55149 ^ t55149;
    wire t55151 = t55150 ^ t55150;
    wire t55152 = t55151 ^ t55151;
    wire t55153 = t55152 ^ t55152;
    wire t55154 = t55153 ^ t55153;
    wire t55155 = t55154 ^ t55154;
    wire t55156 = t55155 ^ t55155;
    wire t55157 = t55156 ^ t55156;
    wire t55158 = t55157 ^ t55157;
    wire t55159 = t55158 ^ t55158;
    wire t55160 = t55159 ^ t55159;
    wire t55161 = t55160 ^ t55160;
    wire t55162 = t55161 ^ t55161;
    wire t55163 = t55162 ^ t55162;
    wire t55164 = t55163 ^ t55163;
    wire t55165 = t55164 ^ t55164;
    wire t55166 = t55165 ^ t55165;
    wire t55167 = t55166 ^ t55166;
    wire t55168 = t55167 ^ t55167;
    wire t55169 = t55168 ^ t55168;
    wire t55170 = t55169 ^ t55169;
    wire t55171 = t55170 ^ t55170;
    wire t55172 = t55171 ^ t55171;
    wire t55173 = t55172 ^ t55172;
    wire t55174 = t55173 ^ t55173;
    wire t55175 = t55174 ^ t55174;
    wire t55176 = t55175 ^ t55175;
    wire t55177 = t55176 ^ t55176;
    wire t55178 = t55177 ^ t55177;
    wire t55179 = t55178 ^ t55178;
    wire t55180 = t55179 ^ t55179;
    wire t55181 = t55180 ^ t55180;
    wire t55182 = t55181 ^ t55181;
    wire t55183 = t55182 ^ t55182;
    wire t55184 = t55183 ^ t55183;
    wire t55185 = t55184 ^ t55184;
    wire t55186 = t55185 ^ t55185;
    wire t55187 = t55186 ^ t55186;
    wire t55188 = t55187 ^ t55187;
    wire t55189 = t55188 ^ t55188;
    wire t55190 = t55189 ^ t55189;
    wire t55191 = t55190 ^ t55190;
    wire t55192 = t55191 ^ t55191;
    wire t55193 = t55192 ^ t55192;
    wire t55194 = t55193 ^ t55193;
    wire t55195 = t55194 ^ t55194;
    wire t55196 = t55195 ^ t55195;
    wire t55197 = t55196 ^ t55196;
    wire t55198 = t55197 ^ t55197;
    wire t55199 = t55198 ^ t55198;
    wire t55200 = t55199 ^ t55199;
    wire t55201 = t55200 ^ t55200;
    wire t55202 = t55201 ^ t55201;
    wire t55203 = t55202 ^ t55202;
    wire t55204 = t55203 ^ t55203;
    wire t55205 = t55204 ^ t55204;
    wire t55206 = t55205 ^ t55205;
    wire t55207 = t55206 ^ t55206;
    wire t55208 = t55207 ^ t55207;
    wire t55209 = t55208 ^ t55208;
    wire t55210 = t55209 ^ t55209;
    wire t55211 = t55210 ^ t55210;
    wire t55212 = t55211 ^ t55211;
    wire t55213 = t55212 ^ t55212;
    wire t55214 = t55213 ^ t55213;
    wire t55215 = t55214 ^ t55214;
    wire t55216 = t55215 ^ t55215;
    wire t55217 = t55216 ^ t55216;
    wire t55218 = t55217 ^ t55217;
    wire t55219 = t55218 ^ t55218;
    wire t55220 = t55219 ^ t55219;
    wire t55221 = t55220 ^ t55220;
    wire t55222 = t55221 ^ t55221;
    wire t55223 = t55222 ^ t55222;
    wire t55224 = t55223 ^ t55223;
    wire t55225 = t55224 ^ t55224;
    wire t55226 = t55225 ^ t55225;
    wire t55227 = t55226 ^ t55226;
    wire t55228 = t55227 ^ t55227;
    wire t55229 = t55228 ^ t55228;
    wire t55230 = t55229 ^ t55229;
    wire t55231 = t55230 ^ t55230;
    wire t55232 = t55231 ^ t55231;
    wire t55233 = t55232 ^ t55232;
    wire t55234 = t55233 ^ t55233;
    wire t55235 = t55234 ^ t55234;
    wire t55236 = t55235 ^ t55235;
    wire t55237 = t55236 ^ t55236;
    wire t55238 = t55237 ^ t55237;
    wire t55239 = t55238 ^ t55238;
    wire t55240 = t55239 ^ t55239;
    wire t55241 = t55240 ^ t55240;
    wire t55242 = t55241 ^ t55241;
    wire t55243 = t55242 ^ t55242;
    wire t55244 = t55243 ^ t55243;
    wire t55245 = t55244 ^ t55244;
    wire t55246 = t55245 ^ t55245;
    wire t55247 = t55246 ^ t55246;
    wire t55248 = t55247 ^ t55247;
    wire t55249 = t55248 ^ t55248;
    wire t55250 = t55249 ^ t55249;
    wire t55251 = t55250 ^ t55250;
    wire t55252 = t55251 ^ t55251;
    wire t55253 = t55252 ^ t55252;
    wire t55254 = t55253 ^ t55253;
    wire t55255 = t55254 ^ t55254;
    wire t55256 = t55255 ^ t55255;
    wire t55257 = t55256 ^ t55256;
    wire t55258 = t55257 ^ t55257;
    wire t55259 = t55258 ^ t55258;
    wire t55260 = t55259 ^ t55259;
    wire t55261 = t55260 ^ t55260;
    wire t55262 = t55261 ^ t55261;
    wire t55263 = t55262 ^ t55262;
    wire t55264 = t55263 ^ t55263;
    wire t55265 = t55264 ^ t55264;
    wire t55266 = t55265 ^ t55265;
    wire t55267 = t55266 ^ t55266;
    wire t55268 = t55267 ^ t55267;
    wire t55269 = t55268 ^ t55268;
    wire t55270 = t55269 ^ t55269;
    wire t55271 = t55270 ^ t55270;
    wire t55272 = t55271 ^ t55271;
    wire t55273 = t55272 ^ t55272;
    wire t55274 = t55273 ^ t55273;
    wire t55275 = t55274 ^ t55274;
    wire t55276 = t55275 ^ t55275;
    wire t55277 = t55276 ^ t55276;
    wire t55278 = t55277 ^ t55277;
    wire t55279 = t55278 ^ t55278;
    wire t55280 = t55279 ^ t55279;
    wire t55281 = t55280 ^ t55280;
    wire t55282 = t55281 ^ t55281;
    wire t55283 = t55282 ^ t55282;
    wire t55284 = t55283 ^ t55283;
    wire t55285 = t55284 ^ t55284;
    wire t55286 = t55285 ^ t55285;
    wire t55287 = t55286 ^ t55286;
    wire t55288 = t55287 ^ t55287;
    wire t55289 = t55288 ^ t55288;
    wire t55290 = t55289 ^ t55289;
    wire t55291 = t55290 ^ t55290;
    wire t55292 = t55291 ^ t55291;
    wire t55293 = t55292 ^ t55292;
    wire t55294 = t55293 ^ t55293;
    wire t55295 = t55294 ^ t55294;
    wire t55296 = t55295 ^ t55295;
    wire t55297 = t55296 ^ t55296;
    wire t55298 = t55297 ^ t55297;
    wire t55299 = t55298 ^ t55298;
    wire t55300 = t55299 ^ t55299;
    wire t55301 = t55300 ^ t55300;
    wire t55302 = t55301 ^ t55301;
    wire t55303 = t55302 ^ t55302;
    wire t55304 = t55303 ^ t55303;
    wire t55305 = t55304 ^ t55304;
    wire t55306 = t55305 ^ t55305;
    wire t55307 = t55306 ^ t55306;
    wire t55308 = t55307 ^ t55307;
    wire t55309 = t55308 ^ t55308;
    wire t55310 = t55309 ^ t55309;
    wire t55311 = t55310 ^ t55310;
    wire t55312 = t55311 ^ t55311;
    wire t55313 = t55312 ^ t55312;
    wire t55314 = t55313 ^ t55313;
    wire t55315 = t55314 ^ t55314;
    wire t55316 = t55315 ^ t55315;
    wire t55317 = t55316 ^ t55316;
    wire t55318 = t55317 ^ t55317;
    wire t55319 = t55318 ^ t55318;
    wire t55320 = t55319 ^ t55319;
    wire t55321 = t55320 ^ t55320;
    wire t55322 = t55321 ^ t55321;
    wire t55323 = t55322 ^ t55322;
    wire t55324 = t55323 ^ t55323;
    wire t55325 = t55324 ^ t55324;
    wire t55326 = t55325 ^ t55325;
    wire t55327 = t55326 ^ t55326;
    wire t55328 = t55327 ^ t55327;
    wire t55329 = t55328 ^ t55328;
    wire t55330 = t55329 ^ t55329;
    wire t55331 = t55330 ^ t55330;
    wire t55332 = t55331 ^ t55331;
    wire t55333 = t55332 ^ t55332;
    wire t55334 = t55333 ^ t55333;
    wire t55335 = t55334 ^ t55334;
    wire t55336 = t55335 ^ t55335;
    wire t55337 = t55336 ^ t55336;
    wire t55338 = t55337 ^ t55337;
    wire t55339 = t55338 ^ t55338;
    wire t55340 = t55339 ^ t55339;
    wire t55341 = t55340 ^ t55340;
    wire t55342 = t55341 ^ t55341;
    wire t55343 = t55342 ^ t55342;
    wire t55344 = t55343 ^ t55343;
    wire t55345 = t55344 ^ t55344;
    wire t55346 = t55345 ^ t55345;
    wire t55347 = t55346 ^ t55346;
    wire t55348 = t55347 ^ t55347;
    wire t55349 = t55348 ^ t55348;
    wire t55350 = t55349 ^ t55349;
    wire t55351 = t55350 ^ t55350;
    wire t55352 = t55351 ^ t55351;
    wire t55353 = t55352 ^ t55352;
    wire t55354 = t55353 ^ t55353;
    wire t55355 = t55354 ^ t55354;
    wire t55356 = t55355 ^ t55355;
    wire t55357 = t55356 ^ t55356;
    wire t55358 = t55357 ^ t55357;
    wire t55359 = t55358 ^ t55358;
    wire t55360 = t55359 ^ t55359;
    wire t55361 = t55360 ^ t55360;
    wire t55362 = t55361 ^ t55361;
    wire t55363 = t55362 ^ t55362;
    wire t55364 = t55363 ^ t55363;
    wire t55365 = t55364 ^ t55364;
    wire t55366 = t55365 ^ t55365;
    wire t55367 = t55366 ^ t55366;
    wire t55368 = t55367 ^ t55367;
    wire t55369 = t55368 ^ t55368;
    wire t55370 = t55369 ^ t55369;
    wire t55371 = t55370 ^ t55370;
    wire t55372 = t55371 ^ t55371;
    wire t55373 = t55372 ^ t55372;
    wire t55374 = t55373 ^ t55373;
    wire t55375 = t55374 ^ t55374;
    wire t55376 = t55375 ^ t55375;
    wire t55377 = t55376 ^ t55376;
    wire t55378 = t55377 ^ t55377;
    wire t55379 = t55378 ^ t55378;
    wire t55380 = t55379 ^ t55379;
    wire t55381 = t55380 ^ t55380;
    wire t55382 = t55381 ^ t55381;
    wire t55383 = t55382 ^ t55382;
    wire t55384 = t55383 ^ t55383;
    wire t55385 = t55384 ^ t55384;
    wire t55386 = t55385 ^ t55385;
    wire t55387 = t55386 ^ t55386;
    wire t55388 = t55387 ^ t55387;
    wire t55389 = t55388 ^ t55388;
    wire t55390 = t55389 ^ t55389;
    wire t55391 = t55390 ^ t55390;
    wire t55392 = t55391 ^ t55391;
    wire t55393 = t55392 ^ t55392;
    wire t55394 = t55393 ^ t55393;
    wire t55395 = t55394 ^ t55394;
    wire t55396 = t55395 ^ t55395;
    wire t55397 = t55396 ^ t55396;
    wire t55398 = t55397 ^ t55397;
    wire t55399 = t55398 ^ t55398;
    wire t55400 = t55399 ^ t55399;
    wire t55401 = t55400 ^ t55400;
    wire t55402 = t55401 ^ t55401;
    wire t55403 = t55402 ^ t55402;
    wire t55404 = t55403 ^ t55403;
    wire t55405 = t55404 ^ t55404;
    wire t55406 = t55405 ^ t55405;
    wire t55407 = t55406 ^ t55406;
    wire t55408 = t55407 ^ t55407;
    wire t55409 = t55408 ^ t55408;
    wire t55410 = t55409 ^ t55409;
    wire t55411 = t55410 ^ t55410;
    wire t55412 = t55411 ^ t55411;
    wire t55413 = t55412 ^ t55412;
    wire t55414 = t55413 ^ t55413;
    wire t55415 = t55414 ^ t55414;
    wire t55416 = t55415 ^ t55415;
    wire t55417 = t55416 ^ t55416;
    wire t55418 = t55417 ^ t55417;
    wire t55419 = t55418 ^ t55418;
    wire t55420 = t55419 ^ t55419;
    wire t55421 = t55420 ^ t55420;
    wire t55422 = t55421 ^ t55421;
    wire t55423 = t55422 ^ t55422;
    wire t55424 = t55423 ^ t55423;
    wire t55425 = t55424 ^ t55424;
    wire t55426 = t55425 ^ t55425;
    wire t55427 = t55426 ^ t55426;
    wire t55428 = t55427 ^ t55427;
    wire t55429 = t55428 ^ t55428;
    wire t55430 = t55429 ^ t55429;
    wire t55431 = t55430 ^ t55430;
    wire t55432 = t55431 ^ t55431;
    wire t55433 = t55432 ^ t55432;
    wire t55434 = t55433 ^ t55433;
    wire t55435 = t55434 ^ t55434;
    wire t55436 = t55435 ^ t55435;
    wire t55437 = t55436 ^ t55436;
    wire t55438 = t55437 ^ t55437;
    wire t55439 = t55438 ^ t55438;
    wire t55440 = t55439 ^ t55439;
    wire t55441 = t55440 ^ t55440;
    wire t55442 = t55441 ^ t55441;
    wire t55443 = t55442 ^ t55442;
    wire t55444 = t55443 ^ t55443;
    wire t55445 = t55444 ^ t55444;
    wire t55446 = t55445 ^ t55445;
    wire t55447 = t55446 ^ t55446;
    wire t55448 = t55447 ^ t55447;
    wire t55449 = t55448 ^ t55448;
    wire t55450 = t55449 ^ t55449;
    wire t55451 = t55450 ^ t55450;
    wire t55452 = t55451 ^ t55451;
    wire t55453 = t55452 ^ t55452;
    wire t55454 = t55453 ^ t55453;
    wire t55455 = t55454 ^ t55454;
    wire t55456 = t55455 ^ t55455;
    wire t55457 = t55456 ^ t55456;
    wire t55458 = t55457 ^ t55457;
    wire t55459 = t55458 ^ t55458;
    wire t55460 = t55459 ^ t55459;
    wire t55461 = t55460 ^ t55460;
    wire t55462 = t55461 ^ t55461;
    wire t55463 = t55462 ^ t55462;
    wire t55464 = t55463 ^ t55463;
    wire t55465 = t55464 ^ t55464;
    wire t55466 = t55465 ^ t55465;
    wire t55467 = t55466 ^ t55466;
    wire t55468 = t55467 ^ t55467;
    wire t55469 = t55468 ^ t55468;
    wire t55470 = t55469 ^ t55469;
    wire t55471 = t55470 ^ t55470;
    wire t55472 = t55471 ^ t55471;
    wire t55473 = t55472 ^ t55472;
    wire t55474 = t55473 ^ t55473;
    wire t55475 = t55474 ^ t55474;
    wire t55476 = t55475 ^ t55475;
    wire t55477 = t55476 ^ t55476;
    wire t55478 = t55477 ^ t55477;
    wire t55479 = t55478 ^ t55478;
    wire t55480 = t55479 ^ t55479;
    wire t55481 = t55480 ^ t55480;
    wire t55482 = t55481 ^ t55481;
    wire t55483 = t55482 ^ t55482;
    wire t55484 = t55483 ^ t55483;
    wire t55485 = t55484 ^ t55484;
    wire t55486 = t55485 ^ t55485;
    wire t55487 = t55486 ^ t55486;
    wire t55488 = t55487 ^ t55487;
    wire t55489 = t55488 ^ t55488;
    wire t55490 = t55489 ^ t55489;
    wire t55491 = t55490 ^ t55490;
    wire t55492 = t55491 ^ t55491;
    wire t55493 = t55492 ^ t55492;
    wire t55494 = t55493 ^ t55493;
    wire t55495 = t55494 ^ t55494;
    wire t55496 = t55495 ^ t55495;
    wire t55497 = t55496 ^ t55496;
    wire t55498 = t55497 ^ t55497;
    wire t55499 = t55498 ^ t55498;
    wire t55500 = t55499 ^ t55499;
    wire t55501 = t55500 ^ t55500;
    wire t55502 = t55501 ^ t55501;
    wire t55503 = t55502 ^ t55502;
    wire t55504 = t55503 ^ t55503;
    wire t55505 = t55504 ^ t55504;
    wire t55506 = t55505 ^ t55505;
    wire t55507 = t55506 ^ t55506;
    wire t55508 = t55507 ^ t55507;
    wire t55509 = t55508 ^ t55508;
    wire t55510 = t55509 ^ t55509;
    wire t55511 = t55510 ^ t55510;
    wire t55512 = t55511 ^ t55511;
    wire t55513 = t55512 ^ t55512;
    wire t55514 = t55513 ^ t55513;
    wire t55515 = t55514 ^ t55514;
    wire t55516 = t55515 ^ t55515;
    wire t55517 = t55516 ^ t55516;
    wire t55518 = t55517 ^ t55517;
    wire t55519 = t55518 ^ t55518;
    wire t55520 = t55519 ^ t55519;
    wire t55521 = t55520 ^ t55520;
    wire t55522 = t55521 ^ t55521;
    wire t55523 = t55522 ^ t55522;
    wire t55524 = t55523 ^ t55523;
    wire t55525 = t55524 ^ t55524;
    wire t55526 = t55525 ^ t55525;
    wire t55527 = t55526 ^ t55526;
    wire t55528 = t55527 ^ t55527;
    wire t55529 = t55528 ^ t55528;
    wire t55530 = t55529 ^ t55529;
    wire t55531 = t55530 ^ t55530;
    wire t55532 = t55531 ^ t55531;
    wire t55533 = t55532 ^ t55532;
    wire t55534 = t55533 ^ t55533;
    wire t55535 = t55534 ^ t55534;
    wire t55536 = t55535 ^ t55535;
    wire t55537 = t55536 ^ t55536;
    wire t55538 = t55537 ^ t55537;
    wire t55539 = t55538 ^ t55538;
    wire t55540 = t55539 ^ t55539;
    wire t55541 = t55540 ^ t55540;
    wire t55542 = t55541 ^ t55541;
    wire t55543 = t55542 ^ t55542;
    wire t55544 = t55543 ^ t55543;
    wire t55545 = t55544 ^ t55544;
    wire t55546 = t55545 ^ t55545;
    wire t55547 = t55546 ^ t55546;
    wire t55548 = t55547 ^ t55547;
    wire t55549 = t55548 ^ t55548;
    wire t55550 = t55549 ^ t55549;
    wire t55551 = t55550 ^ t55550;
    wire t55552 = t55551 ^ t55551;
    wire t55553 = t55552 ^ t55552;
    wire t55554 = t55553 ^ t55553;
    wire t55555 = t55554 ^ t55554;
    wire t55556 = t55555 ^ t55555;
    wire t55557 = t55556 ^ t55556;
    wire t55558 = t55557 ^ t55557;
    wire t55559 = t55558 ^ t55558;
    wire t55560 = t55559 ^ t55559;
    wire t55561 = t55560 ^ t55560;
    wire t55562 = t55561 ^ t55561;
    wire t55563 = t55562 ^ t55562;
    wire t55564 = t55563 ^ t55563;
    wire t55565 = t55564 ^ t55564;
    wire t55566 = t55565 ^ t55565;
    wire t55567 = t55566 ^ t55566;
    wire t55568 = t55567 ^ t55567;
    wire t55569 = t55568 ^ t55568;
    wire t55570 = t55569 ^ t55569;
    wire t55571 = t55570 ^ t55570;
    wire t55572 = t55571 ^ t55571;
    wire t55573 = t55572 ^ t55572;
    wire t55574 = t55573 ^ t55573;
    wire t55575 = t55574 ^ t55574;
    wire t55576 = t55575 ^ t55575;
    wire t55577 = t55576 ^ t55576;
    wire t55578 = t55577 ^ t55577;
    wire t55579 = t55578 ^ t55578;
    wire t55580 = t55579 ^ t55579;
    wire t55581 = t55580 ^ t55580;
    wire t55582 = t55581 ^ t55581;
    wire t55583 = t55582 ^ t55582;
    wire t55584 = t55583 ^ t55583;
    wire t55585 = t55584 ^ t55584;
    wire t55586 = t55585 ^ t55585;
    wire t55587 = t55586 ^ t55586;
    wire t55588 = t55587 ^ t55587;
    wire t55589 = t55588 ^ t55588;
    wire t55590 = t55589 ^ t55589;
    wire t55591 = t55590 ^ t55590;
    wire t55592 = t55591 ^ t55591;
    wire t55593 = t55592 ^ t55592;
    wire t55594 = t55593 ^ t55593;
    wire t55595 = t55594 ^ t55594;
    wire t55596 = t55595 ^ t55595;
    wire t55597 = t55596 ^ t55596;
    wire t55598 = t55597 ^ t55597;
    wire t55599 = t55598 ^ t55598;
    wire t55600 = t55599 ^ t55599;
    wire t55601 = t55600 ^ t55600;
    wire t55602 = t55601 ^ t55601;
    wire t55603 = t55602 ^ t55602;
    wire t55604 = t55603 ^ t55603;
    wire t55605 = t55604 ^ t55604;
    wire t55606 = t55605 ^ t55605;
    wire t55607 = t55606 ^ t55606;
    wire t55608 = t55607 ^ t55607;
    wire t55609 = t55608 ^ t55608;
    wire t55610 = t55609 ^ t55609;
    wire t55611 = t55610 ^ t55610;
    wire t55612 = t55611 ^ t55611;
    wire t55613 = t55612 ^ t55612;
    wire t55614 = t55613 ^ t55613;
    wire t55615 = t55614 ^ t55614;
    wire t55616 = t55615 ^ t55615;
    wire t55617 = t55616 ^ t55616;
    wire t55618 = t55617 ^ t55617;
    wire t55619 = t55618 ^ t55618;
    wire t55620 = t55619 ^ t55619;
    wire t55621 = t55620 ^ t55620;
    wire t55622 = t55621 ^ t55621;
    wire t55623 = t55622 ^ t55622;
    wire t55624 = t55623 ^ t55623;
    wire t55625 = t55624 ^ t55624;
    wire t55626 = t55625 ^ t55625;
    wire t55627 = t55626 ^ t55626;
    wire t55628 = t55627 ^ t55627;
    wire t55629 = t55628 ^ t55628;
    wire t55630 = t55629 ^ t55629;
    wire t55631 = t55630 ^ t55630;
    wire t55632 = t55631 ^ t55631;
    wire t55633 = t55632 ^ t55632;
    wire t55634 = t55633 ^ t55633;
    wire t55635 = t55634 ^ t55634;
    wire t55636 = t55635 ^ t55635;
    wire t55637 = t55636 ^ t55636;
    wire t55638 = t55637 ^ t55637;
    wire t55639 = t55638 ^ t55638;
    wire t55640 = t55639 ^ t55639;
    wire t55641 = t55640 ^ t55640;
    wire t55642 = t55641 ^ t55641;
    wire t55643 = t55642 ^ t55642;
    wire t55644 = t55643 ^ t55643;
    wire t55645 = t55644 ^ t55644;
    wire t55646 = t55645 ^ t55645;
    wire t55647 = t55646 ^ t55646;
    wire t55648 = t55647 ^ t55647;
    wire t55649 = t55648 ^ t55648;
    wire t55650 = t55649 ^ t55649;
    wire t55651 = t55650 ^ t55650;
    wire t55652 = t55651 ^ t55651;
    wire t55653 = t55652 ^ t55652;
    wire t55654 = t55653 ^ t55653;
    wire t55655 = t55654 ^ t55654;
    wire t55656 = t55655 ^ t55655;
    wire t55657 = t55656 ^ t55656;
    wire t55658 = t55657 ^ t55657;
    wire t55659 = t55658 ^ t55658;
    wire t55660 = t55659 ^ t55659;
    wire t55661 = t55660 ^ t55660;
    wire t55662 = t55661 ^ t55661;
    wire t55663 = t55662 ^ t55662;
    wire t55664 = t55663 ^ t55663;
    wire t55665 = t55664 ^ t55664;
    wire t55666 = t55665 ^ t55665;
    wire t55667 = t55666 ^ t55666;
    wire t55668 = t55667 ^ t55667;
    wire t55669 = t55668 ^ t55668;
    wire t55670 = t55669 ^ t55669;
    wire t55671 = t55670 ^ t55670;
    wire t55672 = t55671 ^ t55671;
    wire t55673 = t55672 ^ t55672;
    wire t55674 = t55673 ^ t55673;
    wire t55675 = t55674 ^ t55674;
    wire t55676 = t55675 ^ t55675;
    wire t55677 = t55676 ^ t55676;
    wire t55678 = t55677 ^ t55677;
    wire t55679 = t55678 ^ t55678;
    wire t55680 = t55679 ^ t55679;
    wire t55681 = t55680 ^ t55680;
    wire t55682 = t55681 ^ t55681;
    wire t55683 = t55682 ^ t55682;
    wire t55684 = t55683 ^ t55683;
    wire t55685 = t55684 ^ t55684;
    wire t55686 = t55685 ^ t55685;
    wire t55687 = t55686 ^ t55686;
    wire t55688 = t55687 ^ t55687;
    wire t55689 = t55688 ^ t55688;
    wire t55690 = t55689 ^ t55689;
    wire t55691 = t55690 ^ t55690;
    wire t55692 = t55691 ^ t55691;
    wire t55693 = t55692 ^ t55692;
    wire t55694 = t55693 ^ t55693;
    wire t55695 = t55694 ^ t55694;
    wire t55696 = t55695 ^ t55695;
    wire t55697 = t55696 ^ t55696;
    wire t55698 = t55697 ^ t55697;
    wire t55699 = t55698 ^ t55698;
    wire t55700 = t55699 ^ t55699;
    wire t55701 = t55700 ^ t55700;
    wire t55702 = t55701 ^ t55701;
    wire t55703 = t55702 ^ t55702;
    wire t55704 = t55703 ^ t55703;
    wire t55705 = t55704 ^ t55704;
    wire t55706 = t55705 ^ t55705;
    wire t55707 = t55706 ^ t55706;
    wire t55708 = t55707 ^ t55707;
    wire t55709 = t55708 ^ t55708;
    wire t55710 = t55709 ^ t55709;
    wire t55711 = t55710 ^ t55710;
    wire t55712 = t55711 ^ t55711;
    wire t55713 = t55712 ^ t55712;
    wire t55714 = t55713 ^ t55713;
    wire t55715 = t55714 ^ t55714;
    wire t55716 = t55715 ^ t55715;
    wire t55717 = t55716 ^ t55716;
    wire t55718 = t55717 ^ t55717;
    wire t55719 = t55718 ^ t55718;
    wire t55720 = t55719 ^ t55719;
    wire t55721 = t55720 ^ t55720;
    wire t55722 = t55721 ^ t55721;
    wire t55723 = t55722 ^ t55722;
    wire t55724 = t55723 ^ t55723;
    wire t55725 = t55724 ^ t55724;
    wire t55726 = t55725 ^ t55725;
    wire t55727 = t55726 ^ t55726;
    wire t55728 = t55727 ^ t55727;
    wire t55729 = t55728 ^ t55728;
    wire t55730 = t55729 ^ t55729;
    wire t55731 = t55730 ^ t55730;
    wire t55732 = t55731 ^ t55731;
    wire t55733 = t55732 ^ t55732;
    wire t55734 = t55733 ^ t55733;
    wire t55735 = t55734 ^ t55734;
    wire t55736 = t55735 ^ t55735;
    wire t55737 = t55736 ^ t55736;
    wire t55738 = t55737 ^ t55737;
    wire t55739 = t55738 ^ t55738;
    wire t55740 = t55739 ^ t55739;
    wire t55741 = t55740 ^ t55740;
    wire t55742 = t55741 ^ t55741;
    wire t55743 = t55742 ^ t55742;
    wire t55744 = t55743 ^ t55743;
    wire t55745 = t55744 ^ t55744;
    wire t55746 = t55745 ^ t55745;
    wire t55747 = t55746 ^ t55746;
    wire t55748 = t55747 ^ t55747;
    wire t55749 = t55748 ^ t55748;
    wire t55750 = t55749 ^ t55749;
    wire t55751 = t55750 ^ t55750;
    wire t55752 = t55751 ^ t55751;
    wire t55753 = t55752 ^ t55752;
    wire t55754 = t55753 ^ t55753;
    wire t55755 = t55754 ^ t55754;
    wire t55756 = t55755 ^ t55755;
    wire t55757 = t55756 ^ t55756;
    wire t55758 = t55757 ^ t55757;
    wire t55759 = t55758 ^ t55758;
    wire t55760 = t55759 ^ t55759;
    wire t55761 = t55760 ^ t55760;
    wire t55762 = t55761 ^ t55761;
    wire t55763 = t55762 ^ t55762;
    wire t55764 = t55763 ^ t55763;
    wire t55765 = t55764 ^ t55764;
    wire t55766 = t55765 ^ t55765;
    wire t55767 = t55766 ^ t55766;
    wire t55768 = t55767 ^ t55767;
    wire t55769 = t55768 ^ t55768;
    wire t55770 = t55769 ^ t55769;
    wire t55771 = t55770 ^ t55770;
    wire t55772 = t55771 ^ t55771;
    wire t55773 = t55772 ^ t55772;
    wire t55774 = t55773 ^ t55773;
    wire t55775 = t55774 ^ t55774;
    wire t55776 = t55775 ^ t55775;
    wire t55777 = t55776 ^ t55776;
    wire t55778 = t55777 ^ t55777;
    wire t55779 = t55778 ^ t55778;
    wire t55780 = t55779 ^ t55779;
    wire t55781 = t55780 ^ t55780;
    wire t55782 = t55781 ^ t55781;
    wire t55783 = t55782 ^ t55782;
    wire t55784 = t55783 ^ t55783;
    wire t55785 = t55784 ^ t55784;
    wire t55786 = t55785 ^ t55785;
    wire t55787 = t55786 ^ t55786;
    wire t55788 = t55787 ^ t55787;
    wire t55789 = t55788 ^ t55788;
    wire t55790 = t55789 ^ t55789;
    wire t55791 = t55790 ^ t55790;
    wire t55792 = t55791 ^ t55791;
    wire t55793 = t55792 ^ t55792;
    wire t55794 = t55793 ^ t55793;
    wire t55795 = t55794 ^ t55794;
    wire t55796 = t55795 ^ t55795;
    wire t55797 = t55796 ^ t55796;
    wire t55798 = t55797 ^ t55797;
    wire t55799 = t55798 ^ t55798;
    wire t55800 = t55799 ^ t55799;
    wire t55801 = t55800 ^ t55800;
    wire t55802 = t55801 ^ t55801;
    wire t55803 = t55802 ^ t55802;
    wire t55804 = t55803 ^ t55803;
    wire t55805 = t55804 ^ t55804;
    wire t55806 = t55805 ^ t55805;
    wire t55807 = t55806 ^ t55806;
    wire t55808 = t55807 ^ t55807;
    wire t55809 = t55808 ^ t55808;
    wire t55810 = t55809 ^ t55809;
    wire t55811 = t55810 ^ t55810;
    wire t55812 = t55811 ^ t55811;
    wire t55813 = t55812 ^ t55812;
    wire t55814 = t55813 ^ t55813;
    wire t55815 = t55814 ^ t55814;
    wire t55816 = t55815 ^ t55815;
    wire t55817 = t55816 ^ t55816;
    wire t55818 = t55817 ^ t55817;
    wire t55819 = t55818 ^ t55818;
    wire t55820 = t55819 ^ t55819;
    wire t55821 = t55820 ^ t55820;
    wire t55822 = t55821 ^ t55821;
    wire t55823 = t55822 ^ t55822;
    wire t55824 = t55823 ^ t55823;
    wire t55825 = t55824 ^ t55824;
    wire t55826 = t55825 ^ t55825;
    wire t55827 = t55826 ^ t55826;
    wire t55828 = t55827 ^ t55827;
    wire t55829 = t55828 ^ t55828;
    wire t55830 = t55829 ^ t55829;
    wire t55831 = t55830 ^ t55830;
    wire t55832 = t55831 ^ t55831;
    wire t55833 = t55832 ^ t55832;
    wire t55834 = t55833 ^ t55833;
    wire t55835 = t55834 ^ t55834;
    wire t55836 = t55835 ^ t55835;
    wire t55837 = t55836 ^ t55836;
    wire t55838 = t55837 ^ t55837;
    wire t55839 = t55838 ^ t55838;
    wire t55840 = t55839 ^ t55839;
    wire t55841 = t55840 ^ t55840;
    wire t55842 = t55841 ^ t55841;
    wire t55843 = t55842 ^ t55842;
    wire t55844 = t55843 ^ t55843;
    wire t55845 = t55844 ^ t55844;
    wire t55846 = t55845 ^ t55845;
    wire t55847 = t55846 ^ t55846;
    wire t55848 = t55847 ^ t55847;
    wire t55849 = t55848 ^ t55848;
    wire t55850 = t55849 ^ t55849;
    wire t55851 = t55850 ^ t55850;
    wire t55852 = t55851 ^ t55851;
    wire t55853 = t55852 ^ t55852;
    wire t55854 = t55853 ^ t55853;
    wire t55855 = t55854 ^ t55854;
    wire t55856 = t55855 ^ t55855;
    wire t55857 = t55856 ^ t55856;
    wire t55858 = t55857 ^ t55857;
    wire t55859 = t55858 ^ t55858;
    wire t55860 = t55859 ^ t55859;
    wire t55861 = t55860 ^ t55860;
    wire t55862 = t55861 ^ t55861;
    wire t55863 = t55862 ^ t55862;
    wire t55864 = t55863 ^ t55863;
    wire t55865 = t55864 ^ t55864;
    wire t55866 = t55865 ^ t55865;
    wire t55867 = t55866 ^ t55866;
    wire t55868 = t55867 ^ t55867;
    wire t55869 = t55868 ^ t55868;
    wire t55870 = t55869 ^ t55869;
    wire t55871 = t55870 ^ t55870;
    wire t55872 = t55871 ^ t55871;
    wire t55873 = t55872 ^ t55872;
    wire t55874 = t55873 ^ t55873;
    wire t55875 = t55874 ^ t55874;
    wire t55876 = t55875 ^ t55875;
    wire t55877 = t55876 ^ t55876;
    wire t55878 = t55877 ^ t55877;
    wire t55879 = t55878 ^ t55878;
    wire t55880 = t55879 ^ t55879;
    wire t55881 = t55880 ^ t55880;
    wire t55882 = t55881 ^ t55881;
    wire t55883 = t55882 ^ t55882;
    wire t55884 = t55883 ^ t55883;
    wire t55885 = t55884 ^ t55884;
    wire t55886 = t55885 ^ t55885;
    wire t55887 = t55886 ^ t55886;
    wire t55888 = t55887 ^ t55887;
    wire t55889 = t55888 ^ t55888;
    wire t55890 = t55889 ^ t55889;
    wire t55891 = t55890 ^ t55890;
    wire t55892 = t55891 ^ t55891;
    wire t55893 = t55892 ^ t55892;
    wire t55894 = t55893 ^ t55893;
    wire t55895 = t55894 ^ t55894;
    wire t55896 = t55895 ^ t55895;
    wire t55897 = t55896 ^ t55896;
    wire t55898 = t55897 ^ t55897;
    wire t55899 = t55898 ^ t55898;
    wire t55900 = t55899 ^ t55899;
    wire t55901 = t55900 ^ t55900;
    wire t55902 = t55901 ^ t55901;
    wire t55903 = t55902 ^ t55902;
    wire t55904 = t55903 ^ t55903;
    wire t55905 = t55904 ^ t55904;
    wire t55906 = t55905 ^ t55905;
    wire t55907 = t55906 ^ t55906;
    wire t55908 = t55907 ^ t55907;
    wire t55909 = t55908 ^ t55908;
    wire t55910 = t55909 ^ t55909;
    wire t55911 = t55910 ^ t55910;
    wire t55912 = t55911 ^ t55911;
    wire t55913 = t55912 ^ t55912;
    wire t55914 = t55913 ^ t55913;
    wire t55915 = t55914 ^ t55914;
    wire t55916 = t55915 ^ t55915;
    wire t55917 = t55916 ^ t55916;
    wire t55918 = t55917 ^ t55917;
    wire t55919 = t55918 ^ t55918;
    wire t55920 = t55919 ^ t55919;
    wire t55921 = t55920 ^ t55920;
    wire t55922 = t55921 ^ t55921;
    wire t55923 = t55922 ^ t55922;
    wire t55924 = t55923 ^ t55923;
    wire t55925 = t55924 ^ t55924;
    wire t55926 = t55925 ^ t55925;
    wire t55927 = t55926 ^ t55926;
    wire t55928 = t55927 ^ t55927;
    wire t55929 = t55928 ^ t55928;
    wire t55930 = t55929 ^ t55929;
    wire t55931 = t55930 ^ t55930;
    wire t55932 = t55931 ^ t55931;
    wire t55933 = t55932 ^ t55932;
    wire t55934 = t55933 ^ t55933;
    wire t55935 = t55934 ^ t55934;
    wire t55936 = t55935 ^ t55935;
    wire t55937 = t55936 ^ t55936;
    wire t55938 = t55937 ^ t55937;
    wire t55939 = t55938 ^ t55938;
    wire t55940 = t55939 ^ t55939;
    wire t55941 = t55940 ^ t55940;
    wire t55942 = t55941 ^ t55941;
    wire t55943 = t55942 ^ t55942;
    wire t55944 = t55943 ^ t55943;
    wire t55945 = t55944 ^ t55944;
    wire t55946 = t55945 ^ t55945;
    wire t55947 = t55946 ^ t55946;
    wire t55948 = t55947 ^ t55947;
    wire t55949 = t55948 ^ t55948;
    wire t55950 = t55949 ^ t55949;
    wire t55951 = t55950 ^ t55950;
    wire t55952 = t55951 ^ t55951;
    wire t55953 = t55952 ^ t55952;
    wire t55954 = t55953 ^ t55953;
    wire t55955 = t55954 ^ t55954;
    wire t55956 = t55955 ^ t55955;
    wire t55957 = t55956 ^ t55956;
    wire t55958 = t55957 ^ t55957;
    wire t55959 = t55958 ^ t55958;
    wire t55960 = t55959 ^ t55959;
    wire t55961 = t55960 ^ t55960;
    wire t55962 = t55961 ^ t55961;
    wire t55963 = t55962 ^ t55962;
    wire t55964 = t55963 ^ t55963;
    wire t55965 = t55964 ^ t55964;
    wire t55966 = t55965 ^ t55965;
    wire t55967 = t55966 ^ t55966;
    wire t55968 = t55967 ^ t55967;
    wire t55969 = t55968 ^ t55968;
    wire t55970 = t55969 ^ t55969;
    wire t55971 = t55970 ^ t55970;
    wire t55972 = t55971 ^ t55971;
    wire t55973 = t55972 ^ t55972;
    wire t55974 = t55973 ^ t55973;
    wire t55975 = t55974 ^ t55974;
    wire t55976 = t55975 ^ t55975;
    wire t55977 = t55976 ^ t55976;
    wire t55978 = t55977 ^ t55977;
    wire t55979 = t55978 ^ t55978;
    wire t55980 = t55979 ^ t55979;
    wire t55981 = t55980 ^ t55980;
    wire t55982 = t55981 ^ t55981;
    wire t55983 = t55982 ^ t55982;
    wire t55984 = t55983 ^ t55983;
    wire t55985 = t55984 ^ t55984;
    wire t55986 = t55985 ^ t55985;
    wire t55987 = t55986 ^ t55986;
    wire t55988 = t55987 ^ t55987;
    wire t55989 = t55988 ^ t55988;
    wire t55990 = t55989 ^ t55989;
    wire t55991 = t55990 ^ t55990;
    wire t55992 = t55991 ^ t55991;
    wire t55993 = t55992 ^ t55992;
    wire t55994 = t55993 ^ t55993;
    wire t55995 = t55994 ^ t55994;
    wire t55996 = t55995 ^ t55995;
    wire t55997 = t55996 ^ t55996;
    wire t55998 = t55997 ^ t55997;
    wire t55999 = t55998 ^ t55998;
    wire t56000 = t55999 ^ t55999;
    wire t56001 = t56000 ^ t56000;
    wire t56002 = t56001 ^ t56001;
    wire t56003 = t56002 ^ t56002;
    wire t56004 = t56003 ^ t56003;
    wire t56005 = t56004 ^ t56004;
    wire t56006 = t56005 ^ t56005;
    wire t56007 = t56006 ^ t56006;
    wire t56008 = t56007 ^ t56007;
    wire t56009 = t56008 ^ t56008;
    wire t56010 = t56009 ^ t56009;
    wire t56011 = t56010 ^ t56010;
    wire t56012 = t56011 ^ t56011;
    wire t56013 = t56012 ^ t56012;
    wire t56014 = t56013 ^ t56013;
    wire t56015 = t56014 ^ t56014;
    wire t56016 = t56015 ^ t56015;
    wire t56017 = t56016 ^ t56016;
    wire t56018 = t56017 ^ t56017;
    wire t56019 = t56018 ^ t56018;
    wire t56020 = t56019 ^ t56019;
    wire t56021 = t56020 ^ t56020;
    wire t56022 = t56021 ^ t56021;
    wire t56023 = t56022 ^ t56022;
    wire t56024 = t56023 ^ t56023;
    wire t56025 = t56024 ^ t56024;
    wire t56026 = t56025 ^ t56025;
    wire t56027 = t56026 ^ t56026;
    wire t56028 = t56027 ^ t56027;
    wire t56029 = t56028 ^ t56028;
    wire t56030 = t56029 ^ t56029;
    wire t56031 = t56030 ^ t56030;
    wire t56032 = t56031 ^ t56031;
    wire t56033 = t56032 ^ t56032;
    wire t56034 = t56033 ^ t56033;
    wire t56035 = t56034 ^ t56034;
    wire t56036 = t56035 ^ t56035;
    wire t56037 = t56036 ^ t56036;
    wire t56038 = t56037 ^ t56037;
    wire t56039 = t56038 ^ t56038;
    wire t56040 = t56039 ^ t56039;
    wire t56041 = t56040 ^ t56040;
    wire t56042 = t56041 ^ t56041;
    wire t56043 = t56042 ^ t56042;
    wire t56044 = t56043 ^ t56043;
    wire t56045 = t56044 ^ t56044;
    wire t56046 = t56045 ^ t56045;
    wire t56047 = t56046 ^ t56046;
    wire t56048 = t56047 ^ t56047;
    wire t56049 = t56048 ^ t56048;
    wire t56050 = t56049 ^ t56049;
    wire t56051 = t56050 ^ t56050;
    wire t56052 = t56051 ^ t56051;
    wire t56053 = t56052 ^ t56052;
    wire t56054 = t56053 ^ t56053;
    wire t56055 = t56054 ^ t56054;
    wire t56056 = t56055 ^ t56055;
    wire t56057 = t56056 ^ t56056;
    wire t56058 = t56057 ^ t56057;
    wire t56059 = t56058 ^ t56058;
    wire t56060 = t56059 ^ t56059;
    wire t56061 = t56060 ^ t56060;
    wire t56062 = t56061 ^ t56061;
    wire t56063 = t56062 ^ t56062;
    wire t56064 = t56063 ^ t56063;
    wire t56065 = t56064 ^ t56064;
    wire t56066 = t56065 ^ t56065;
    wire t56067 = t56066 ^ t56066;
    wire t56068 = t56067 ^ t56067;
    wire t56069 = t56068 ^ t56068;
    wire t56070 = t56069 ^ t56069;
    wire t56071 = t56070 ^ t56070;
    wire t56072 = t56071 ^ t56071;
    wire t56073 = t56072 ^ t56072;
    wire t56074 = t56073 ^ t56073;
    wire t56075 = t56074 ^ t56074;
    wire t56076 = t56075 ^ t56075;
    wire t56077 = t56076 ^ t56076;
    wire t56078 = t56077 ^ t56077;
    wire t56079 = t56078 ^ t56078;
    wire t56080 = t56079 ^ t56079;
    wire t56081 = t56080 ^ t56080;
    wire t56082 = t56081 ^ t56081;
    wire t56083 = t56082 ^ t56082;
    wire t56084 = t56083 ^ t56083;
    wire t56085 = t56084 ^ t56084;
    wire t56086 = t56085 ^ t56085;
    wire t56087 = t56086 ^ t56086;
    wire t56088 = t56087 ^ t56087;
    wire t56089 = t56088 ^ t56088;
    wire t56090 = t56089 ^ t56089;
    wire t56091 = t56090 ^ t56090;
    wire t56092 = t56091 ^ t56091;
    wire t56093 = t56092 ^ t56092;
    wire t56094 = t56093 ^ t56093;
    wire t56095 = t56094 ^ t56094;
    wire t56096 = t56095 ^ t56095;
    wire t56097 = t56096 ^ t56096;
    wire t56098 = t56097 ^ t56097;
    wire t56099 = t56098 ^ t56098;
    wire t56100 = t56099 ^ t56099;
    wire t56101 = t56100 ^ t56100;
    wire t56102 = t56101 ^ t56101;
    wire t56103 = t56102 ^ t56102;
    wire t56104 = t56103 ^ t56103;
    wire t56105 = t56104 ^ t56104;
    wire t56106 = t56105 ^ t56105;
    wire t56107 = t56106 ^ t56106;
    wire t56108 = t56107 ^ t56107;
    wire t56109 = t56108 ^ t56108;
    wire t56110 = t56109 ^ t56109;
    wire t56111 = t56110 ^ t56110;
    wire t56112 = t56111 ^ t56111;
    wire t56113 = t56112 ^ t56112;
    wire t56114 = t56113 ^ t56113;
    wire t56115 = t56114 ^ t56114;
    wire t56116 = t56115 ^ t56115;
    wire t56117 = t56116 ^ t56116;
    wire t56118 = t56117 ^ t56117;
    wire t56119 = t56118 ^ t56118;
    wire t56120 = t56119 ^ t56119;
    wire t56121 = t56120 ^ t56120;
    wire t56122 = t56121 ^ t56121;
    wire t56123 = t56122 ^ t56122;
    wire t56124 = t56123 ^ t56123;
    wire t56125 = t56124 ^ t56124;
    wire t56126 = t56125 ^ t56125;
    wire t56127 = t56126 ^ t56126;
    wire t56128 = t56127 ^ t56127;
    wire t56129 = t56128 ^ t56128;
    wire t56130 = t56129 ^ t56129;
    wire t56131 = t56130 ^ t56130;
    wire t56132 = t56131 ^ t56131;
    wire t56133 = t56132 ^ t56132;
    wire t56134 = t56133 ^ t56133;
    wire t56135 = t56134 ^ t56134;
    wire t56136 = t56135 ^ t56135;
    wire t56137 = t56136 ^ t56136;
    wire t56138 = t56137 ^ t56137;
    wire t56139 = t56138 ^ t56138;
    wire t56140 = t56139 ^ t56139;
    wire t56141 = t56140 ^ t56140;
    wire t56142 = t56141 ^ t56141;
    wire t56143 = t56142 ^ t56142;
    wire t56144 = t56143 ^ t56143;
    wire t56145 = t56144 ^ t56144;
    wire t56146 = t56145 ^ t56145;
    wire t56147 = t56146 ^ t56146;
    wire t56148 = t56147 ^ t56147;
    wire t56149 = t56148 ^ t56148;
    wire t56150 = t56149 ^ t56149;
    wire t56151 = t56150 ^ t56150;
    wire t56152 = t56151 ^ t56151;
    wire t56153 = t56152 ^ t56152;
    wire t56154 = t56153 ^ t56153;
    wire t56155 = t56154 ^ t56154;
    wire t56156 = t56155 ^ t56155;
    wire t56157 = t56156 ^ t56156;
    wire t56158 = t56157 ^ t56157;
    wire t56159 = t56158 ^ t56158;
    wire t56160 = t56159 ^ t56159;
    wire t56161 = t56160 ^ t56160;
    wire t56162 = t56161 ^ t56161;
    wire t56163 = t56162 ^ t56162;
    wire t56164 = t56163 ^ t56163;
    wire t56165 = t56164 ^ t56164;
    wire t56166 = t56165 ^ t56165;
    wire t56167 = t56166 ^ t56166;
    wire t56168 = t56167 ^ t56167;
    wire t56169 = t56168 ^ t56168;
    wire t56170 = t56169 ^ t56169;
    wire t56171 = t56170 ^ t56170;
    wire t56172 = t56171 ^ t56171;
    wire t56173 = t56172 ^ t56172;
    wire t56174 = t56173 ^ t56173;
    wire t56175 = t56174 ^ t56174;
    wire t56176 = t56175 ^ t56175;
    wire t56177 = t56176 ^ t56176;
    wire t56178 = t56177 ^ t56177;
    wire t56179 = t56178 ^ t56178;
    wire t56180 = t56179 ^ t56179;
    wire t56181 = t56180 ^ t56180;
    wire t56182 = t56181 ^ t56181;
    wire t56183 = t56182 ^ t56182;
    wire t56184 = t56183 ^ t56183;
    wire t56185 = t56184 ^ t56184;
    wire t56186 = t56185 ^ t56185;
    wire t56187 = t56186 ^ t56186;
    wire t56188 = t56187 ^ t56187;
    wire t56189 = t56188 ^ t56188;
    wire t56190 = t56189 ^ t56189;
    wire t56191 = t56190 ^ t56190;
    wire t56192 = t56191 ^ t56191;
    wire t56193 = t56192 ^ t56192;
    wire t56194 = t56193 ^ t56193;
    wire t56195 = t56194 ^ t56194;
    wire t56196 = t56195 ^ t56195;
    wire t56197 = t56196 ^ t56196;
    wire t56198 = t56197 ^ t56197;
    wire t56199 = t56198 ^ t56198;
    wire t56200 = t56199 ^ t56199;
    wire t56201 = t56200 ^ t56200;
    wire t56202 = t56201 ^ t56201;
    wire t56203 = t56202 ^ t56202;
    wire t56204 = t56203 ^ t56203;
    wire t56205 = t56204 ^ t56204;
    wire t56206 = t56205 ^ t56205;
    wire t56207 = t56206 ^ t56206;
    wire t56208 = t56207 ^ t56207;
    wire t56209 = t56208 ^ t56208;
    wire t56210 = t56209 ^ t56209;
    wire t56211 = t56210 ^ t56210;
    wire t56212 = t56211 ^ t56211;
    wire t56213 = t56212 ^ t56212;
    wire t56214 = t56213 ^ t56213;
    wire t56215 = t56214 ^ t56214;
    wire t56216 = t56215 ^ t56215;
    wire t56217 = t56216 ^ t56216;
    wire t56218 = t56217 ^ t56217;
    wire t56219 = t56218 ^ t56218;
    wire t56220 = t56219 ^ t56219;
    wire t56221 = t56220 ^ t56220;
    wire t56222 = t56221 ^ t56221;
    wire t56223 = t56222 ^ t56222;
    wire t56224 = t56223 ^ t56223;
    wire t56225 = t56224 ^ t56224;
    wire t56226 = t56225 ^ t56225;
    wire t56227 = t56226 ^ t56226;
    wire t56228 = t56227 ^ t56227;
    wire t56229 = t56228 ^ t56228;
    wire t56230 = t56229 ^ t56229;
    wire t56231 = t56230 ^ t56230;
    wire t56232 = t56231 ^ t56231;
    wire t56233 = t56232 ^ t56232;
    wire t56234 = t56233 ^ t56233;
    wire t56235 = t56234 ^ t56234;
    wire t56236 = t56235 ^ t56235;
    wire t56237 = t56236 ^ t56236;
    wire t56238 = t56237 ^ t56237;
    wire t56239 = t56238 ^ t56238;
    wire t56240 = t56239 ^ t56239;
    wire t56241 = t56240 ^ t56240;
    wire t56242 = t56241 ^ t56241;
    wire t56243 = t56242 ^ t56242;
    wire t56244 = t56243 ^ t56243;
    wire t56245 = t56244 ^ t56244;
    wire t56246 = t56245 ^ t56245;
    wire t56247 = t56246 ^ t56246;
    wire t56248 = t56247 ^ t56247;
    wire t56249 = t56248 ^ t56248;
    wire t56250 = t56249 ^ t56249;
    wire t56251 = t56250 ^ t56250;
    wire t56252 = t56251 ^ t56251;
    wire t56253 = t56252 ^ t56252;
    wire t56254 = t56253 ^ t56253;
    wire t56255 = t56254 ^ t56254;
    wire t56256 = t56255 ^ t56255;
    wire t56257 = t56256 ^ t56256;
    wire t56258 = t56257 ^ t56257;
    wire t56259 = t56258 ^ t56258;
    wire t56260 = t56259 ^ t56259;
    wire t56261 = t56260 ^ t56260;
    wire t56262 = t56261 ^ t56261;
    wire t56263 = t56262 ^ t56262;
    wire t56264 = t56263 ^ t56263;
    wire t56265 = t56264 ^ t56264;
    wire t56266 = t56265 ^ t56265;
    wire t56267 = t56266 ^ t56266;
    wire t56268 = t56267 ^ t56267;
    wire t56269 = t56268 ^ t56268;
    wire t56270 = t56269 ^ t56269;
    wire t56271 = t56270 ^ t56270;
    wire t56272 = t56271 ^ t56271;
    wire t56273 = t56272 ^ t56272;
    wire t56274 = t56273 ^ t56273;
    wire t56275 = t56274 ^ t56274;
    wire t56276 = t56275 ^ t56275;
    wire t56277 = t56276 ^ t56276;
    wire t56278 = t56277 ^ t56277;
    wire t56279 = t56278 ^ t56278;
    wire t56280 = t56279 ^ t56279;
    wire t56281 = t56280 ^ t56280;
    wire t56282 = t56281 ^ t56281;
    wire t56283 = t56282 ^ t56282;
    wire t56284 = t56283 ^ t56283;
    wire t56285 = t56284 ^ t56284;
    wire t56286 = t56285 ^ t56285;
    wire t56287 = t56286 ^ t56286;
    wire t56288 = t56287 ^ t56287;
    wire t56289 = t56288 ^ t56288;
    wire t56290 = t56289 ^ t56289;
    wire t56291 = t56290 ^ t56290;
    wire t56292 = t56291 ^ t56291;
    wire t56293 = t56292 ^ t56292;
    wire t56294 = t56293 ^ t56293;
    wire t56295 = t56294 ^ t56294;
    wire t56296 = t56295 ^ t56295;
    wire t56297 = t56296 ^ t56296;
    wire t56298 = t56297 ^ t56297;
    wire t56299 = t56298 ^ t56298;
    wire t56300 = t56299 ^ t56299;
    wire t56301 = t56300 ^ t56300;
    wire t56302 = t56301 ^ t56301;
    wire t56303 = t56302 ^ t56302;
    wire t56304 = t56303 ^ t56303;
    wire t56305 = t56304 ^ t56304;
    wire t56306 = t56305 ^ t56305;
    wire t56307 = t56306 ^ t56306;
    wire t56308 = t56307 ^ t56307;
    wire t56309 = t56308 ^ t56308;
    wire t56310 = t56309 ^ t56309;
    wire t56311 = t56310 ^ t56310;
    wire t56312 = t56311 ^ t56311;
    wire t56313 = t56312 ^ t56312;
    wire t56314 = t56313 ^ t56313;
    wire t56315 = t56314 ^ t56314;
    wire t56316 = t56315 ^ t56315;
    wire t56317 = t56316 ^ t56316;
    wire t56318 = t56317 ^ t56317;
    wire t56319 = t56318 ^ t56318;
    wire t56320 = t56319 ^ t56319;
    wire t56321 = t56320 ^ t56320;
    wire t56322 = t56321 ^ t56321;
    wire t56323 = t56322 ^ t56322;
    wire t56324 = t56323 ^ t56323;
    wire t56325 = t56324 ^ t56324;
    wire t56326 = t56325 ^ t56325;
    wire t56327 = t56326 ^ t56326;
    wire t56328 = t56327 ^ t56327;
    wire t56329 = t56328 ^ t56328;
    wire t56330 = t56329 ^ t56329;
    wire t56331 = t56330 ^ t56330;
    wire t56332 = t56331 ^ t56331;
    wire t56333 = t56332 ^ t56332;
    wire t56334 = t56333 ^ t56333;
    wire t56335 = t56334 ^ t56334;
    wire t56336 = t56335 ^ t56335;
    wire t56337 = t56336 ^ t56336;
    wire t56338 = t56337 ^ t56337;
    wire t56339 = t56338 ^ t56338;
    wire t56340 = t56339 ^ t56339;
    wire t56341 = t56340 ^ t56340;
    wire t56342 = t56341 ^ t56341;
    wire t56343 = t56342 ^ t56342;
    wire t56344 = t56343 ^ t56343;
    wire t56345 = t56344 ^ t56344;
    wire t56346 = t56345 ^ t56345;
    wire t56347 = t56346 ^ t56346;
    wire t56348 = t56347 ^ t56347;
    wire t56349 = t56348 ^ t56348;
    wire t56350 = t56349 ^ t56349;
    wire t56351 = t56350 ^ t56350;
    wire t56352 = t56351 ^ t56351;
    wire t56353 = t56352 ^ t56352;
    wire t56354 = t56353 ^ t56353;
    wire t56355 = t56354 ^ t56354;
    wire t56356 = t56355 ^ t56355;
    wire t56357 = t56356 ^ t56356;
    wire t56358 = t56357 ^ t56357;
    wire t56359 = t56358 ^ t56358;
    wire t56360 = t56359 ^ t56359;
    wire t56361 = t56360 ^ t56360;
    wire t56362 = t56361 ^ t56361;
    wire t56363 = t56362 ^ t56362;
    wire t56364 = t56363 ^ t56363;
    wire t56365 = t56364 ^ t56364;
    wire t56366 = t56365 ^ t56365;
    wire t56367 = t56366 ^ t56366;
    wire t56368 = t56367 ^ t56367;
    wire t56369 = t56368 ^ t56368;
    wire t56370 = t56369 ^ t56369;
    wire t56371 = t56370 ^ t56370;
    wire t56372 = t56371 ^ t56371;
    wire t56373 = t56372 ^ t56372;
    wire t56374 = t56373 ^ t56373;
    wire t56375 = t56374 ^ t56374;
    wire t56376 = t56375 ^ t56375;
    wire t56377 = t56376 ^ t56376;
    wire t56378 = t56377 ^ t56377;
    wire t56379 = t56378 ^ t56378;
    wire t56380 = t56379 ^ t56379;
    wire t56381 = t56380 ^ t56380;
    wire t56382 = t56381 ^ t56381;
    wire t56383 = t56382 ^ t56382;
    wire t56384 = t56383 ^ t56383;
    wire t56385 = t56384 ^ t56384;
    wire t56386 = t56385 ^ t56385;
    wire t56387 = t56386 ^ t56386;
    wire t56388 = t56387 ^ t56387;
    wire t56389 = t56388 ^ t56388;
    wire t56390 = t56389 ^ t56389;
    wire t56391 = t56390 ^ t56390;
    wire t56392 = t56391 ^ t56391;
    wire t56393 = t56392 ^ t56392;
    wire t56394 = t56393 ^ t56393;
    wire t56395 = t56394 ^ t56394;
    wire t56396 = t56395 ^ t56395;
    wire t56397 = t56396 ^ t56396;
    wire t56398 = t56397 ^ t56397;
    wire t56399 = t56398 ^ t56398;
    wire t56400 = t56399 ^ t56399;
    wire t56401 = t56400 ^ t56400;
    wire t56402 = t56401 ^ t56401;
    wire t56403 = t56402 ^ t56402;
    wire t56404 = t56403 ^ t56403;
    wire t56405 = t56404 ^ t56404;
    wire t56406 = t56405 ^ t56405;
    wire t56407 = t56406 ^ t56406;
    wire t56408 = t56407 ^ t56407;
    wire t56409 = t56408 ^ t56408;
    wire t56410 = t56409 ^ t56409;
    wire t56411 = t56410 ^ t56410;
    wire t56412 = t56411 ^ t56411;
    wire t56413 = t56412 ^ t56412;
    wire t56414 = t56413 ^ t56413;
    wire t56415 = t56414 ^ t56414;
    wire t56416 = t56415 ^ t56415;
    wire t56417 = t56416 ^ t56416;
    wire t56418 = t56417 ^ t56417;
    wire t56419 = t56418 ^ t56418;
    wire t56420 = t56419 ^ t56419;
    wire t56421 = t56420 ^ t56420;
    wire t56422 = t56421 ^ t56421;
    wire t56423 = t56422 ^ t56422;
    wire t56424 = t56423 ^ t56423;
    wire t56425 = t56424 ^ t56424;
    wire t56426 = t56425 ^ t56425;
    wire t56427 = t56426 ^ t56426;
    wire t56428 = t56427 ^ t56427;
    wire t56429 = t56428 ^ t56428;
    wire t56430 = t56429 ^ t56429;
    wire t56431 = t56430 ^ t56430;
    wire t56432 = t56431 ^ t56431;
    wire t56433 = t56432 ^ t56432;
    wire t56434 = t56433 ^ t56433;
    wire t56435 = t56434 ^ t56434;
    wire t56436 = t56435 ^ t56435;
    wire t56437 = t56436 ^ t56436;
    wire t56438 = t56437 ^ t56437;
    wire t56439 = t56438 ^ t56438;
    wire t56440 = t56439 ^ t56439;
    wire t56441 = t56440 ^ t56440;
    wire t56442 = t56441 ^ t56441;
    wire t56443 = t56442 ^ t56442;
    wire t56444 = t56443 ^ t56443;
    wire t56445 = t56444 ^ t56444;
    wire t56446 = t56445 ^ t56445;
    wire t56447 = t56446 ^ t56446;
    wire t56448 = t56447 ^ t56447;
    wire t56449 = t56448 ^ t56448;
    wire t56450 = t56449 ^ t56449;
    wire t56451 = t56450 ^ t56450;
    wire t56452 = t56451 ^ t56451;
    wire t56453 = t56452 ^ t56452;
    wire t56454 = t56453 ^ t56453;
    wire t56455 = t56454 ^ t56454;
    wire t56456 = t56455 ^ t56455;
    wire t56457 = t56456 ^ t56456;
    wire t56458 = t56457 ^ t56457;
    wire t56459 = t56458 ^ t56458;
    wire t56460 = t56459 ^ t56459;
    wire t56461 = t56460 ^ t56460;
    wire t56462 = t56461 ^ t56461;
    wire t56463 = t56462 ^ t56462;
    wire t56464 = t56463 ^ t56463;
    wire t56465 = t56464 ^ t56464;
    wire t56466 = t56465 ^ t56465;
    wire t56467 = t56466 ^ t56466;
    wire t56468 = t56467 ^ t56467;
    wire t56469 = t56468 ^ t56468;
    wire t56470 = t56469 ^ t56469;
    wire t56471 = t56470 ^ t56470;
    wire t56472 = t56471 ^ t56471;
    wire t56473 = t56472 ^ t56472;
    wire t56474 = t56473 ^ t56473;
    wire t56475 = t56474 ^ t56474;
    wire t56476 = t56475 ^ t56475;
    wire t56477 = t56476 ^ t56476;
    wire t56478 = t56477 ^ t56477;
    wire t56479 = t56478 ^ t56478;
    wire t56480 = t56479 ^ t56479;
    wire t56481 = t56480 ^ t56480;
    wire t56482 = t56481 ^ t56481;
    wire t56483 = t56482 ^ t56482;
    wire t56484 = t56483 ^ t56483;
    wire t56485 = t56484 ^ t56484;
    wire t56486 = t56485 ^ t56485;
    wire t56487 = t56486 ^ t56486;
    wire t56488 = t56487 ^ t56487;
    wire t56489 = t56488 ^ t56488;
    wire t56490 = t56489 ^ t56489;
    wire t56491 = t56490 ^ t56490;
    wire t56492 = t56491 ^ t56491;
    wire t56493 = t56492 ^ t56492;
    wire t56494 = t56493 ^ t56493;
    wire t56495 = t56494 ^ t56494;
    wire t56496 = t56495 ^ t56495;
    wire t56497 = t56496 ^ t56496;
    wire t56498 = t56497 ^ t56497;
    wire t56499 = t56498 ^ t56498;
    wire t56500 = t56499 ^ t56499;
    wire t56501 = t56500 ^ t56500;
    wire t56502 = t56501 ^ t56501;
    wire t56503 = t56502 ^ t56502;
    wire t56504 = t56503 ^ t56503;
    wire t56505 = t56504 ^ t56504;
    wire t56506 = t56505 ^ t56505;
    wire t56507 = t56506 ^ t56506;
    wire t56508 = t56507 ^ t56507;
    wire t56509 = t56508 ^ t56508;
    wire t56510 = t56509 ^ t56509;
    wire t56511 = t56510 ^ t56510;
    wire t56512 = t56511 ^ t56511;
    wire t56513 = t56512 ^ t56512;
    wire t56514 = t56513 ^ t56513;
    wire t56515 = t56514 ^ t56514;
    wire t56516 = t56515 ^ t56515;
    wire t56517 = t56516 ^ t56516;
    wire t56518 = t56517 ^ t56517;
    wire t56519 = t56518 ^ t56518;
    wire t56520 = t56519 ^ t56519;
    wire t56521 = t56520 ^ t56520;
    wire t56522 = t56521 ^ t56521;
    wire t56523 = t56522 ^ t56522;
    wire t56524 = t56523 ^ t56523;
    wire t56525 = t56524 ^ t56524;
    wire t56526 = t56525 ^ t56525;
    wire t56527 = t56526 ^ t56526;
    wire t56528 = t56527 ^ t56527;
    wire t56529 = t56528 ^ t56528;
    wire t56530 = t56529 ^ t56529;
    wire t56531 = t56530 ^ t56530;
    wire t56532 = t56531 ^ t56531;
    wire t56533 = t56532 ^ t56532;
    wire t56534 = t56533 ^ t56533;
    wire t56535 = t56534 ^ t56534;
    wire t56536 = t56535 ^ t56535;
    wire t56537 = t56536 ^ t56536;
    wire t56538 = t56537 ^ t56537;
    wire t56539 = t56538 ^ t56538;
    wire t56540 = t56539 ^ t56539;
    wire t56541 = t56540 ^ t56540;
    wire t56542 = t56541 ^ t56541;
    wire t56543 = t56542 ^ t56542;
    wire t56544 = t56543 ^ t56543;
    wire t56545 = t56544 ^ t56544;
    wire t56546 = t56545 ^ t56545;
    wire t56547 = t56546 ^ t56546;
    wire t56548 = t56547 ^ t56547;
    wire t56549 = t56548 ^ t56548;
    wire t56550 = t56549 ^ t56549;
    wire t56551 = t56550 ^ t56550;
    wire t56552 = t56551 ^ t56551;
    wire t56553 = t56552 ^ t56552;
    wire t56554 = t56553 ^ t56553;
    wire t56555 = t56554 ^ t56554;
    wire t56556 = t56555 ^ t56555;
    wire t56557 = t56556 ^ t56556;
    wire t56558 = t56557 ^ t56557;
    wire t56559 = t56558 ^ t56558;
    wire t56560 = t56559 ^ t56559;
    wire t56561 = t56560 ^ t56560;
    wire t56562 = t56561 ^ t56561;
    wire t56563 = t56562 ^ t56562;
    wire t56564 = t56563 ^ t56563;
    wire t56565 = t56564 ^ t56564;
    wire t56566 = t56565 ^ t56565;
    wire t56567 = t56566 ^ t56566;
    wire t56568 = t56567 ^ t56567;
    wire t56569 = t56568 ^ t56568;
    wire t56570 = t56569 ^ t56569;
    wire t56571 = t56570 ^ t56570;
    wire t56572 = t56571 ^ t56571;
    wire t56573 = t56572 ^ t56572;
    wire t56574 = t56573 ^ t56573;
    wire t56575 = t56574 ^ t56574;
    wire t56576 = t56575 ^ t56575;
    wire t56577 = t56576 ^ t56576;
    wire t56578 = t56577 ^ t56577;
    wire t56579 = t56578 ^ t56578;
    wire t56580 = t56579 ^ t56579;
    wire t56581 = t56580 ^ t56580;
    wire t56582 = t56581 ^ t56581;
    wire t56583 = t56582 ^ t56582;
    wire t56584 = t56583 ^ t56583;
    wire t56585 = t56584 ^ t56584;
    wire t56586 = t56585 ^ t56585;
    wire t56587 = t56586 ^ t56586;
    wire t56588 = t56587 ^ t56587;
    wire t56589 = t56588 ^ t56588;
    wire t56590 = t56589 ^ t56589;
    wire t56591 = t56590 ^ t56590;
    wire t56592 = t56591 ^ t56591;
    wire t56593 = t56592 ^ t56592;
    wire t56594 = t56593 ^ t56593;
    wire t56595 = t56594 ^ t56594;
    wire t56596 = t56595 ^ t56595;
    wire t56597 = t56596 ^ t56596;
    wire t56598 = t56597 ^ t56597;
    wire t56599 = t56598 ^ t56598;
    wire t56600 = t56599 ^ t56599;
    wire t56601 = t56600 ^ t56600;
    wire t56602 = t56601 ^ t56601;
    wire t56603 = t56602 ^ t56602;
    wire t56604 = t56603 ^ t56603;
    wire t56605 = t56604 ^ t56604;
    wire t56606 = t56605 ^ t56605;
    wire t56607 = t56606 ^ t56606;
    wire t56608 = t56607 ^ t56607;
    wire t56609 = t56608 ^ t56608;
    wire t56610 = t56609 ^ t56609;
    wire t56611 = t56610 ^ t56610;
    wire t56612 = t56611 ^ t56611;
    wire t56613 = t56612 ^ t56612;
    wire t56614 = t56613 ^ t56613;
    wire t56615 = t56614 ^ t56614;
    wire t56616 = t56615 ^ t56615;
    wire t56617 = t56616 ^ t56616;
    wire t56618 = t56617 ^ t56617;
    wire t56619 = t56618 ^ t56618;
    wire t56620 = t56619 ^ t56619;
    wire t56621 = t56620 ^ t56620;
    wire t56622 = t56621 ^ t56621;
    wire t56623 = t56622 ^ t56622;
    wire t56624 = t56623 ^ t56623;
    wire t56625 = t56624 ^ t56624;
    wire t56626 = t56625 ^ t56625;
    wire t56627 = t56626 ^ t56626;
    wire t56628 = t56627 ^ t56627;
    wire t56629 = t56628 ^ t56628;
    wire t56630 = t56629 ^ t56629;
    wire t56631 = t56630 ^ t56630;
    wire t56632 = t56631 ^ t56631;
    wire t56633 = t56632 ^ t56632;
    wire t56634 = t56633 ^ t56633;
    wire t56635 = t56634 ^ t56634;
    wire t56636 = t56635 ^ t56635;
    wire t56637 = t56636 ^ t56636;
    wire t56638 = t56637 ^ t56637;
    wire t56639 = t56638 ^ t56638;
    wire t56640 = t56639 ^ t56639;
    wire t56641 = t56640 ^ t56640;
    wire t56642 = t56641 ^ t56641;
    wire t56643 = t56642 ^ t56642;
    wire t56644 = t56643 ^ t56643;
    wire t56645 = t56644 ^ t56644;
    wire t56646 = t56645 ^ t56645;
    wire t56647 = t56646 ^ t56646;
    wire t56648 = t56647 ^ t56647;
    wire t56649 = t56648 ^ t56648;
    wire t56650 = t56649 ^ t56649;
    wire t56651 = t56650 ^ t56650;
    wire t56652 = t56651 ^ t56651;
    wire t56653 = t56652 ^ t56652;
    wire t56654 = t56653 ^ t56653;
    wire t56655 = t56654 ^ t56654;
    wire t56656 = t56655 ^ t56655;
    wire t56657 = t56656 ^ t56656;
    wire t56658 = t56657 ^ t56657;
    wire t56659 = t56658 ^ t56658;
    wire t56660 = t56659 ^ t56659;
    wire t56661 = t56660 ^ t56660;
    wire t56662 = t56661 ^ t56661;
    wire t56663 = t56662 ^ t56662;
    wire t56664 = t56663 ^ t56663;
    wire t56665 = t56664 ^ t56664;
    wire t56666 = t56665 ^ t56665;
    wire t56667 = t56666 ^ t56666;
    wire t56668 = t56667 ^ t56667;
    wire t56669 = t56668 ^ t56668;
    wire t56670 = t56669 ^ t56669;
    wire t56671 = t56670 ^ t56670;
    wire t56672 = t56671 ^ t56671;
    wire t56673 = t56672 ^ t56672;
    wire t56674 = t56673 ^ t56673;
    wire t56675 = t56674 ^ t56674;
    wire t56676 = t56675 ^ t56675;
    wire t56677 = t56676 ^ t56676;
    wire t56678 = t56677 ^ t56677;
    wire t56679 = t56678 ^ t56678;
    wire t56680 = t56679 ^ t56679;
    wire t56681 = t56680 ^ t56680;
    wire t56682 = t56681 ^ t56681;
    wire t56683 = t56682 ^ t56682;
    wire t56684 = t56683 ^ t56683;
    wire t56685 = t56684 ^ t56684;
    wire t56686 = t56685 ^ t56685;
    wire t56687 = t56686 ^ t56686;
    wire t56688 = t56687 ^ t56687;
    wire t56689 = t56688 ^ t56688;
    wire t56690 = t56689 ^ t56689;
    wire t56691 = t56690 ^ t56690;
    wire t56692 = t56691 ^ t56691;
    wire t56693 = t56692 ^ t56692;
    wire t56694 = t56693 ^ t56693;
    wire t56695 = t56694 ^ t56694;
    wire t56696 = t56695 ^ t56695;
    wire t56697 = t56696 ^ t56696;
    wire t56698 = t56697 ^ t56697;
    wire t56699 = t56698 ^ t56698;
    wire t56700 = t56699 ^ t56699;
    wire t56701 = t56700 ^ t56700;
    wire t56702 = t56701 ^ t56701;
    wire t56703 = t56702 ^ t56702;
    wire t56704 = t56703 ^ t56703;
    wire t56705 = t56704 ^ t56704;
    wire t56706 = t56705 ^ t56705;
    wire t56707 = t56706 ^ t56706;
    wire t56708 = t56707 ^ t56707;
    wire t56709 = t56708 ^ t56708;
    wire t56710 = t56709 ^ t56709;
    wire t56711 = t56710 ^ t56710;
    wire t56712 = t56711 ^ t56711;
    wire t56713 = t56712 ^ t56712;
    wire t56714 = t56713 ^ t56713;
    wire t56715 = t56714 ^ t56714;
    wire t56716 = t56715 ^ t56715;
    wire t56717 = t56716 ^ t56716;
    wire t56718 = t56717 ^ t56717;
    wire t56719 = t56718 ^ t56718;
    wire t56720 = t56719 ^ t56719;
    wire t56721 = t56720 ^ t56720;
    wire t56722 = t56721 ^ t56721;
    wire t56723 = t56722 ^ t56722;
    wire t56724 = t56723 ^ t56723;
    wire t56725 = t56724 ^ t56724;
    wire t56726 = t56725 ^ t56725;
    wire t56727 = t56726 ^ t56726;
    wire t56728 = t56727 ^ t56727;
    wire t56729 = t56728 ^ t56728;
    wire t56730 = t56729 ^ t56729;
    wire t56731 = t56730 ^ t56730;
    wire t56732 = t56731 ^ t56731;
    wire t56733 = t56732 ^ t56732;
    wire t56734 = t56733 ^ t56733;
    wire t56735 = t56734 ^ t56734;
    wire t56736 = t56735 ^ t56735;
    wire t56737 = t56736 ^ t56736;
    wire t56738 = t56737 ^ t56737;
    wire t56739 = t56738 ^ t56738;
    wire t56740 = t56739 ^ t56739;
    wire t56741 = t56740 ^ t56740;
    wire t56742 = t56741 ^ t56741;
    wire t56743 = t56742 ^ t56742;
    wire t56744 = t56743 ^ t56743;
    wire t56745 = t56744 ^ t56744;
    wire t56746 = t56745 ^ t56745;
    wire t56747 = t56746 ^ t56746;
    wire t56748 = t56747 ^ t56747;
    wire t56749 = t56748 ^ t56748;
    wire t56750 = t56749 ^ t56749;
    wire t56751 = t56750 ^ t56750;
    wire t56752 = t56751 ^ t56751;
    wire t56753 = t56752 ^ t56752;
    wire t56754 = t56753 ^ t56753;
    wire t56755 = t56754 ^ t56754;
    wire t56756 = t56755 ^ t56755;
    wire t56757 = t56756 ^ t56756;
    wire t56758 = t56757 ^ t56757;
    wire t56759 = t56758 ^ t56758;
    wire t56760 = t56759 ^ t56759;
    wire t56761 = t56760 ^ t56760;
    wire t56762 = t56761 ^ t56761;
    wire t56763 = t56762 ^ t56762;
    wire t56764 = t56763 ^ t56763;
    wire t56765 = t56764 ^ t56764;
    wire t56766 = t56765 ^ t56765;
    wire t56767 = t56766 ^ t56766;
    wire t56768 = t56767 ^ t56767;
    wire t56769 = t56768 ^ t56768;
    wire t56770 = t56769 ^ t56769;
    wire t56771 = t56770 ^ t56770;
    wire t56772 = t56771 ^ t56771;
    wire t56773 = t56772 ^ t56772;
    wire t56774 = t56773 ^ t56773;
    wire t56775 = t56774 ^ t56774;
    wire t56776 = t56775 ^ t56775;
    wire t56777 = t56776 ^ t56776;
    wire t56778 = t56777 ^ t56777;
    wire t56779 = t56778 ^ t56778;
    wire t56780 = t56779 ^ t56779;
    wire t56781 = t56780 ^ t56780;
    wire t56782 = t56781 ^ t56781;
    wire t56783 = t56782 ^ t56782;
    wire t56784 = t56783 ^ t56783;
    wire t56785 = t56784 ^ t56784;
    wire t56786 = t56785 ^ t56785;
    wire t56787 = t56786 ^ t56786;
    wire t56788 = t56787 ^ t56787;
    wire t56789 = t56788 ^ t56788;
    wire t56790 = t56789 ^ t56789;
    wire t56791 = t56790 ^ t56790;
    wire t56792 = t56791 ^ t56791;
    wire t56793 = t56792 ^ t56792;
    wire t56794 = t56793 ^ t56793;
    wire t56795 = t56794 ^ t56794;
    wire t56796 = t56795 ^ t56795;
    wire t56797 = t56796 ^ t56796;
    wire t56798 = t56797 ^ t56797;
    wire t56799 = t56798 ^ t56798;
    wire t56800 = t56799 ^ t56799;
    wire t56801 = t56800 ^ t56800;
    wire t56802 = t56801 ^ t56801;
    wire t56803 = t56802 ^ t56802;
    wire t56804 = t56803 ^ t56803;
    wire t56805 = t56804 ^ t56804;
    wire t56806 = t56805 ^ t56805;
    wire t56807 = t56806 ^ t56806;
    wire t56808 = t56807 ^ t56807;
    wire t56809 = t56808 ^ t56808;
    wire t56810 = t56809 ^ t56809;
    wire t56811 = t56810 ^ t56810;
    wire t56812 = t56811 ^ t56811;
    wire t56813 = t56812 ^ t56812;
    wire t56814 = t56813 ^ t56813;
    wire t56815 = t56814 ^ t56814;
    wire t56816 = t56815 ^ t56815;
    wire t56817 = t56816 ^ t56816;
    wire t56818 = t56817 ^ t56817;
    wire t56819 = t56818 ^ t56818;
    wire t56820 = t56819 ^ t56819;
    wire t56821 = t56820 ^ t56820;
    wire t56822 = t56821 ^ t56821;
    wire t56823 = t56822 ^ t56822;
    wire t56824 = t56823 ^ t56823;
    wire t56825 = t56824 ^ t56824;
    wire t56826 = t56825 ^ t56825;
    wire t56827 = t56826 ^ t56826;
    wire t56828 = t56827 ^ t56827;
    wire t56829 = t56828 ^ t56828;
    wire t56830 = t56829 ^ t56829;
    wire t56831 = t56830 ^ t56830;
    wire t56832 = t56831 ^ t56831;
    wire t56833 = t56832 ^ t56832;
    wire t56834 = t56833 ^ t56833;
    wire t56835 = t56834 ^ t56834;
    wire t56836 = t56835 ^ t56835;
    wire t56837 = t56836 ^ t56836;
    wire t56838 = t56837 ^ t56837;
    wire t56839 = t56838 ^ t56838;
    wire t56840 = t56839 ^ t56839;
    wire t56841 = t56840 ^ t56840;
    wire t56842 = t56841 ^ t56841;
    wire t56843 = t56842 ^ t56842;
    wire t56844 = t56843 ^ t56843;
    wire t56845 = t56844 ^ t56844;
    wire t56846 = t56845 ^ t56845;
    wire t56847 = t56846 ^ t56846;
    wire t56848 = t56847 ^ t56847;
    wire t56849 = t56848 ^ t56848;
    wire t56850 = t56849 ^ t56849;
    wire t56851 = t56850 ^ t56850;
    wire t56852 = t56851 ^ t56851;
    wire t56853 = t56852 ^ t56852;
    wire t56854 = t56853 ^ t56853;
    wire t56855 = t56854 ^ t56854;
    wire t56856 = t56855 ^ t56855;
    wire t56857 = t56856 ^ t56856;
    wire t56858 = t56857 ^ t56857;
    wire t56859 = t56858 ^ t56858;
    wire t56860 = t56859 ^ t56859;
    wire t56861 = t56860 ^ t56860;
    wire t56862 = t56861 ^ t56861;
    wire t56863 = t56862 ^ t56862;
    wire t56864 = t56863 ^ t56863;
    wire t56865 = t56864 ^ t56864;
    wire t56866 = t56865 ^ t56865;
    wire t56867 = t56866 ^ t56866;
    wire t56868 = t56867 ^ t56867;
    wire t56869 = t56868 ^ t56868;
    wire t56870 = t56869 ^ t56869;
    wire t56871 = t56870 ^ t56870;
    wire t56872 = t56871 ^ t56871;
    wire t56873 = t56872 ^ t56872;
    wire t56874 = t56873 ^ t56873;
    wire t56875 = t56874 ^ t56874;
    wire t56876 = t56875 ^ t56875;
    wire t56877 = t56876 ^ t56876;
    wire t56878 = t56877 ^ t56877;
    wire t56879 = t56878 ^ t56878;
    wire t56880 = t56879 ^ t56879;
    wire t56881 = t56880 ^ t56880;
    wire t56882 = t56881 ^ t56881;
    wire t56883 = t56882 ^ t56882;
    wire t56884 = t56883 ^ t56883;
    wire t56885 = t56884 ^ t56884;
    wire t56886 = t56885 ^ t56885;
    wire t56887 = t56886 ^ t56886;
    wire t56888 = t56887 ^ t56887;
    wire t56889 = t56888 ^ t56888;
    wire t56890 = t56889 ^ t56889;
    wire t56891 = t56890 ^ t56890;
    wire t56892 = t56891 ^ t56891;
    wire t56893 = t56892 ^ t56892;
    wire t56894 = t56893 ^ t56893;
    wire t56895 = t56894 ^ t56894;
    wire t56896 = t56895 ^ t56895;
    wire t56897 = t56896 ^ t56896;
    wire t56898 = t56897 ^ t56897;
    wire t56899 = t56898 ^ t56898;
    wire t56900 = t56899 ^ t56899;
    wire t56901 = t56900 ^ t56900;
    wire t56902 = t56901 ^ t56901;
    wire t56903 = t56902 ^ t56902;
    wire t56904 = t56903 ^ t56903;
    wire t56905 = t56904 ^ t56904;
    wire t56906 = t56905 ^ t56905;
    wire t56907 = t56906 ^ t56906;
    wire t56908 = t56907 ^ t56907;
    wire t56909 = t56908 ^ t56908;
    wire t56910 = t56909 ^ t56909;
    wire t56911 = t56910 ^ t56910;
    wire t56912 = t56911 ^ t56911;
    wire t56913 = t56912 ^ t56912;
    wire t56914 = t56913 ^ t56913;
    wire t56915 = t56914 ^ t56914;
    wire t56916 = t56915 ^ t56915;
    wire t56917 = t56916 ^ t56916;
    wire t56918 = t56917 ^ t56917;
    wire t56919 = t56918 ^ t56918;
    wire t56920 = t56919 ^ t56919;
    wire t56921 = t56920 ^ t56920;
    wire t56922 = t56921 ^ t56921;
    wire t56923 = t56922 ^ t56922;
    wire t56924 = t56923 ^ t56923;
    wire t56925 = t56924 ^ t56924;
    wire t56926 = t56925 ^ t56925;
    wire t56927 = t56926 ^ t56926;
    wire t56928 = t56927 ^ t56927;
    wire t56929 = t56928 ^ t56928;
    wire t56930 = t56929 ^ t56929;
    wire t56931 = t56930 ^ t56930;
    wire t56932 = t56931 ^ t56931;
    wire t56933 = t56932 ^ t56932;
    wire t56934 = t56933 ^ t56933;
    wire t56935 = t56934 ^ t56934;
    wire t56936 = t56935 ^ t56935;
    wire t56937 = t56936 ^ t56936;
    wire t56938 = t56937 ^ t56937;
    wire t56939 = t56938 ^ t56938;
    wire t56940 = t56939 ^ t56939;
    wire t56941 = t56940 ^ t56940;
    wire t56942 = t56941 ^ t56941;
    wire t56943 = t56942 ^ t56942;
    wire t56944 = t56943 ^ t56943;
    wire t56945 = t56944 ^ t56944;
    wire t56946 = t56945 ^ t56945;
    wire t56947 = t56946 ^ t56946;
    wire t56948 = t56947 ^ t56947;
    wire t56949 = t56948 ^ t56948;
    wire t56950 = t56949 ^ t56949;
    wire t56951 = t56950 ^ t56950;
    wire t56952 = t56951 ^ t56951;
    wire t56953 = t56952 ^ t56952;
    wire t56954 = t56953 ^ t56953;
    wire t56955 = t56954 ^ t56954;
    wire t56956 = t56955 ^ t56955;
    wire t56957 = t56956 ^ t56956;
    wire t56958 = t56957 ^ t56957;
    wire t56959 = t56958 ^ t56958;
    wire t56960 = t56959 ^ t56959;
    wire t56961 = t56960 ^ t56960;
    wire t56962 = t56961 ^ t56961;
    wire t56963 = t56962 ^ t56962;
    wire t56964 = t56963 ^ t56963;
    wire t56965 = t56964 ^ t56964;
    wire t56966 = t56965 ^ t56965;
    wire t56967 = t56966 ^ t56966;
    wire t56968 = t56967 ^ t56967;
    wire t56969 = t56968 ^ t56968;
    wire t56970 = t56969 ^ t56969;
    wire t56971 = t56970 ^ t56970;
    wire t56972 = t56971 ^ t56971;
    wire t56973 = t56972 ^ t56972;
    wire t56974 = t56973 ^ t56973;
    wire t56975 = t56974 ^ t56974;
    wire t56976 = t56975 ^ t56975;
    wire t56977 = t56976 ^ t56976;
    wire t56978 = t56977 ^ t56977;
    wire t56979 = t56978 ^ t56978;
    wire t56980 = t56979 ^ t56979;
    wire t56981 = t56980 ^ t56980;
    wire t56982 = t56981 ^ t56981;
    wire t56983 = t56982 ^ t56982;
    wire t56984 = t56983 ^ t56983;
    wire t56985 = t56984 ^ t56984;
    wire t56986 = t56985 ^ t56985;
    wire t56987 = t56986 ^ t56986;
    wire t56988 = t56987 ^ t56987;
    wire t56989 = t56988 ^ t56988;
    wire t56990 = t56989 ^ t56989;
    wire t56991 = t56990 ^ t56990;
    wire t56992 = t56991 ^ t56991;
    wire t56993 = t56992 ^ t56992;
    wire t56994 = t56993 ^ t56993;
    wire t56995 = t56994 ^ t56994;
    wire t56996 = t56995 ^ t56995;
    wire t56997 = t56996 ^ t56996;
    wire t56998 = t56997 ^ t56997;
    wire t56999 = t56998 ^ t56998;
    wire t57000 = t56999 ^ t56999;
    wire t57001 = t57000 ^ t57000;
    wire t57002 = t57001 ^ t57001;
    wire t57003 = t57002 ^ t57002;
    wire t57004 = t57003 ^ t57003;
    wire t57005 = t57004 ^ t57004;
    wire t57006 = t57005 ^ t57005;
    wire t57007 = t57006 ^ t57006;
    wire t57008 = t57007 ^ t57007;
    wire t57009 = t57008 ^ t57008;
    wire t57010 = t57009 ^ t57009;
    wire t57011 = t57010 ^ t57010;
    wire t57012 = t57011 ^ t57011;
    wire t57013 = t57012 ^ t57012;
    wire t57014 = t57013 ^ t57013;
    wire t57015 = t57014 ^ t57014;
    wire t57016 = t57015 ^ t57015;
    wire t57017 = t57016 ^ t57016;
    wire t57018 = t57017 ^ t57017;
    wire t57019 = t57018 ^ t57018;
    wire t57020 = t57019 ^ t57019;
    wire t57021 = t57020 ^ t57020;
    wire t57022 = t57021 ^ t57021;
    wire t57023 = t57022 ^ t57022;
    wire t57024 = t57023 ^ t57023;
    wire t57025 = t57024 ^ t57024;
    wire t57026 = t57025 ^ t57025;
    wire t57027 = t57026 ^ t57026;
    wire t57028 = t57027 ^ t57027;
    wire t57029 = t57028 ^ t57028;
    wire t57030 = t57029 ^ t57029;
    wire t57031 = t57030 ^ t57030;
    wire t57032 = t57031 ^ t57031;
    wire t57033 = t57032 ^ t57032;
    wire t57034 = t57033 ^ t57033;
    wire t57035 = t57034 ^ t57034;
    wire t57036 = t57035 ^ t57035;
    wire t57037 = t57036 ^ t57036;
    wire t57038 = t57037 ^ t57037;
    wire t57039 = t57038 ^ t57038;
    wire t57040 = t57039 ^ t57039;
    wire t57041 = t57040 ^ t57040;
    wire t57042 = t57041 ^ t57041;
    wire t57043 = t57042 ^ t57042;
    wire t57044 = t57043 ^ t57043;
    wire t57045 = t57044 ^ t57044;
    wire t57046 = t57045 ^ t57045;
    wire t57047 = t57046 ^ t57046;
    wire t57048 = t57047 ^ t57047;
    wire t57049 = t57048 ^ t57048;
    wire t57050 = t57049 ^ t57049;
    wire t57051 = t57050 ^ t57050;
    wire t57052 = t57051 ^ t57051;
    wire t57053 = t57052 ^ t57052;
    wire t57054 = t57053 ^ t57053;
    wire t57055 = t57054 ^ t57054;
    wire t57056 = t57055 ^ t57055;
    wire t57057 = t57056 ^ t57056;
    wire t57058 = t57057 ^ t57057;
    wire t57059 = t57058 ^ t57058;
    wire t57060 = t57059 ^ t57059;
    wire t57061 = t57060 ^ t57060;
    wire t57062 = t57061 ^ t57061;
    wire t57063 = t57062 ^ t57062;
    wire t57064 = t57063 ^ t57063;
    wire t57065 = t57064 ^ t57064;
    wire t57066 = t57065 ^ t57065;
    wire t57067 = t57066 ^ t57066;
    wire t57068 = t57067 ^ t57067;
    wire t57069 = t57068 ^ t57068;
    wire t57070 = t57069 ^ t57069;
    wire t57071 = t57070 ^ t57070;
    wire t57072 = t57071 ^ t57071;
    wire t57073 = t57072 ^ t57072;
    wire t57074 = t57073 ^ t57073;
    wire t57075 = t57074 ^ t57074;
    wire t57076 = t57075 ^ t57075;
    wire t57077 = t57076 ^ t57076;
    wire t57078 = t57077 ^ t57077;
    wire t57079 = t57078 ^ t57078;
    wire t57080 = t57079 ^ t57079;
    wire t57081 = t57080 ^ t57080;
    wire t57082 = t57081 ^ t57081;
    wire t57083 = t57082 ^ t57082;
    wire t57084 = t57083 ^ t57083;
    wire t57085 = t57084 ^ t57084;
    wire t57086 = t57085 ^ t57085;
    wire t57087 = t57086 ^ t57086;
    wire t57088 = t57087 ^ t57087;
    wire t57089 = t57088 ^ t57088;
    wire t57090 = t57089 ^ t57089;
    wire t57091 = t57090 ^ t57090;
    wire t57092 = t57091 ^ t57091;
    wire t57093 = t57092 ^ t57092;
    wire t57094 = t57093 ^ t57093;
    wire t57095 = t57094 ^ t57094;
    wire t57096 = t57095 ^ t57095;
    wire t57097 = t57096 ^ t57096;
    wire t57098 = t57097 ^ t57097;
    wire t57099 = t57098 ^ t57098;
    wire t57100 = t57099 ^ t57099;
    wire t57101 = t57100 ^ t57100;
    wire t57102 = t57101 ^ t57101;
    wire t57103 = t57102 ^ t57102;
    wire t57104 = t57103 ^ t57103;
    wire t57105 = t57104 ^ t57104;
    wire t57106 = t57105 ^ t57105;
    wire t57107 = t57106 ^ t57106;
    wire t57108 = t57107 ^ t57107;
    wire t57109 = t57108 ^ t57108;
    wire t57110 = t57109 ^ t57109;
    wire t57111 = t57110 ^ t57110;
    wire t57112 = t57111 ^ t57111;
    wire t57113 = t57112 ^ t57112;
    wire t57114 = t57113 ^ t57113;
    wire t57115 = t57114 ^ t57114;
    wire t57116 = t57115 ^ t57115;
    wire t57117 = t57116 ^ t57116;
    wire t57118 = t57117 ^ t57117;
    wire t57119 = t57118 ^ t57118;
    wire t57120 = t57119 ^ t57119;
    wire t57121 = t57120 ^ t57120;
    wire t57122 = t57121 ^ t57121;
    wire t57123 = t57122 ^ t57122;
    wire t57124 = t57123 ^ t57123;
    wire t57125 = t57124 ^ t57124;
    wire t57126 = t57125 ^ t57125;
    wire t57127 = t57126 ^ t57126;
    wire t57128 = t57127 ^ t57127;
    wire t57129 = t57128 ^ t57128;
    wire t57130 = t57129 ^ t57129;
    wire t57131 = t57130 ^ t57130;
    wire t57132 = t57131 ^ t57131;
    wire t57133 = t57132 ^ t57132;
    wire t57134 = t57133 ^ t57133;
    wire t57135 = t57134 ^ t57134;
    wire t57136 = t57135 ^ t57135;
    wire t57137 = t57136 ^ t57136;
    wire t57138 = t57137 ^ t57137;
    wire t57139 = t57138 ^ t57138;
    wire t57140 = t57139 ^ t57139;
    wire t57141 = t57140 ^ t57140;
    wire t57142 = t57141 ^ t57141;
    wire t57143 = t57142 ^ t57142;
    wire t57144 = t57143 ^ t57143;
    wire t57145 = t57144 ^ t57144;
    wire t57146 = t57145 ^ t57145;
    wire t57147 = t57146 ^ t57146;
    wire t57148 = t57147 ^ t57147;
    wire t57149 = t57148 ^ t57148;
    wire t57150 = t57149 ^ t57149;
    wire t57151 = t57150 ^ t57150;
    wire t57152 = t57151 ^ t57151;
    wire t57153 = t57152 ^ t57152;
    wire t57154 = t57153 ^ t57153;
    wire t57155 = t57154 ^ t57154;
    wire t57156 = t57155 ^ t57155;
    wire t57157 = t57156 ^ t57156;
    wire t57158 = t57157 ^ t57157;
    wire t57159 = t57158 ^ t57158;
    wire t57160 = t57159 ^ t57159;
    wire t57161 = t57160 ^ t57160;
    wire t57162 = t57161 ^ t57161;
    wire t57163 = t57162 ^ t57162;
    wire t57164 = t57163 ^ t57163;
    wire t57165 = t57164 ^ t57164;
    wire t57166 = t57165 ^ t57165;
    wire t57167 = t57166 ^ t57166;
    wire t57168 = t57167 ^ t57167;
    wire t57169 = t57168 ^ t57168;
    wire t57170 = t57169 ^ t57169;
    wire t57171 = t57170 ^ t57170;
    wire t57172 = t57171 ^ t57171;
    wire t57173 = t57172 ^ t57172;
    wire t57174 = t57173 ^ t57173;
    wire t57175 = t57174 ^ t57174;
    wire t57176 = t57175 ^ t57175;
    wire t57177 = t57176 ^ t57176;
    wire t57178 = t57177 ^ t57177;
    wire t57179 = t57178 ^ t57178;
    wire t57180 = t57179 ^ t57179;
    wire t57181 = t57180 ^ t57180;
    wire t57182 = t57181 ^ t57181;
    wire t57183 = t57182 ^ t57182;
    wire t57184 = t57183 ^ t57183;
    wire t57185 = t57184 ^ t57184;
    wire t57186 = t57185 ^ t57185;
    wire t57187 = t57186 ^ t57186;
    wire t57188 = t57187 ^ t57187;
    wire t57189 = t57188 ^ t57188;
    wire t57190 = t57189 ^ t57189;
    wire t57191 = t57190 ^ t57190;
    wire t57192 = t57191 ^ t57191;
    wire t57193 = t57192 ^ t57192;
    wire t57194 = t57193 ^ t57193;
    wire t57195 = t57194 ^ t57194;
    wire t57196 = t57195 ^ t57195;
    wire t57197 = t57196 ^ t57196;
    wire t57198 = t57197 ^ t57197;
    wire t57199 = t57198 ^ t57198;
    wire t57200 = t57199 ^ t57199;
    wire t57201 = t57200 ^ t57200;
    wire t57202 = t57201 ^ t57201;
    wire t57203 = t57202 ^ t57202;
    wire t57204 = t57203 ^ t57203;
    wire t57205 = t57204 ^ t57204;
    wire t57206 = t57205 ^ t57205;
    wire t57207 = t57206 ^ t57206;
    wire t57208 = t57207 ^ t57207;
    wire t57209 = t57208 ^ t57208;
    wire t57210 = t57209 ^ t57209;
    wire t57211 = t57210 ^ t57210;
    wire t57212 = t57211 ^ t57211;
    wire t57213 = t57212 ^ t57212;
    wire t57214 = t57213 ^ t57213;
    wire t57215 = t57214 ^ t57214;
    wire t57216 = t57215 ^ t57215;
    wire t57217 = t57216 ^ t57216;
    wire t57218 = t57217 ^ t57217;
    wire t57219 = t57218 ^ t57218;
    wire t57220 = t57219 ^ t57219;
    wire t57221 = t57220 ^ t57220;
    wire t57222 = t57221 ^ t57221;
    wire t57223 = t57222 ^ t57222;
    wire t57224 = t57223 ^ t57223;
    wire t57225 = t57224 ^ t57224;
    wire t57226 = t57225 ^ t57225;
    wire t57227 = t57226 ^ t57226;
    wire t57228 = t57227 ^ t57227;
    wire t57229 = t57228 ^ t57228;
    wire t57230 = t57229 ^ t57229;
    wire t57231 = t57230 ^ t57230;
    wire t57232 = t57231 ^ t57231;
    wire t57233 = t57232 ^ t57232;
    wire t57234 = t57233 ^ t57233;
    wire t57235 = t57234 ^ t57234;
    wire t57236 = t57235 ^ t57235;
    wire t57237 = t57236 ^ t57236;
    wire t57238 = t57237 ^ t57237;
    wire t57239 = t57238 ^ t57238;
    wire t57240 = t57239 ^ t57239;
    wire t57241 = t57240 ^ t57240;
    wire t57242 = t57241 ^ t57241;
    wire t57243 = t57242 ^ t57242;
    wire t57244 = t57243 ^ t57243;
    wire t57245 = t57244 ^ t57244;
    wire t57246 = t57245 ^ t57245;
    wire t57247 = t57246 ^ t57246;
    wire t57248 = t57247 ^ t57247;
    wire t57249 = t57248 ^ t57248;
    wire t57250 = t57249 ^ t57249;
    wire t57251 = t57250 ^ t57250;
    wire t57252 = t57251 ^ t57251;
    wire t57253 = t57252 ^ t57252;
    wire t57254 = t57253 ^ t57253;
    wire t57255 = t57254 ^ t57254;
    wire t57256 = t57255 ^ t57255;
    wire t57257 = t57256 ^ t57256;
    wire t57258 = t57257 ^ t57257;
    wire t57259 = t57258 ^ t57258;
    wire t57260 = t57259 ^ t57259;
    wire t57261 = t57260 ^ t57260;
    wire t57262 = t57261 ^ t57261;
    wire t57263 = t57262 ^ t57262;
    wire t57264 = t57263 ^ t57263;
    wire t57265 = t57264 ^ t57264;
    wire t57266 = t57265 ^ t57265;
    wire t57267 = t57266 ^ t57266;
    wire t57268 = t57267 ^ t57267;
    wire t57269 = t57268 ^ t57268;
    wire t57270 = t57269 ^ t57269;
    wire t57271 = t57270 ^ t57270;
    wire t57272 = t57271 ^ t57271;
    wire t57273 = t57272 ^ t57272;
    wire t57274 = t57273 ^ t57273;
    wire t57275 = t57274 ^ t57274;
    wire t57276 = t57275 ^ t57275;
    wire t57277 = t57276 ^ t57276;
    wire t57278 = t57277 ^ t57277;
    wire t57279 = t57278 ^ t57278;
    wire t57280 = t57279 ^ t57279;
    wire t57281 = t57280 ^ t57280;
    wire t57282 = t57281 ^ t57281;
    wire t57283 = t57282 ^ t57282;
    wire t57284 = t57283 ^ t57283;
    wire t57285 = t57284 ^ t57284;
    wire t57286 = t57285 ^ t57285;
    wire t57287 = t57286 ^ t57286;
    wire t57288 = t57287 ^ t57287;
    wire t57289 = t57288 ^ t57288;
    wire t57290 = t57289 ^ t57289;
    wire t57291 = t57290 ^ t57290;
    wire t57292 = t57291 ^ t57291;
    wire t57293 = t57292 ^ t57292;
    wire t57294 = t57293 ^ t57293;
    wire t57295 = t57294 ^ t57294;
    wire t57296 = t57295 ^ t57295;
    wire t57297 = t57296 ^ t57296;
    wire t57298 = t57297 ^ t57297;
    wire t57299 = t57298 ^ t57298;
    wire t57300 = t57299 ^ t57299;
    wire t57301 = t57300 ^ t57300;
    wire t57302 = t57301 ^ t57301;
    wire t57303 = t57302 ^ t57302;
    wire t57304 = t57303 ^ t57303;
    wire t57305 = t57304 ^ t57304;
    wire t57306 = t57305 ^ t57305;
    wire t57307 = t57306 ^ t57306;
    wire t57308 = t57307 ^ t57307;
    wire t57309 = t57308 ^ t57308;
    wire t57310 = t57309 ^ t57309;
    wire t57311 = t57310 ^ t57310;
    wire t57312 = t57311 ^ t57311;
    wire t57313 = t57312 ^ t57312;
    wire t57314 = t57313 ^ t57313;
    wire t57315 = t57314 ^ t57314;
    wire t57316 = t57315 ^ t57315;
    wire t57317 = t57316 ^ t57316;
    wire t57318 = t57317 ^ t57317;
    wire t57319 = t57318 ^ t57318;
    wire t57320 = t57319 ^ t57319;
    wire t57321 = t57320 ^ t57320;
    wire t57322 = t57321 ^ t57321;
    wire t57323 = t57322 ^ t57322;
    wire t57324 = t57323 ^ t57323;
    wire t57325 = t57324 ^ t57324;
    wire t57326 = t57325 ^ t57325;
    wire t57327 = t57326 ^ t57326;
    wire t57328 = t57327 ^ t57327;
    wire t57329 = t57328 ^ t57328;
    wire t57330 = t57329 ^ t57329;
    wire t57331 = t57330 ^ t57330;
    wire t57332 = t57331 ^ t57331;
    wire t57333 = t57332 ^ t57332;
    wire t57334 = t57333 ^ t57333;
    wire t57335 = t57334 ^ t57334;
    wire t57336 = t57335 ^ t57335;
    wire t57337 = t57336 ^ t57336;
    wire t57338 = t57337 ^ t57337;
    wire t57339 = t57338 ^ t57338;
    wire t57340 = t57339 ^ t57339;
    wire t57341 = t57340 ^ t57340;
    wire t57342 = t57341 ^ t57341;
    wire t57343 = t57342 ^ t57342;
    wire t57344 = t57343 ^ t57343;
    wire t57345 = t57344 ^ t57344;
    wire t57346 = t57345 ^ t57345;
    wire t57347 = t57346 ^ t57346;
    wire t57348 = t57347 ^ t57347;
    wire t57349 = t57348 ^ t57348;
    wire t57350 = t57349 ^ t57349;
    wire t57351 = t57350 ^ t57350;
    wire t57352 = t57351 ^ t57351;
    wire t57353 = t57352 ^ t57352;
    wire t57354 = t57353 ^ t57353;
    wire t57355 = t57354 ^ t57354;
    wire t57356 = t57355 ^ t57355;
    wire t57357 = t57356 ^ t57356;
    wire t57358 = t57357 ^ t57357;
    wire t57359 = t57358 ^ t57358;
    wire t57360 = t57359 ^ t57359;
    wire t57361 = t57360 ^ t57360;
    wire t57362 = t57361 ^ t57361;
    wire t57363 = t57362 ^ t57362;
    wire t57364 = t57363 ^ t57363;
    wire t57365 = t57364 ^ t57364;
    wire t57366 = t57365 ^ t57365;
    wire t57367 = t57366 ^ t57366;
    wire t57368 = t57367 ^ t57367;
    wire t57369 = t57368 ^ t57368;
    wire t57370 = t57369 ^ t57369;
    wire t57371 = t57370 ^ t57370;
    wire t57372 = t57371 ^ t57371;
    wire t57373 = t57372 ^ t57372;
    wire t57374 = t57373 ^ t57373;
    wire t57375 = t57374 ^ t57374;
    wire t57376 = t57375 ^ t57375;
    wire t57377 = t57376 ^ t57376;
    wire t57378 = t57377 ^ t57377;
    wire t57379 = t57378 ^ t57378;
    wire t57380 = t57379 ^ t57379;
    wire t57381 = t57380 ^ t57380;
    wire t57382 = t57381 ^ t57381;
    wire t57383 = t57382 ^ t57382;
    wire t57384 = t57383 ^ t57383;
    wire t57385 = t57384 ^ t57384;
    wire t57386 = t57385 ^ t57385;
    wire t57387 = t57386 ^ t57386;
    wire t57388 = t57387 ^ t57387;
    wire t57389 = t57388 ^ t57388;
    wire t57390 = t57389 ^ t57389;
    wire t57391 = t57390 ^ t57390;
    wire t57392 = t57391 ^ t57391;
    wire t57393 = t57392 ^ t57392;
    wire t57394 = t57393 ^ t57393;
    wire t57395 = t57394 ^ t57394;
    wire t57396 = t57395 ^ t57395;
    wire t57397 = t57396 ^ t57396;
    wire t57398 = t57397 ^ t57397;
    wire t57399 = t57398 ^ t57398;
    wire t57400 = t57399 ^ t57399;
    wire t57401 = t57400 ^ t57400;
    wire t57402 = t57401 ^ t57401;
    wire t57403 = t57402 ^ t57402;
    wire t57404 = t57403 ^ t57403;
    wire t57405 = t57404 ^ t57404;
    wire t57406 = t57405 ^ t57405;
    wire t57407 = t57406 ^ t57406;
    wire t57408 = t57407 ^ t57407;
    wire t57409 = t57408 ^ t57408;
    wire t57410 = t57409 ^ t57409;
    wire t57411 = t57410 ^ t57410;
    wire t57412 = t57411 ^ t57411;
    wire t57413 = t57412 ^ t57412;
    wire t57414 = t57413 ^ t57413;
    wire t57415 = t57414 ^ t57414;
    wire t57416 = t57415 ^ t57415;
    wire t57417 = t57416 ^ t57416;
    wire t57418 = t57417 ^ t57417;
    wire t57419 = t57418 ^ t57418;
    wire t57420 = t57419 ^ t57419;
    wire t57421 = t57420 ^ t57420;
    wire t57422 = t57421 ^ t57421;
    wire t57423 = t57422 ^ t57422;
    wire t57424 = t57423 ^ t57423;
    wire t57425 = t57424 ^ t57424;
    wire t57426 = t57425 ^ t57425;
    wire t57427 = t57426 ^ t57426;
    wire t57428 = t57427 ^ t57427;
    wire t57429 = t57428 ^ t57428;
    wire t57430 = t57429 ^ t57429;
    wire t57431 = t57430 ^ t57430;
    wire t57432 = t57431 ^ t57431;
    wire t57433 = t57432 ^ t57432;
    wire t57434 = t57433 ^ t57433;
    wire t57435 = t57434 ^ t57434;
    wire t57436 = t57435 ^ t57435;
    wire t57437 = t57436 ^ t57436;
    wire t57438 = t57437 ^ t57437;
    wire t57439 = t57438 ^ t57438;
    wire t57440 = t57439 ^ t57439;
    wire t57441 = t57440 ^ t57440;
    wire t57442 = t57441 ^ t57441;
    wire t57443 = t57442 ^ t57442;
    wire t57444 = t57443 ^ t57443;
    wire t57445 = t57444 ^ t57444;
    wire t57446 = t57445 ^ t57445;
    wire t57447 = t57446 ^ t57446;
    wire t57448 = t57447 ^ t57447;
    wire t57449 = t57448 ^ t57448;
    wire t57450 = t57449 ^ t57449;
    wire t57451 = t57450 ^ t57450;
    wire t57452 = t57451 ^ t57451;
    wire t57453 = t57452 ^ t57452;
    wire t57454 = t57453 ^ t57453;
    wire t57455 = t57454 ^ t57454;
    wire t57456 = t57455 ^ t57455;
    wire t57457 = t57456 ^ t57456;
    wire t57458 = t57457 ^ t57457;
    wire t57459 = t57458 ^ t57458;
    wire t57460 = t57459 ^ t57459;
    wire t57461 = t57460 ^ t57460;
    wire t57462 = t57461 ^ t57461;
    wire t57463 = t57462 ^ t57462;
    wire t57464 = t57463 ^ t57463;
    wire t57465 = t57464 ^ t57464;
    wire t57466 = t57465 ^ t57465;
    wire t57467 = t57466 ^ t57466;
    wire t57468 = t57467 ^ t57467;
    wire t57469 = t57468 ^ t57468;
    wire t57470 = t57469 ^ t57469;
    wire t57471 = t57470 ^ t57470;
    wire t57472 = t57471 ^ t57471;
    wire t57473 = t57472 ^ t57472;
    wire t57474 = t57473 ^ t57473;
    wire t57475 = t57474 ^ t57474;
    wire t57476 = t57475 ^ t57475;
    wire t57477 = t57476 ^ t57476;
    wire t57478 = t57477 ^ t57477;
    wire t57479 = t57478 ^ t57478;
    wire t57480 = t57479 ^ t57479;
    wire t57481 = t57480 ^ t57480;
    wire t57482 = t57481 ^ t57481;
    wire t57483 = t57482 ^ t57482;
    wire t57484 = t57483 ^ t57483;
    wire t57485 = t57484 ^ t57484;
    wire t57486 = t57485 ^ t57485;
    wire t57487 = t57486 ^ t57486;
    wire t57488 = t57487 ^ t57487;
    wire t57489 = t57488 ^ t57488;
    wire t57490 = t57489 ^ t57489;
    wire t57491 = t57490 ^ t57490;
    wire t57492 = t57491 ^ t57491;
    wire t57493 = t57492 ^ t57492;
    wire t57494 = t57493 ^ t57493;
    wire t57495 = t57494 ^ t57494;
    wire t57496 = t57495 ^ t57495;
    wire t57497 = t57496 ^ t57496;
    wire t57498 = t57497 ^ t57497;
    wire t57499 = t57498 ^ t57498;
    wire t57500 = t57499 ^ t57499;
    wire t57501 = t57500 ^ t57500;
    wire t57502 = t57501 ^ t57501;
    wire t57503 = t57502 ^ t57502;
    wire t57504 = t57503 ^ t57503;
    wire t57505 = t57504 ^ t57504;
    wire t57506 = t57505 ^ t57505;
    wire t57507 = t57506 ^ t57506;
    wire t57508 = t57507 ^ t57507;
    wire t57509 = t57508 ^ t57508;
    wire t57510 = t57509 ^ t57509;
    wire t57511 = t57510 ^ t57510;
    wire t57512 = t57511 ^ t57511;
    wire t57513 = t57512 ^ t57512;
    wire t57514 = t57513 ^ t57513;
    wire t57515 = t57514 ^ t57514;
    wire t57516 = t57515 ^ t57515;
    wire t57517 = t57516 ^ t57516;
    wire t57518 = t57517 ^ t57517;
    wire t57519 = t57518 ^ t57518;
    wire t57520 = t57519 ^ t57519;
    wire t57521 = t57520 ^ t57520;
    wire t57522 = t57521 ^ t57521;
    wire t57523 = t57522 ^ t57522;
    wire t57524 = t57523 ^ t57523;
    wire t57525 = t57524 ^ t57524;
    wire t57526 = t57525 ^ t57525;
    wire t57527 = t57526 ^ t57526;
    wire t57528 = t57527 ^ t57527;
    wire t57529 = t57528 ^ t57528;
    wire t57530 = t57529 ^ t57529;
    wire t57531 = t57530 ^ t57530;
    wire t57532 = t57531 ^ t57531;
    wire t57533 = t57532 ^ t57532;
    wire t57534 = t57533 ^ t57533;
    wire t57535 = t57534 ^ t57534;
    wire t57536 = t57535 ^ t57535;
    wire t57537 = t57536 ^ t57536;
    wire t57538 = t57537 ^ t57537;
    wire t57539 = t57538 ^ t57538;
    wire t57540 = t57539 ^ t57539;
    wire t57541 = t57540 ^ t57540;
    wire t57542 = t57541 ^ t57541;
    wire t57543 = t57542 ^ t57542;
    wire t57544 = t57543 ^ t57543;
    wire t57545 = t57544 ^ t57544;
    wire t57546 = t57545 ^ t57545;
    wire t57547 = t57546 ^ t57546;
    wire t57548 = t57547 ^ t57547;
    wire t57549 = t57548 ^ t57548;
    wire t57550 = t57549 ^ t57549;
    wire t57551 = t57550 ^ t57550;
    wire t57552 = t57551 ^ t57551;
    wire t57553 = t57552 ^ t57552;
    wire t57554 = t57553 ^ t57553;
    wire t57555 = t57554 ^ t57554;
    wire t57556 = t57555 ^ t57555;
    wire t57557 = t57556 ^ t57556;
    wire t57558 = t57557 ^ t57557;
    wire t57559 = t57558 ^ t57558;
    wire t57560 = t57559 ^ t57559;
    wire t57561 = t57560 ^ t57560;
    wire t57562 = t57561 ^ t57561;
    wire t57563 = t57562 ^ t57562;
    wire t57564 = t57563 ^ t57563;
    wire t57565 = t57564 ^ t57564;
    wire t57566 = t57565 ^ t57565;
    wire t57567 = t57566 ^ t57566;
    wire t57568 = t57567 ^ t57567;
    wire t57569 = t57568 ^ t57568;
    wire t57570 = t57569 ^ t57569;
    wire t57571 = t57570 ^ t57570;
    wire t57572 = t57571 ^ t57571;
    wire t57573 = t57572 ^ t57572;
    wire t57574 = t57573 ^ t57573;
    wire t57575 = t57574 ^ t57574;
    wire t57576 = t57575 ^ t57575;
    wire t57577 = t57576 ^ t57576;
    wire t57578 = t57577 ^ t57577;
    wire t57579 = t57578 ^ t57578;
    wire t57580 = t57579 ^ t57579;
    wire t57581 = t57580 ^ t57580;
    wire t57582 = t57581 ^ t57581;
    wire t57583 = t57582 ^ t57582;
    wire t57584 = t57583 ^ t57583;
    wire t57585 = t57584 ^ t57584;
    wire t57586 = t57585 ^ t57585;
    wire t57587 = t57586 ^ t57586;
    wire t57588 = t57587 ^ t57587;
    wire t57589 = t57588 ^ t57588;
    wire t57590 = t57589 ^ t57589;
    wire t57591 = t57590 ^ t57590;
    wire t57592 = t57591 ^ t57591;
    wire t57593 = t57592 ^ t57592;
    wire t57594 = t57593 ^ t57593;
    wire t57595 = t57594 ^ t57594;
    wire t57596 = t57595 ^ t57595;
    wire t57597 = t57596 ^ t57596;
    wire t57598 = t57597 ^ t57597;
    wire t57599 = t57598 ^ t57598;
    wire t57600 = t57599 ^ t57599;
    wire t57601 = t57600 ^ t57600;
    wire t57602 = t57601 ^ t57601;
    wire t57603 = t57602 ^ t57602;
    wire t57604 = t57603 ^ t57603;
    wire t57605 = t57604 ^ t57604;
    wire t57606 = t57605 ^ t57605;
    wire t57607 = t57606 ^ t57606;
    wire t57608 = t57607 ^ t57607;
    wire t57609 = t57608 ^ t57608;
    wire t57610 = t57609 ^ t57609;
    wire t57611 = t57610 ^ t57610;
    wire t57612 = t57611 ^ t57611;
    wire t57613 = t57612 ^ t57612;
    wire t57614 = t57613 ^ t57613;
    wire t57615 = t57614 ^ t57614;
    wire t57616 = t57615 ^ t57615;
    wire t57617 = t57616 ^ t57616;
    wire t57618 = t57617 ^ t57617;
    wire t57619 = t57618 ^ t57618;
    wire t57620 = t57619 ^ t57619;
    wire t57621 = t57620 ^ t57620;
    wire t57622 = t57621 ^ t57621;
    wire t57623 = t57622 ^ t57622;
    wire t57624 = t57623 ^ t57623;
    wire t57625 = t57624 ^ t57624;
    wire t57626 = t57625 ^ t57625;
    wire t57627 = t57626 ^ t57626;
    wire t57628 = t57627 ^ t57627;
    wire t57629 = t57628 ^ t57628;
    wire t57630 = t57629 ^ t57629;
    wire t57631 = t57630 ^ t57630;
    wire t57632 = t57631 ^ t57631;
    wire t57633 = t57632 ^ t57632;
    wire t57634 = t57633 ^ t57633;
    wire t57635 = t57634 ^ t57634;
    wire t57636 = t57635 ^ t57635;
    wire t57637 = t57636 ^ t57636;
    wire t57638 = t57637 ^ t57637;
    wire t57639 = t57638 ^ t57638;
    wire t57640 = t57639 ^ t57639;
    wire t57641 = t57640 ^ t57640;
    wire t57642 = t57641 ^ t57641;
    wire t57643 = t57642 ^ t57642;
    wire t57644 = t57643 ^ t57643;
    wire t57645 = t57644 ^ t57644;
    wire t57646 = t57645 ^ t57645;
    wire t57647 = t57646 ^ t57646;
    wire t57648 = t57647 ^ t57647;
    wire t57649 = t57648 ^ t57648;
    wire t57650 = t57649 ^ t57649;
    wire t57651 = t57650 ^ t57650;
    wire t57652 = t57651 ^ t57651;
    wire t57653 = t57652 ^ t57652;
    wire t57654 = t57653 ^ t57653;
    wire t57655 = t57654 ^ t57654;
    wire t57656 = t57655 ^ t57655;
    wire t57657 = t57656 ^ t57656;
    wire t57658 = t57657 ^ t57657;
    wire t57659 = t57658 ^ t57658;
    wire t57660 = t57659 ^ t57659;
    wire t57661 = t57660 ^ t57660;
    wire t57662 = t57661 ^ t57661;
    wire t57663 = t57662 ^ t57662;
    wire t57664 = t57663 ^ t57663;
    wire t57665 = t57664 ^ t57664;
    wire t57666 = t57665 ^ t57665;
    wire t57667 = t57666 ^ t57666;
    wire t57668 = t57667 ^ t57667;
    wire t57669 = t57668 ^ t57668;
    wire t57670 = t57669 ^ t57669;
    wire t57671 = t57670 ^ t57670;
    wire t57672 = t57671 ^ t57671;
    wire t57673 = t57672 ^ t57672;
    wire t57674 = t57673 ^ t57673;
    wire t57675 = t57674 ^ t57674;
    wire t57676 = t57675 ^ t57675;
    wire t57677 = t57676 ^ t57676;
    wire t57678 = t57677 ^ t57677;
    wire t57679 = t57678 ^ t57678;
    wire t57680 = t57679 ^ t57679;
    wire t57681 = t57680 ^ t57680;
    wire t57682 = t57681 ^ t57681;
    wire t57683 = t57682 ^ t57682;
    wire t57684 = t57683 ^ t57683;
    wire t57685 = t57684 ^ t57684;
    wire t57686 = t57685 ^ t57685;
    wire t57687 = t57686 ^ t57686;
    wire t57688 = t57687 ^ t57687;
    wire t57689 = t57688 ^ t57688;
    wire t57690 = t57689 ^ t57689;
    wire t57691 = t57690 ^ t57690;
    wire t57692 = t57691 ^ t57691;
    wire t57693 = t57692 ^ t57692;
    wire t57694 = t57693 ^ t57693;
    wire t57695 = t57694 ^ t57694;
    wire t57696 = t57695 ^ t57695;
    wire t57697 = t57696 ^ t57696;
    wire t57698 = t57697 ^ t57697;
    wire t57699 = t57698 ^ t57698;
    wire t57700 = t57699 ^ t57699;
    wire t57701 = t57700 ^ t57700;
    wire t57702 = t57701 ^ t57701;
    wire t57703 = t57702 ^ t57702;
    wire t57704 = t57703 ^ t57703;
    wire t57705 = t57704 ^ t57704;
    wire t57706 = t57705 ^ t57705;
    wire t57707 = t57706 ^ t57706;
    wire t57708 = t57707 ^ t57707;
    wire t57709 = t57708 ^ t57708;
    wire t57710 = t57709 ^ t57709;
    wire t57711 = t57710 ^ t57710;
    wire t57712 = t57711 ^ t57711;
    wire t57713 = t57712 ^ t57712;
    wire t57714 = t57713 ^ t57713;
    wire t57715 = t57714 ^ t57714;
    wire t57716 = t57715 ^ t57715;
    wire t57717 = t57716 ^ t57716;
    wire t57718 = t57717 ^ t57717;
    wire t57719 = t57718 ^ t57718;
    wire t57720 = t57719 ^ t57719;
    wire t57721 = t57720 ^ t57720;
    wire t57722 = t57721 ^ t57721;
    wire t57723 = t57722 ^ t57722;
    wire t57724 = t57723 ^ t57723;
    wire t57725 = t57724 ^ t57724;
    wire t57726 = t57725 ^ t57725;
    wire t57727 = t57726 ^ t57726;
    wire t57728 = t57727 ^ t57727;
    wire t57729 = t57728 ^ t57728;
    wire t57730 = t57729 ^ t57729;
    wire t57731 = t57730 ^ t57730;
    wire t57732 = t57731 ^ t57731;
    wire t57733 = t57732 ^ t57732;
    wire t57734 = t57733 ^ t57733;
    wire t57735 = t57734 ^ t57734;
    wire t57736 = t57735 ^ t57735;
    wire t57737 = t57736 ^ t57736;
    wire t57738 = t57737 ^ t57737;
    wire t57739 = t57738 ^ t57738;
    wire t57740 = t57739 ^ t57739;
    wire t57741 = t57740 ^ t57740;
    wire t57742 = t57741 ^ t57741;
    wire t57743 = t57742 ^ t57742;
    wire t57744 = t57743 ^ t57743;
    wire t57745 = t57744 ^ t57744;
    wire t57746 = t57745 ^ t57745;
    wire t57747 = t57746 ^ t57746;
    wire t57748 = t57747 ^ t57747;
    wire t57749 = t57748 ^ t57748;
    wire t57750 = t57749 ^ t57749;
    wire t57751 = t57750 ^ t57750;
    wire t57752 = t57751 ^ t57751;
    wire t57753 = t57752 ^ t57752;
    wire t57754 = t57753 ^ t57753;
    wire t57755 = t57754 ^ t57754;
    wire t57756 = t57755 ^ t57755;
    wire t57757 = t57756 ^ t57756;
    wire t57758 = t57757 ^ t57757;
    wire t57759 = t57758 ^ t57758;
    wire t57760 = t57759 ^ t57759;
    wire t57761 = t57760 ^ t57760;
    wire t57762 = t57761 ^ t57761;
    wire t57763 = t57762 ^ t57762;
    wire t57764 = t57763 ^ t57763;
    wire t57765 = t57764 ^ t57764;
    wire t57766 = t57765 ^ t57765;
    wire t57767 = t57766 ^ t57766;
    wire t57768 = t57767 ^ t57767;
    wire t57769 = t57768 ^ t57768;
    wire t57770 = t57769 ^ t57769;
    wire t57771 = t57770 ^ t57770;
    wire t57772 = t57771 ^ t57771;
    wire t57773 = t57772 ^ t57772;
    wire t57774 = t57773 ^ t57773;
    wire t57775 = t57774 ^ t57774;
    wire t57776 = t57775 ^ t57775;
    wire t57777 = t57776 ^ t57776;
    wire t57778 = t57777 ^ t57777;
    wire t57779 = t57778 ^ t57778;
    wire t57780 = t57779 ^ t57779;
    wire t57781 = t57780 ^ t57780;
    wire t57782 = t57781 ^ t57781;
    wire t57783 = t57782 ^ t57782;
    wire t57784 = t57783 ^ t57783;
    wire t57785 = t57784 ^ t57784;
    wire t57786 = t57785 ^ t57785;
    wire t57787 = t57786 ^ t57786;
    wire t57788 = t57787 ^ t57787;
    wire t57789 = t57788 ^ t57788;
    wire t57790 = t57789 ^ t57789;
    wire t57791 = t57790 ^ t57790;
    wire t57792 = t57791 ^ t57791;
    wire t57793 = t57792 ^ t57792;
    wire t57794 = t57793 ^ t57793;
    wire t57795 = t57794 ^ t57794;
    wire t57796 = t57795 ^ t57795;
    wire t57797 = t57796 ^ t57796;
    wire t57798 = t57797 ^ t57797;
    wire t57799 = t57798 ^ t57798;
    wire t57800 = t57799 ^ t57799;
    wire t57801 = t57800 ^ t57800;
    wire t57802 = t57801 ^ t57801;
    wire t57803 = t57802 ^ t57802;
    wire t57804 = t57803 ^ t57803;
    wire t57805 = t57804 ^ t57804;
    wire t57806 = t57805 ^ t57805;
    wire t57807 = t57806 ^ t57806;
    wire t57808 = t57807 ^ t57807;
    wire t57809 = t57808 ^ t57808;
    wire t57810 = t57809 ^ t57809;
    wire t57811 = t57810 ^ t57810;
    wire t57812 = t57811 ^ t57811;
    wire t57813 = t57812 ^ t57812;
    wire t57814 = t57813 ^ t57813;
    wire t57815 = t57814 ^ t57814;
    wire t57816 = t57815 ^ t57815;
    wire t57817 = t57816 ^ t57816;
    wire t57818 = t57817 ^ t57817;
    wire t57819 = t57818 ^ t57818;
    wire t57820 = t57819 ^ t57819;
    wire t57821 = t57820 ^ t57820;
    wire t57822 = t57821 ^ t57821;
    wire t57823 = t57822 ^ t57822;
    wire t57824 = t57823 ^ t57823;
    wire t57825 = t57824 ^ t57824;
    wire t57826 = t57825 ^ t57825;
    wire t57827 = t57826 ^ t57826;
    wire t57828 = t57827 ^ t57827;
    wire t57829 = t57828 ^ t57828;
    wire t57830 = t57829 ^ t57829;
    wire t57831 = t57830 ^ t57830;
    wire t57832 = t57831 ^ t57831;
    wire t57833 = t57832 ^ t57832;
    wire t57834 = t57833 ^ t57833;
    wire t57835 = t57834 ^ t57834;
    wire t57836 = t57835 ^ t57835;
    wire t57837 = t57836 ^ t57836;
    wire t57838 = t57837 ^ t57837;
    wire t57839 = t57838 ^ t57838;
    wire t57840 = t57839 ^ t57839;
    wire t57841 = t57840 ^ t57840;
    wire t57842 = t57841 ^ t57841;
    wire t57843 = t57842 ^ t57842;
    wire t57844 = t57843 ^ t57843;
    wire t57845 = t57844 ^ t57844;
    wire t57846 = t57845 ^ t57845;
    wire t57847 = t57846 ^ t57846;
    wire t57848 = t57847 ^ t57847;
    wire t57849 = t57848 ^ t57848;
    wire t57850 = t57849 ^ t57849;
    wire t57851 = t57850 ^ t57850;
    wire t57852 = t57851 ^ t57851;
    wire t57853 = t57852 ^ t57852;
    wire t57854 = t57853 ^ t57853;
    wire t57855 = t57854 ^ t57854;
    wire t57856 = t57855 ^ t57855;
    wire t57857 = t57856 ^ t57856;
    wire t57858 = t57857 ^ t57857;
    wire t57859 = t57858 ^ t57858;
    wire t57860 = t57859 ^ t57859;
    wire t57861 = t57860 ^ t57860;
    wire t57862 = t57861 ^ t57861;
    wire t57863 = t57862 ^ t57862;
    wire t57864 = t57863 ^ t57863;
    wire t57865 = t57864 ^ t57864;
    wire t57866 = t57865 ^ t57865;
    wire t57867 = t57866 ^ t57866;
    wire t57868 = t57867 ^ t57867;
    wire t57869 = t57868 ^ t57868;
    wire t57870 = t57869 ^ t57869;
    wire t57871 = t57870 ^ t57870;
    wire t57872 = t57871 ^ t57871;
    wire t57873 = t57872 ^ t57872;
    wire t57874 = t57873 ^ t57873;
    wire t57875 = t57874 ^ t57874;
    wire t57876 = t57875 ^ t57875;
    wire t57877 = t57876 ^ t57876;
    wire t57878 = t57877 ^ t57877;
    wire t57879 = t57878 ^ t57878;
    wire t57880 = t57879 ^ t57879;
    wire t57881 = t57880 ^ t57880;
    wire t57882 = t57881 ^ t57881;
    wire t57883 = t57882 ^ t57882;
    wire t57884 = t57883 ^ t57883;
    wire t57885 = t57884 ^ t57884;
    wire t57886 = t57885 ^ t57885;
    wire t57887 = t57886 ^ t57886;
    wire t57888 = t57887 ^ t57887;
    wire t57889 = t57888 ^ t57888;
    wire t57890 = t57889 ^ t57889;
    wire t57891 = t57890 ^ t57890;
    wire t57892 = t57891 ^ t57891;
    wire t57893 = t57892 ^ t57892;
    wire t57894 = t57893 ^ t57893;
    wire t57895 = t57894 ^ t57894;
    wire t57896 = t57895 ^ t57895;
    wire t57897 = t57896 ^ t57896;
    wire t57898 = t57897 ^ t57897;
    wire t57899 = t57898 ^ t57898;
    wire t57900 = t57899 ^ t57899;
    wire t57901 = t57900 ^ t57900;
    wire t57902 = t57901 ^ t57901;
    wire t57903 = t57902 ^ t57902;
    wire t57904 = t57903 ^ t57903;
    wire t57905 = t57904 ^ t57904;
    wire t57906 = t57905 ^ t57905;
    wire t57907 = t57906 ^ t57906;
    wire t57908 = t57907 ^ t57907;
    wire t57909 = t57908 ^ t57908;
    wire t57910 = t57909 ^ t57909;
    wire t57911 = t57910 ^ t57910;
    wire t57912 = t57911 ^ t57911;
    wire t57913 = t57912 ^ t57912;
    wire t57914 = t57913 ^ t57913;
    wire t57915 = t57914 ^ t57914;
    wire t57916 = t57915 ^ t57915;
    wire t57917 = t57916 ^ t57916;
    wire t57918 = t57917 ^ t57917;
    wire t57919 = t57918 ^ t57918;
    wire t57920 = t57919 ^ t57919;
    wire t57921 = t57920 ^ t57920;
    wire t57922 = t57921 ^ t57921;
    wire t57923 = t57922 ^ t57922;
    wire t57924 = t57923 ^ t57923;
    wire t57925 = t57924 ^ t57924;
    wire t57926 = t57925 ^ t57925;
    wire t57927 = t57926 ^ t57926;
    wire t57928 = t57927 ^ t57927;
    wire t57929 = t57928 ^ t57928;
    wire t57930 = t57929 ^ t57929;
    wire t57931 = t57930 ^ t57930;
    wire t57932 = t57931 ^ t57931;
    wire t57933 = t57932 ^ t57932;
    wire t57934 = t57933 ^ t57933;
    wire t57935 = t57934 ^ t57934;
    wire t57936 = t57935 ^ t57935;
    wire t57937 = t57936 ^ t57936;
    wire t57938 = t57937 ^ t57937;
    wire t57939 = t57938 ^ t57938;
    wire t57940 = t57939 ^ t57939;
    wire t57941 = t57940 ^ t57940;
    wire t57942 = t57941 ^ t57941;
    wire t57943 = t57942 ^ t57942;
    wire t57944 = t57943 ^ t57943;
    wire t57945 = t57944 ^ t57944;
    wire t57946 = t57945 ^ t57945;
    wire t57947 = t57946 ^ t57946;
    wire t57948 = t57947 ^ t57947;
    wire t57949 = t57948 ^ t57948;
    wire t57950 = t57949 ^ t57949;
    wire t57951 = t57950 ^ t57950;
    wire t57952 = t57951 ^ t57951;
    wire t57953 = t57952 ^ t57952;
    wire t57954 = t57953 ^ t57953;
    wire t57955 = t57954 ^ t57954;
    wire t57956 = t57955 ^ t57955;
    wire t57957 = t57956 ^ t57956;
    wire t57958 = t57957 ^ t57957;
    wire t57959 = t57958 ^ t57958;
    wire t57960 = t57959 ^ t57959;
    wire t57961 = t57960 ^ t57960;
    wire t57962 = t57961 ^ t57961;
    wire t57963 = t57962 ^ t57962;
    wire t57964 = t57963 ^ t57963;
    wire t57965 = t57964 ^ t57964;
    wire t57966 = t57965 ^ t57965;
    wire t57967 = t57966 ^ t57966;
    wire t57968 = t57967 ^ t57967;
    wire t57969 = t57968 ^ t57968;
    wire t57970 = t57969 ^ t57969;
    wire t57971 = t57970 ^ t57970;
    wire t57972 = t57971 ^ t57971;
    wire t57973 = t57972 ^ t57972;
    wire t57974 = t57973 ^ t57973;
    wire t57975 = t57974 ^ t57974;
    wire t57976 = t57975 ^ t57975;
    wire t57977 = t57976 ^ t57976;
    wire t57978 = t57977 ^ t57977;
    wire t57979 = t57978 ^ t57978;
    wire t57980 = t57979 ^ t57979;
    wire t57981 = t57980 ^ t57980;
    wire t57982 = t57981 ^ t57981;
    wire t57983 = t57982 ^ t57982;
    wire t57984 = t57983 ^ t57983;
    wire t57985 = t57984 ^ t57984;
    wire t57986 = t57985 ^ t57985;
    wire t57987 = t57986 ^ t57986;
    wire t57988 = t57987 ^ t57987;
    wire t57989 = t57988 ^ t57988;
    wire t57990 = t57989 ^ t57989;
    wire t57991 = t57990 ^ t57990;
    wire t57992 = t57991 ^ t57991;
    wire t57993 = t57992 ^ t57992;
    wire t57994 = t57993 ^ t57993;
    wire t57995 = t57994 ^ t57994;
    wire t57996 = t57995 ^ t57995;
    wire t57997 = t57996 ^ t57996;
    wire t57998 = t57997 ^ t57997;
    wire t57999 = t57998 ^ t57998;
    wire t58000 = t57999 ^ t57999;
    wire t58001 = t58000 ^ t58000;
    wire t58002 = t58001 ^ t58001;
    wire t58003 = t58002 ^ t58002;
    wire t58004 = t58003 ^ t58003;
    wire t58005 = t58004 ^ t58004;
    wire t58006 = t58005 ^ t58005;
    wire t58007 = t58006 ^ t58006;
    wire t58008 = t58007 ^ t58007;
    wire t58009 = t58008 ^ t58008;
    wire t58010 = t58009 ^ t58009;
    wire t58011 = t58010 ^ t58010;
    wire t58012 = t58011 ^ t58011;
    wire t58013 = t58012 ^ t58012;
    wire t58014 = t58013 ^ t58013;
    wire t58015 = t58014 ^ t58014;
    wire t58016 = t58015 ^ t58015;
    wire t58017 = t58016 ^ t58016;
    wire t58018 = t58017 ^ t58017;
    wire t58019 = t58018 ^ t58018;
    wire t58020 = t58019 ^ t58019;
    wire t58021 = t58020 ^ t58020;
    wire t58022 = t58021 ^ t58021;
    wire t58023 = t58022 ^ t58022;
    wire t58024 = t58023 ^ t58023;
    wire t58025 = t58024 ^ t58024;
    wire t58026 = t58025 ^ t58025;
    wire t58027 = t58026 ^ t58026;
    wire t58028 = t58027 ^ t58027;
    wire t58029 = t58028 ^ t58028;
    wire t58030 = t58029 ^ t58029;
    wire t58031 = t58030 ^ t58030;
    wire t58032 = t58031 ^ t58031;
    wire t58033 = t58032 ^ t58032;
    wire t58034 = t58033 ^ t58033;
    wire t58035 = t58034 ^ t58034;
    wire t58036 = t58035 ^ t58035;
    wire t58037 = t58036 ^ t58036;
    wire t58038 = t58037 ^ t58037;
    wire t58039 = t58038 ^ t58038;
    wire t58040 = t58039 ^ t58039;
    wire t58041 = t58040 ^ t58040;
    wire t58042 = t58041 ^ t58041;
    wire t58043 = t58042 ^ t58042;
    wire t58044 = t58043 ^ t58043;
    wire t58045 = t58044 ^ t58044;
    wire t58046 = t58045 ^ t58045;
    wire t58047 = t58046 ^ t58046;
    wire t58048 = t58047 ^ t58047;
    wire t58049 = t58048 ^ t58048;
    wire t58050 = t58049 ^ t58049;
    wire t58051 = t58050 ^ t58050;
    wire t58052 = t58051 ^ t58051;
    wire t58053 = t58052 ^ t58052;
    wire t58054 = t58053 ^ t58053;
    wire t58055 = t58054 ^ t58054;
    wire t58056 = t58055 ^ t58055;
    wire t58057 = t58056 ^ t58056;
    wire t58058 = t58057 ^ t58057;
    wire t58059 = t58058 ^ t58058;
    wire t58060 = t58059 ^ t58059;
    wire t58061 = t58060 ^ t58060;
    wire t58062 = t58061 ^ t58061;
    wire t58063 = t58062 ^ t58062;
    wire t58064 = t58063 ^ t58063;
    wire t58065 = t58064 ^ t58064;
    wire t58066 = t58065 ^ t58065;
    wire t58067 = t58066 ^ t58066;
    wire t58068 = t58067 ^ t58067;
    wire t58069 = t58068 ^ t58068;
    wire t58070 = t58069 ^ t58069;
    wire t58071 = t58070 ^ t58070;
    wire t58072 = t58071 ^ t58071;
    wire t58073 = t58072 ^ t58072;
    wire t58074 = t58073 ^ t58073;
    wire t58075 = t58074 ^ t58074;
    wire t58076 = t58075 ^ t58075;
    wire t58077 = t58076 ^ t58076;
    wire t58078 = t58077 ^ t58077;
    wire t58079 = t58078 ^ t58078;
    wire t58080 = t58079 ^ t58079;
    wire t58081 = t58080 ^ t58080;
    wire t58082 = t58081 ^ t58081;
    wire t58083 = t58082 ^ t58082;
    wire t58084 = t58083 ^ t58083;
    wire t58085 = t58084 ^ t58084;
    wire t58086 = t58085 ^ t58085;
    wire t58087 = t58086 ^ t58086;
    wire t58088 = t58087 ^ t58087;
    wire t58089 = t58088 ^ t58088;
    wire t58090 = t58089 ^ t58089;
    wire t58091 = t58090 ^ t58090;
    wire t58092 = t58091 ^ t58091;
    wire t58093 = t58092 ^ t58092;
    wire t58094 = t58093 ^ t58093;
    wire t58095 = t58094 ^ t58094;
    wire t58096 = t58095 ^ t58095;
    wire t58097 = t58096 ^ t58096;
    wire t58098 = t58097 ^ t58097;
    wire t58099 = t58098 ^ t58098;
    wire t58100 = t58099 ^ t58099;
    wire t58101 = t58100 ^ t58100;
    wire t58102 = t58101 ^ t58101;
    wire t58103 = t58102 ^ t58102;
    wire t58104 = t58103 ^ t58103;
    wire t58105 = t58104 ^ t58104;
    wire t58106 = t58105 ^ t58105;
    wire t58107 = t58106 ^ t58106;
    wire t58108 = t58107 ^ t58107;
    wire t58109 = t58108 ^ t58108;
    wire t58110 = t58109 ^ t58109;
    wire t58111 = t58110 ^ t58110;
    wire t58112 = t58111 ^ t58111;
    wire t58113 = t58112 ^ t58112;
    wire t58114 = t58113 ^ t58113;
    wire t58115 = t58114 ^ t58114;
    wire t58116 = t58115 ^ t58115;
    wire t58117 = t58116 ^ t58116;
    wire t58118 = t58117 ^ t58117;
    wire t58119 = t58118 ^ t58118;
    wire t58120 = t58119 ^ t58119;
    wire t58121 = t58120 ^ t58120;
    wire t58122 = t58121 ^ t58121;
    wire t58123 = t58122 ^ t58122;
    wire t58124 = t58123 ^ t58123;
    wire t58125 = t58124 ^ t58124;
    wire t58126 = t58125 ^ t58125;
    wire t58127 = t58126 ^ t58126;
    wire t58128 = t58127 ^ t58127;
    wire t58129 = t58128 ^ t58128;
    wire t58130 = t58129 ^ t58129;
    wire t58131 = t58130 ^ t58130;
    wire t58132 = t58131 ^ t58131;
    wire t58133 = t58132 ^ t58132;
    wire t58134 = t58133 ^ t58133;
    wire t58135 = t58134 ^ t58134;
    wire t58136 = t58135 ^ t58135;
    wire t58137 = t58136 ^ t58136;
    wire t58138 = t58137 ^ t58137;
    wire t58139 = t58138 ^ t58138;
    wire t58140 = t58139 ^ t58139;
    wire t58141 = t58140 ^ t58140;
    wire t58142 = t58141 ^ t58141;
    wire t58143 = t58142 ^ t58142;
    wire t58144 = t58143 ^ t58143;
    wire t58145 = t58144 ^ t58144;
    wire t58146 = t58145 ^ t58145;
    wire t58147 = t58146 ^ t58146;
    wire t58148 = t58147 ^ t58147;
    wire t58149 = t58148 ^ t58148;
    wire t58150 = t58149 ^ t58149;
    wire t58151 = t58150 ^ t58150;
    wire t58152 = t58151 ^ t58151;
    wire t58153 = t58152 ^ t58152;
    wire t58154 = t58153 ^ t58153;
    wire t58155 = t58154 ^ t58154;
    wire t58156 = t58155 ^ t58155;
    wire t58157 = t58156 ^ t58156;
    wire t58158 = t58157 ^ t58157;
    wire t58159 = t58158 ^ t58158;
    wire t58160 = t58159 ^ t58159;
    wire t58161 = t58160 ^ t58160;
    wire t58162 = t58161 ^ t58161;
    wire t58163 = t58162 ^ t58162;
    wire t58164 = t58163 ^ t58163;
    wire t58165 = t58164 ^ t58164;
    wire t58166 = t58165 ^ t58165;
    wire t58167 = t58166 ^ t58166;
    wire t58168 = t58167 ^ t58167;
    wire t58169 = t58168 ^ t58168;
    wire t58170 = t58169 ^ t58169;
    wire t58171 = t58170 ^ t58170;
    wire t58172 = t58171 ^ t58171;
    wire t58173 = t58172 ^ t58172;
    wire t58174 = t58173 ^ t58173;
    wire t58175 = t58174 ^ t58174;
    wire t58176 = t58175 ^ t58175;
    wire t58177 = t58176 ^ t58176;
    wire t58178 = t58177 ^ t58177;
    wire t58179 = t58178 ^ t58178;
    wire t58180 = t58179 ^ t58179;
    wire t58181 = t58180 ^ t58180;
    wire t58182 = t58181 ^ t58181;
    wire t58183 = t58182 ^ t58182;
    wire t58184 = t58183 ^ t58183;
    wire t58185 = t58184 ^ t58184;
    wire t58186 = t58185 ^ t58185;
    wire t58187 = t58186 ^ t58186;
    wire t58188 = t58187 ^ t58187;
    wire t58189 = t58188 ^ t58188;
    wire t58190 = t58189 ^ t58189;
    wire t58191 = t58190 ^ t58190;
    wire t58192 = t58191 ^ t58191;
    wire t58193 = t58192 ^ t58192;
    wire t58194 = t58193 ^ t58193;
    wire t58195 = t58194 ^ t58194;
    wire t58196 = t58195 ^ t58195;
    wire t58197 = t58196 ^ t58196;
    wire t58198 = t58197 ^ t58197;
    wire t58199 = t58198 ^ t58198;
    wire t58200 = t58199 ^ t58199;
    wire t58201 = t58200 ^ t58200;
    wire t58202 = t58201 ^ t58201;
    wire t58203 = t58202 ^ t58202;
    wire t58204 = t58203 ^ t58203;
    wire t58205 = t58204 ^ t58204;
    wire t58206 = t58205 ^ t58205;
    wire t58207 = t58206 ^ t58206;
    wire t58208 = t58207 ^ t58207;
    wire t58209 = t58208 ^ t58208;
    wire t58210 = t58209 ^ t58209;
    wire t58211 = t58210 ^ t58210;
    wire t58212 = t58211 ^ t58211;
    wire t58213 = t58212 ^ t58212;
    wire t58214 = t58213 ^ t58213;
    wire t58215 = t58214 ^ t58214;
    wire t58216 = t58215 ^ t58215;
    wire t58217 = t58216 ^ t58216;
    wire t58218 = t58217 ^ t58217;
    wire t58219 = t58218 ^ t58218;
    wire t58220 = t58219 ^ t58219;
    wire t58221 = t58220 ^ t58220;
    wire t58222 = t58221 ^ t58221;
    wire t58223 = t58222 ^ t58222;
    wire t58224 = t58223 ^ t58223;
    wire t58225 = t58224 ^ t58224;
    wire t58226 = t58225 ^ t58225;
    wire t58227 = t58226 ^ t58226;
    wire t58228 = t58227 ^ t58227;
    wire t58229 = t58228 ^ t58228;
    wire t58230 = t58229 ^ t58229;
    wire t58231 = t58230 ^ t58230;
    wire t58232 = t58231 ^ t58231;
    wire t58233 = t58232 ^ t58232;
    wire t58234 = t58233 ^ t58233;
    wire t58235 = t58234 ^ t58234;
    wire t58236 = t58235 ^ t58235;
    wire t58237 = t58236 ^ t58236;
    wire t58238 = t58237 ^ t58237;
    wire t58239 = t58238 ^ t58238;
    wire t58240 = t58239 ^ t58239;
    wire t58241 = t58240 ^ t58240;
    wire t58242 = t58241 ^ t58241;
    wire t58243 = t58242 ^ t58242;
    wire t58244 = t58243 ^ t58243;
    wire t58245 = t58244 ^ t58244;
    wire t58246 = t58245 ^ t58245;
    wire t58247 = t58246 ^ t58246;
    wire t58248 = t58247 ^ t58247;
    wire t58249 = t58248 ^ t58248;
    wire t58250 = t58249 ^ t58249;
    wire t58251 = t58250 ^ t58250;
    wire t58252 = t58251 ^ t58251;
    wire t58253 = t58252 ^ t58252;
    wire t58254 = t58253 ^ t58253;
    wire t58255 = t58254 ^ t58254;
    wire t58256 = t58255 ^ t58255;
    wire t58257 = t58256 ^ t58256;
    wire t58258 = t58257 ^ t58257;
    wire t58259 = t58258 ^ t58258;
    wire t58260 = t58259 ^ t58259;
    wire t58261 = t58260 ^ t58260;
    wire t58262 = t58261 ^ t58261;
    wire t58263 = t58262 ^ t58262;
    wire t58264 = t58263 ^ t58263;
    wire t58265 = t58264 ^ t58264;
    wire t58266 = t58265 ^ t58265;
    wire t58267 = t58266 ^ t58266;
    wire t58268 = t58267 ^ t58267;
    wire t58269 = t58268 ^ t58268;
    wire t58270 = t58269 ^ t58269;
    wire t58271 = t58270 ^ t58270;
    wire t58272 = t58271 ^ t58271;
    wire t58273 = t58272 ^ t58272;
    wire t58274 = t58273 ^ t58273;
    wire t58275 = t58274 ^ t58274;
    wire t58276 = t58275 ^ t58275;
    wire t58277 = t58276 ^ t58276;
    wire t58278 = t58277 ^ t58277;
    wire t58279 = t58278 ^ t58278;
    wire t58280 = t58279 ^ t58279;
    wire t58281 = t58280 ^ t58280;
    wire t58282 = t58281 ^ t58281;
    wire t58283 = t58282 ^ t58282;
    wire t58284 = t58283 ^ t58283;
    wire t58285 = t58284 ^ t58284;
    wire t58286 = t58285 ^ t58285;
    wire t58287 = t58286 ^ t58286;
    wire t58288 = t58287 ^ t58287;
    wire t58289 = t58288 ^ t58288;
    wire t58290 = t58289 ^ t58289;
    wire t58291 = t58290 ^ t58290;
    wire t58292 = t58291 ^ t58291;
    wire t58293 = t58292 ^ t58292;
    wire t58294 = t58293 ^ t58293;
    wire t58295 = t58294 ^ t58294;
    wire t58296 = t58295 ^ t58295;
    wire t58297 = t58296 ^ t58296;
    wire t58298 = t58297 ^ t58297;
    wire t58299 = t58298 ^ t58298;
    wire t58300 = t58299 ^ t58299;
    wire t58301 = t58300 ^ t58300;
    wire t58302 = t58301 ^ t58301;
    wire t58303 = t58302 ^ t58302;
    wire t58304 = t58303 ^ t58303;
    wire t58305 = t58304 ^ t58304;
    wire t58306 = t58305 ^ t58305;
    wire t58307 = t58306 ^ t58306;
    wire t58308 = t58307 ^ t58307;
    wire t58309 = t58308 ^ t58308;
    wire t58310 = t58309 ^ t58309;
    wire t58311 = t58310 ^ t58310;
    wire t58312 = t58311 ^ t58311;
    wire t58313 = t58312 ^ t58312;
    wire t58314 = t58313 ^ t58313;
    wire t58315 = t58314 ^ t58314;
    wire t58316 = t58315 ^ t58315;
    wire t58317 = t58316 ^ t58316;
    wire t58318 = t58317 ^ t58317;
    wire t58319 = t58318 ^ t58318;
    wire t58320 = t58319 ^ t58319;
    wire t58321 = t58320 ^ t58320;
    wire t58322 = t58321 ^ t58321;
    wire t58323 = t58322 ^ t58322;
    wire t58324 = t58323 ^ t58323;
    wire t58325 = t58324 ^ t58324;
    wire t58326 = t58325 ^ t58325;
    wire t58327 = t58326 ^ t58326;
    wire t58328 = t58327 ^ t58327;
    wire t58329 = t58328 ^ t58328;
    wire t58330 = t58329 ^ t58329;
    wire t58331 = t58330 ^ t58330;
    wire t58332 = t58331 ^ t58331;
    wire t58333 = t58332 ^ t58332;
    wire t58334 = t58333 ^ t58333;
    wire t58335 = t58334 ^ t58334;
    wire t58336 = t58335 ^ t58335;
    wire t58337 = t58336 ^ t58336;
    wire t58338 = t58337 ^ t58337;
    wire t58339 = t58338 ^ t58338;
    wire t58340 = t58339 ^ t58339;
    wire t58341 = t58340 ^ t58340;
    wire t58342 = t58341 ^ t58341;
    wire t58343 = t58342 ^ t58342;
    wire t58344 = t58343 ^ t58343;
    wire t58345 = t58344 ^ t58344;
    wire t58346 = t58345 ^ t58345;
    wire t58347 = t58346 ^ t58346;
    wire t58348 = t58347 ^ t58347;
    wire t58349 = t58348 ^ t58348;
    wire t58350 = t58349 ^ t58349;
    wire t58351 = t58350 ^ t58350;
    wire t58352 = t58351 ^ t58351;
    wire t58353 = t58352 ^ t58352;
    wire t58354 = t58353 ^ t58353;
    wire t58355 = t58354 ^ t58354;
    wire t58356 = t58355 ^ t58355;
    wire t58357 = t58356 ^ t58356;
    wire t58358 = t58357 ^ t58357;
    wire t58359 = t58358 ^ t58358;
    wire t58360 = t58359 ^ t58359;
    wire t58361 = t58360 ^ t58360;
    wire t58362 = t58361 ^ t58361;
    wire t58363 = t58362 ^ t58362;
    wire t58364 = t58363 ^ t58363;
    wire t58365 = t58364 ^ t58364;
    wire t58366 = t58365 ^ t58365;
    wire t58367 = t58366 ^ t58366;
    wire t58368 = t58367 ^ t58367;
    wire t58369 = t58368 ^ t58368;
    wire t58370 = t58369 ^ t58369;
    wire t58371 = t58370 ^ t58370;
    wire t58372 = t58371 ^ t58371;
    wire t58373 = t58372 ^ t58372;
    wire t58374 = t58373 ^ t58373;
    wire t58375 = t58374 ^ t58374;
    wire t58376 = t58375 ^ t58375;
    wire t58377 = t58376 ^ t58376;
    wire t58378 = t58377 ^ t58377;
    wire t58379 = t58378 ^ t58378;
    wire t58380 = t58379 ^ t58379;
    wire t58381 = t58380 ^ t58380;
    wire t58382 = t58381 ^ t58381;
    wire t58383 = t58382 ^ t58382;
    wire t58384 = t58383 ^ t58383;
    wire t58385 = t58384 ^ t58384;
    wire t58386 = t58385 ^ t58385;
    wire t58387 = t58386 ^ t58386;
    wire t58388 = t58387 ^ t58387;
    wire t58389 = t58388 ^ t58388;
    wire t58390 = t58389 ^ t58389;
    wire t58391 = t58390 ^ t58390;
    wire t58392 = t58391 ^ t58391;
    wire t58393 = t58392 ^ t58392;
    wire t58394 = t58393 ^ t58393;
    wire t58395 = t58394 ^ t58394;
    wire t58396 = t58395 ^ t58395;
    wire t58397 = t58396 ^ t58396;
    wire t58398 = t58397 ^ t58397;
    wire t58399 = t58398 ^ t58398;
    wire t58400 = t58399 ^ t58399;
    wire t58401 = t58400 ^ t58400;
    wire t58402 = t58401 ^ t58401;
    wire t58403 = t58402 ^ t58402;
    wire t58404 = t58403 ^ t58403;
    wire t58405 = t58404 ^ t58404;
    wire t58406 = t58405 ^ t58405;
    wire t58407 = t58406 ^ t58406;
    wire t58408 = t58407 ^ t58407;
    wire t58409 = t58408 ^ t58408;
    wire t58410 = t58409 ^ t58409;
    wire t58411 = t58410 ^ t58410;
    wire t58412 = t58411 ^ t58411;
    wire t58413 = t58412 ^ t58412;
    wire t58414 = t58413 ^ t58413;
    wire t58415 = t58414 ^ t58414;
    wire t58416 = t58415 ^ t58415;
    wire t58417 = t58416 ^ t58416;
    wire t58418 = t58417 ^ t58417;
    wire t58419 = t58418 ^ t58418;
    wire t58420 = t58419 ^ t58419;
    wire t58421 = t58420 ^ t58420;
    wire t58422 = t58421 ^ t58421;
    wire t58423 = t58422 ^ t58422;
    wire t58424 = t58423 ^ t58423;
    wire t58425 = t58424 ^ t58424;
    wire t58426 = t58425 ^ t58425;
    wire t58427 = t58426 ^ t58426;
    wire t58428 = t58427 ^ t58427;
    wire t58429 = t58428 ^ t58428;
    wire t58430 = t58429 ^ t58429;
    wire t58431 = t58430 ^ t58430;
    wire t58432 = t58431 ^ t58431;
    wire t58433 = t58432 ^ t58432;
    wire t58434 = t58433 ^ t58433;
    wire t58435 = t58434 ^ t58434;
    wire t58436 = t58435 ^ t58435;
    wire t58437 = t58436 ^ t58436;
    wire t58438 = t58437 ^ t58437;
    wire t58439 = t58438 ^ t58438;
    wire t58440 = t58439 ^ t58439;
    wire t58441 = t58440 ^ t58440;
    wire t58442 = t58441 ^ t58441;
    wire t58443 = t58442 ^ t58442;
    wire t58444 = t58443 ^ t58443;
    wire t58445 = t58444 ^ t58444;
    wire t58446 = t58445 ^ t58445;
    wire t58447 = t58446 ^ t58446;
    wire t58448 = t58447 ^ t58447;
    wire t58449 = t58448 ^ t58448;
    wire t58450 = t58449 ^ t58449;
    wire t58451 = t58450 ^ t58450;
    wire t58452 = t58451 ^ t58451;
    wire t58453 = t58452 ^ t58452;
    wire t58454 = t58453 ^ t58453;
    wire t58455 = t58454 ^ t58454;
    wire t58456 = t58455 ^ t58455;
    wire t58457 = t58456 ^ t58456;
    wire t58458 = t58457 ^ t58457;
    wire t58459 = t58458 ^ t58458;
    wire t58460 = t58459 ^ t58459;
    wire t58461 = t58460 ^ t58460;
    wire t58462 = t58461 ^ t58461;
    wire t58463 = t58462 ^ t58462;
    wire t58464 = t58463 ^ t58463;
    wire t58465 = t58464 ^ t58464;
    wire t58466 = t58465 ^ t58465;
    wire t58467 = t58466 ^ t58466;
    wire t58468 = t58467 ^ t58467;
    wire t58469 = t58468 ^ t58468;
    wire t58470 = t58469 ^ t58469;
    wire t58471 = t58470 ^ t58470;
    wire t58472 = t58471 ^ t58471;
    wire t58473 = t58472 ^ t58472;
    wire t58474 = t58473 ^ t58473;
    wire t58475 = t58474 ^ t58474;
    wire t58476 = t58475 ^ t58475;
    wire t58477 = t58476 ^ t58476;
    wire t58478 = t58477 ^ t58477;
    wire t58479 = t58478 ^ t58478;
    wire t58480 = t58479 ^ t58479;
    wire t58481 = t58480 ^ t58480;
    wire t58482 = t58481 ^ t58481;
    wire t58483 = t58482 ^ t58482;
    wire t58484 = t58483 ^ t58483;
    wire t58485 = t58484 ^ t58484;
    wire t58486 = t58485 ^ t58485;
    wire t58487 = t58486 ^ t58486;
    wire t58488 = t58487 ^ t58487;
    wire t58489 = t58488 ^ t58488;
    wire t58490 = t58489 ^ t58489;
    wire t58491 = t58490 ^ t58490;
    wire t58492 = t58491 ^ t58491;
    wire t58493 = t58492 ^ t58492;
    wire t58494 = t58493 ^ t58493;
    wire t58495 = t58494 ^ t58494;
    wire t58496 = t58495 ^ t58495;
    wire t58497 = t58496 ^ t58496;
    wire t58498 = t58497 ^ t58497;
    wire t58499 = t58498 ^ t58498;
    wire t58500 = t58499 ^ t58499;
    wire t58501 = t58500 ^ t58500;
    wire t58502 = t58501 ^ t58501;
    wire t58503 = t58502 ^ t58502;
    wire t58504 = t58503 ^ t58503;
    wire t58505 = t58504 ^ t58504;
    wire t58506 = t58505 ^ t58505;
    wire t58507 = t58506 ^ t58506;
    wire t58508 = t58507 ^ t58507;
    wire t58509 = t58508 ^ t58508;
    wire t58510 = t58509 ^ t58509;
    wire t58511 = t58510 ^ t58510;
    wire t58512 = t58511 ^ t58511;
    wire t58513 = t58512 ^ t58512;
    wire t58514 = t58513 ^ t58513;
    wire t58515 = t58514 ^ t58514;
    wire t58516 = t58515 ^ t58515;
    wire t58517 = t58516 ^ t58516;
    wire t58518 = t58517 ^ t58517;
    wire t58519 = t58518 ^ t58518;
    wire t58520 = t58519 ^ t58519;
    wire t58521 = t58520 ^ t58520;
    wire t58522 = t58521 ^ t58521;
    wire t58523 = t58522 ^ t58522;
    wire t58524 = t58523 ^ t58523;
    wire t58525 = t58524 ^ t58524;
    wire t58526 = t58525 ^ t58525;
    wire t58527 = t58526 ^ t58526;
    wire t58528 = t58527 ^ t58527;
    wire t58529 = t58528 ^ t58528;
    wire t58530 = t58529 ^ t58529;
    wire t58531 = t58530 ^ t58530;
    wire t58532 = t58531 ^ t58531;
    wire t58533 = t58532 ^ t58532;
    wire t58534 = t58533 ^ t58533;
    wire t58535 = t58534 ^ t58534;
    wire t58536 = t58535 ^ t58535;
    wire t58537 = t58536 ^ t58536;
    wire t58538 = t58537 ^ t58537;
    wire t58539 = t58538 ^ t58538;
    wire t58540 = t58539 ^ t58539;
    wire t58541 = t58540 ^ t58540;
    wire t58542 = t58541 ^ t58541;
    wire t58543 = t58542 ^ t58542;
    wire t58544 = t58543 ^ t58543;
    wire t58545 = t58544 ^ t58544;
    wire t58546 = t58545 ^ t58545;
    wire t58547 = t58546 ^ t58546;
    wire t58548 = t58547 ^ t58547;
    wire t58549 = t58548 ^ t58548;
    wire t58550 = t58549 ^ t58549;
    wire t58551 = t58550 ^ t58550;
    wire t58552 = t58551 ^ t58551;
    wire t58553 = t58552 ^ t58552;
    wire t58554 = t58553 ^ t58553;
    wire t58555 = t58554 ^ t58554;
    wire t58556 = t58555 ^ t58555;
    wire t58557 = t58556 ^ t58556;
    wire t58558 = t58557 ^ t58557;
    wire t58559 = t58558 ^ t58558;
    wire t58560 = t58559 ^ t58559;
    wire t58561 = t58560 ^ t58560;
    wire t58562 = t58561 ^ t58561;
    wire t58563 = t58562 ^ t58562;
    wire t58564 = t58563 ^ t58563;
    wire t58565 = t58564 ^ t58564;
    wire t58566 = t58565 ^ t58565;
    wire t58567 = t58566 ^ t58566;
    wire t58568 = t58567 ^ t58567;
    wire t58569 = t58568 ^ t58568;
    wire t58570 = t58569 ^ t58569;
    wire t58571 = t58570 ^ t58570;
    wire t58572 = t58571 ^ t58571;
    wire t58573 = t58572 ^ t58572;
    wire t58574 = t58573 ^ t58573;
    wire t58575 = t58574 ^ t58574;
    wire t58576 = t58575 ^ t58575;
    wire t58577 = t58576 ^ t58576;
    wire t58578 = t58577 ^ t58577;
    wire t58579 = t58578 ^ t58578;
    wire t58580 = t58579 ^ t58579;
    wire t58581 = t58580 ^ t58580;
    wire t58582 = t58581 ^ t58581;
    wire t58583 = t58582 ^ t58582;
    wire t58584 = t58583 ^ t58583;
    wire t58585 = t58584 ^ t58584;
    wire t58586 = t58585 ^ t58585;
    wire t58587 = t58586 ^ t58586;
    wire t58588 = t58587 ^ t58587;
    wire t58589 = t58588 ^ t58588;
    wire t58590 = t58589 ^ t58589;
    wire t58591 = t58590 ^ t58590;
    wire t58592 = t58591 ^ t58591;
    wire t58593 = t58592 ^ t58592;
    wire t58594 = t58593 ^ t58593;
    wire t58595 = t58594 ^ t58594;
    wire t58596 = t58595 ^ t58595;
    wire t58597 = t58596 ^ t58596;
    wire t58598 = t58597 ^ t58597;
    wire t58599 = t58598 ^ t58598;
    wire t58600 = t58599 ^ t58599;
    wire t58601 = t58600 ^ t58600;
    wire t58602 = t58601 ^ t58601;
    wire t58603 = t58602 ^ t58602;
    wire t58604 = t58603 ^ t58603;
    wire t58605 = t58604 ^ t58604;
    wire t58606 = t58605 ^ t58605;
    wire t58607 = t58606 ^ t58606;
    wire t58608 = t58607 ^ t58607;
    wire t58609 = t58608 ^ t58608;
    wire t58610 = t58609 ^ t58609;
    wire t58611 = t58610 ^ t58610;
    wire t58612 = t58611 ^ t58611;
    wire t58613 = t58612 ^ t58612;
    wire t58614 = t58613 ^ t58613;
    wire t58615 = t58614 ^ t58614;
    wire t58616 = t58615 ^ t58615;
    wire t58617 = t58616 ^ t58616;
    wire t58618 = t58617 ^ t58617;
    wire t58619 = t58618 ^ t58618;
    wire t58620 = t58619 ^ t58619;
    wire t58621 = t58620 ^ t58620;
    wire t58622 = t58621 ^ t58621;
    wire t58623 = t58622 ^ t58622;
    wire t58624 = t58623 ^ t58623;
    wire t58625 = t58624 ^ t58624;
    wire t58626 = t58625 ^ t58625;
    wire t58627 = t58626 ^ t58626;
    wire t58628 = t58627 ^ t58627;
    wire t58629 = t58628 ^ t58628;
    wire t58630 = t58629 ^ t58629;
    wire t58631 = t58630 ^ t58630;
    wire t58632 = t58631 ^ t58631;
    wire t58633 = t58632 ^ t58632;
    wire t58634 = t58633 ^ t58633;
    wire t58635 = t58634 ^ t58634;
    wire t58636 = t58635 ^ t58635;
    wire t58637 = t58636 ^ t58636;
    wire t58638 = t58637 ^ t58637;
    wire t58639 = t58638 ^ t58638;
    wire t58640 = t58639 ^ t58639;
    wire t58641 = t58640 ^ t58640;
    wire t58642 = t58641 ^ t58641;
    wire t58643 = t58642 ^ t58642;
    wire t58644 = t58643 ^ t58643;
    wire t58645 = t58644 ^ t58644;
    wire t58646 = t58645 ^ t58645;
    wire t58647 = t58646 ^ t58646;
    wire t58648 = t58647 ^ t58647;
    wire t58649 = t58648 ^ t58648;
    wire t58650 = t58649 ^ t58649;
    wire t58651 = t58650 ^ t58650;
    wire t58652 = t58651 ^ t58651;
    wire t58653 = t58652 ^ t58652;
    wire t58654 = t58653 ^ t58653;
    wire t58655 = t58654 ^ t58654;
    wire t58656 = t58655 ^ t58655;
    wire t58657 = t58656 ^ t58656;
    wire t58658 = t58657 ^ t58657;
    wire t58659 = t58658 ^ t58658;
    wire t58660 = t58659 ^ t58659;
    wire t58661 = t58660 ^ t58660;
    wire t58662 = t58661 ^ t58661;
    wire t58663 = t58662 ^ t58662;
    wire t58664 = t58663 ^ t58663;
    wire t58665 = t58664 ^ t58664;
    wire t58666 = t58665 ^ t58665;
    wire t58667 = t58666 ^ t58666;
    wire t58668 = t58667 ^ t58667;
    wire t58669 = t58668 ^ t58668;
    wire t58670 = t58669 ^ t58669;
    wire t58671 = t58670 ^ t58670;
    wire t58672 = t58671 ^ t58671;
    wire t58673 = t58672 ^ t58672;
    wire t58674 = t58673 ^ t58673;
    wire t58675 = t58674 ^ t58674;
    wire t58676 = t58675 ^ t58675;
    wire t58677 = t58676 ^ t58676;
    wire t58678 = t58677 ^ t58677;
    wire t58679 = t58678 ^ t58678;
    wire t58680 = t58679 ^ t58679;
    wire t58681 = t58680 ^ t58680;
    wire t58682 = t58681 ^ t58681;
    wire t58683 = t58682 ^ t58682;
    wire t58684 = t58683 ^ t58683;
    wire t58685 = t58684 ^ t58684;
    wire t58686 = t58685 ^ t58685;
    wire t58687 = t58686 ^ t58686;
    wire t58688 = t58687 ^ t58687;
    wire t58689 = t58688 ^ t58688;
    wire t58690 = t58689 ^ t58689;
    wire t58691 = t58690 ^ t58690;
    wire t58692 = t58691 ^ t58691;
    wire t58693 = t58692 ^ t58692;
    wire t58694 = t58693 ^ t58693;
    wire t58695 = t58694 ^ t58694;
    wire t58696 = t58695 ^ t58695;
    wire t58697 = t58696 ^ t58696;
    wire t58698 = t58697 ^ t58697;
    wire t58699 = t58698 ^ t58698;
    wire t58700 = t58699 ^ t58699;
    wire t58701 = t58700 ^ t58700;
    wire t58702 = t58701 ^ t58701;
    wire t58703 = t58702 ^ t58702;
    wire t58704 = t58703 ^ t58703;
    wire t58705 = t58704 ^ t58704;
    wire t58706 = t58705 ^ t58705;
    wire t58707 = t58706 ^ t58706;
    wire t58708 = t58707 ^ t58707;
    wire t58709 = t58708 ^ t58708;
    wire t58710 = t58709 ^ t58709;
    wire t58711 = t58710 ^ t58710;
    wire t58712 = t58711 ^ t58711;
    wire t58713 = t58712 ^ t58712;
    wire t58714 = t58713 ^ t58713;
    wire t58715 = t58714 ^ t58714;
    wire t58716 = t58715 ^ t58715;
    wire t58717 = t58716 ^ t58716;
    wire t58718 = t58717 ^ t58717;
    wire t58719 = t58718 ^ t58718;
    wire t58720 = t58719 ^ t58719;
    wire t58721 = t58720 ^ t58720;
    wire t58722 = t58721 ^ t58721;
    wire t58723 = t58722 ^ t58722;
    wire t58724 = t58723 ^ t58723;
    wire t58725 = t58724 ^ t58724;
    wire t58726 = t58725 ^ t58725;
    wire t58727 = t58726 ^ t58726;
    wire t58728 = t58727 ^ t58727;
    wire t58729 = t58728 ^ t58728;
    wire t58730 = t58729 ^ t58729;
    wire t58731 = t58730 ^ t58730;
    wire t58732 = t58731 ^ t58731;
    wire t58733 = t58732 ^ t58732;
    wire t58734 = t58733 ^ t58733;
    wire t58735 = t58734 ^ t58734;
    wire t58736 = t58735 ^ t58735;
    wire t58737 = t58736 ^ t58736;
    wire t58738 = t58737 ^ t58737;
    wire t58739 = t58738 ^ t58738;
    wire t58740 = t58739 ^ t58739;
    wire t58741 = t58740 ^ t58740;
    wire t58742 = t58741 ^ t58741;
    wire t58743 = t58742 ^ t58742;
    wire t58744 = t58743 ^ t58743;
    wire t58745 = t58744 ^ t58744;
    wire t58746 = t58745 ^ t58745;
    wire t58747 = t58746 ^ t58746;
    wire t58748 = t58747 ^ t58747;
    wire t58749 = t58748 ^ t58748;
    wire t58750 = t58749 ^ t58749;
    wire t58751 = t58750 ^ t58750;
    wire t58752 = t58751 ^ t58751;
    wire t58753 = t58752 ^ t58752;
    wire t58754 = t58753 ^ t58753;
    wire t58755 = t58754 ^ t58754;
    wire t58756 = t58755 ^ t58755;
    wire t58757 = t58756 ^ t58756;
    wire t58758 = t58757 ^ t58757;
    wire t58759 = t58758 ^ t58758;
    wire t58760 = t58759 ^ t58759;
    wire t58761 = t58760 ^ t58760;
    wire t58762 = t58761 ^ t58761;
    wire t58763 = t58762 ^ t58762;
    wire t58764 = t58763 ^ t58763;
    wire t58765 = t58764 ^ t58764;
    wire t58766 = t58765 ^ t58765;
    wire t58767 = t58766 ^ t58766;
    wire t58768 = t58767 ^ t58767;
    wire t58769 = t58768 ^ t58768;
    wire t58770 = t58769 ^ t58769;
    wire t58771 = t58770 ^ t58770;
    wire t58772 = t58771 ^ t58771;
    wire t58773 = t58772 ^ t58772;
    wire t58774 = t58773 ^ t58773;
    wire t58775 = t58774 ^ t58774;
    wire t58776 = t58775 ^ t58775;
    wire t58777 = t58776 ^ t58776;
    wire t58778 = t58777 ^ t58777;
    wire t58779 = t58778 ^ t58778;
    wire t58780 = t58779 ^ t58779;
    wire t58781 = t58780 ^ t58780;
    wire t58782 = t58781 ^ t58781;
    wire t58783 = t58782 ^ t58782;
    wire t58784 = t58783 ^ t58783;
    wire t58785 = t58784 ^ t58784;
    wire t58786 = t58785 ^ t58785;
    wire t58787 = t58786 ^ t58786;
    wire t58788 = t58787 ^ t58787;
    wire t58789 = t58788 ^ t58788;
    wire t58790 = t58789 ^ t58789;
    wire t58791 = t58790 ^ t58790;
    wire t58792 = t58791 ^ t58791;
    wire t58793 = t58792 ^ t58792;
    wire t58794 = t58793 ^ t58793;
    wire t58795 = t58794 ^ t58794;
    wire t58796 = t58795 ^ t58795;
    wire t58797 = t58796 ^ t58796;
    wire t58798 = t58797 ^ t58797;
    wire t58799 = t58798 ^ t58798;
    wire t58800 = t58799 ^ t58799;
    wire t58801 = t58800 ^ t58800;
    wire t58802 = t58801 ^ t58801;
    wire t58803 = t58802 ^ t58802;
    wire t58804 = t58803 ^ t58803;
    wire t58805 = t58804 ^ t58804;
    wire t58806 = t58805 ^ t58805;
    wire t58807 = t58806 ^ t58806;
    wire t58808 = t58807 ^ t58807;
    wire t58809 = t58808 ^ t58808;
    wire t58810 = t58809 ^ t58809;
    wire t58811 = t58810 ^ t58810;
    wire t58812 = t58811 ^ t58811;
    wire t58813 = t58812 ^ t58812;
    wire t58814 = t58813 ^ t58813;
    wire t58815 = t58814 ^ t58814;
    wire t58816 = t58815 ^ t58815;
    wire t58817 = t58816 ^ t58816;
    wire t58818 = t58817 ^ t58817;
    wire t58819 = t58818 ^ t58818;
    wire t58820 = t58819 ^ t58819;
    wire t58821 = t58820 ^ t58820;
    wire t58822 = t58821 ^ t58821;
    wire t58823 = t58822 ^ t58822;
    wire t58824 = t58823 ^ t58823;
    wire t58825 = t58824 ^ t58824;
    wire t58826 = t58825 ^ t58825;
    wire t58827 = t58826 ^ t58826;
    wire t58828 = t58827 ^ t58827;
    wire t58829 = t58828 ^ t58828;
    wire t58830 = t58829 ^ t58829;
    wire t58831 = t58830 ^ t58830;
    wire t58832 = t58831 ^ t58831;
    wire t58833 = t58832 ^ t58832;
    wire t58834 = t58833 ^ t58833;
    wire t58835 = t58834 ^ t58834;
    wire t58836 = t58835 ^ t58835;
    wire t58837 = t58836 ^ t58836;
    wire t58838 = t58837 ^ t58837;
    wire t58839 = t58838 ^ t58838;
    wire t58840 = t58839 ^ t58839;
    wire t58841 = t58840 ^ t58840;
    wire t58842 = t58841 ^ t58841;
    wire t58843 = t58842 ^ t58842;
    wire t58844 = t58843 ^ t58843;
    wire t58845 = t58844 ^ t58844;
    wire t58846 = t58845 ^ t58845;
    wire t58847 = t58846 ^ t58846;
    wire t58848 = t58847 ^ t58847;
    wire t58849 = t58848 ^ t58848;
    wire t58850 = t58849 ^ t58849;
    wire t58851 = t58850 ^ t58850;
    wire t58852 = t58851 ^ t58851;
    wire t58853 = t58852 ^ t58852;
    wire t58854 = t58853 ^ t58853;
    wire t58855 = t58854 ^ t58854;
    wire t58856 = t58855 ^ t58855;
    wire t58857 = t58856 ^ t58856;
    wire t58858 = t58857 ^ t58857;
    wire t58859 = t58858 ^ t58858;
    wire t58860 = t58859 ^ t58859;
    wire t58861 = t58860 ^ t58860;
    wire t58862 = t58861 ^ t58861;
    wire t58863 = t58862 ^ t58862;
    wire t58864 = t58863 ^ t58863;
    wire t58865 = t58864 ^ t58864;
    wire t58866 = t58865 ^ t58865;
    wire t58867 = t58866 ^ t58866;
    wire t58868 = t58867 ^ t58867;
    wire t58869 = t58868 ^ t58868;
    wire t58870 = t58869 ^ t58869;
    wire t58871 = t58870 ^ t58870;
    wire t58872 = t58871 ^ t58871;
    wire t58873 = t58872 ^ t58872;
    wire t58874 = t58873 ^ t58873;
    wire t58875 = t58874 ^ t58874;
    wire t58876 = t58875 ^ t58875;
    wire t58877 = t58876 ^ t58876;
    wire t58878 = t58877 ^ t58877;
    wire t58879 = t58878 ^ t58878;
    wire t58880 = t58879 ^ t58879;
    wire t58881 = t58880 ^ t58880;
    wire t58882 = t58881 ^ t58881;
    wire t58883 = t58882 ^ t58882;
    wire t58884 = t58883 ^ t58883;
    wire t58885 = t58884 ^ t58884;
    wire t58886 = t58885 ^ t58885;
    wire t58887 = t58886 ^ t58886;
    wire t58888 = t58887 ^ t58887;
    wire t58889 = t58888 ^ t58888;
    wire t58890 = t58889 ^ t58889;
    wire t58891 = t58890 ^ t58890;
    wire t58892 = t58891 ^ t58891;
    wire t58893 = t58892 ^ t58892;
    wire t58894 = t58893 ^ t58893;
    wire t58895 = t58894 ^ t58894;
    wire t58896 = t58895 ^ t58895;
    wire t58897 = t58896 ^ t58896;
    wire t58898 = t58897 ^ t58897;
    wire t58899 = t58898 ^ t58898;
    wire t58900 = t58899 ^ t58899;
    wire t58901 = t58900 ^ t58900;
    wire t58902 = t58901 ^ t58901;
    wire t58903 = t58902 ^ t58902;
    wire t58904 = t58903 ^ t58903;
    wire t58905 = t58904 ^ t58904;
    wire t58906 = t58905 ^ t58905;
    wire t58907 = t58906 ^ t58906;
    wire t58908 = t58907 ^ t58907;
    wire t58909 = t58908 ^ t58908;
    wire t58910 = t58909 ^ t58909;
    wire t58911 = t58910 ^ t58910;
    wire t58912 = t58911 ^ t58911;
    wire t58913 = t58912 ^ t58912;
    wire t58914 = t58913 ^ t58913;
    wire t58915 = t58914 ^ t58914;
    wire t58916 = t58915 ^ t58915;
    wire t58917 = t58916 ^ t58916;
    wire t58918 = t58917 ^ t58917;
    wire t58919 = t58918 ^ t58918;
    wire t58920 = t58919 ^ t58919;
    wire t58921 = t58920 ^ t58920;
    wire t58922 = t58921 ^ t58921;
    wire t58923 = t58922 ^ t58922;
    wire t58924 = t58923 ^ t58923;
    wire t58925 = t58924 ^ t58924;
    wire t58926 = t58925 ^ t58925;
    wire t58927 = t58926 ^ t58926;
    wire t58928 = t58927 ^ t58927;
    wire t58929 = t58928 ^ t58928;
    wire t58930 = t58929 ^ t58929;
    wire t58931 = t58930 ^ t58930;
    wire t58932 = t58931 ^ t58931;
    wire t58933 = t58932 ^ t58932;
    wire t58934 = t58933 ^ t58933;
    wire t58935 = t58934 ^ t58934;
    wire t58936 = t58935 ^ t58935;
    wire t58937 = t58936 ^ t58936;
    wire t58938 = t58937 ^ t58937;
    wire t58939 = t58938 ^ t58938;
    wire t58940 = t58939 ^ t58939;
    wire t58941 = t58940 ^ t58940;
    wire t58942 = t58941 ^ t58941;
    wire t58943 = t58942 ^ t58942;
    wire t58944 = t58943 ^ t58943;
    wire t58945 = t58944 ^ t58944;
    wire t58946 = t58945 ^ t58945;
    wire t58947 = t58946 ^ t58946;
    wire t58948 = t58947 ^ t58947;
    wire t58949 = t58948 ^ t58948;
    wire t58950 = t58949 ^ t58949;
    wire t58951 = t58950 ^ t58950;
    wire t58952 = t58951 ^ t58951;
    wire t58953 = t58952 ^ t58952;
    wire t58954 = t58953 ^ t58953;
    wire t58955 = t58954 ^ t58954;
    wire t58956 = t58955 ^ t58955;
    wire t58957 = t58956 ^ t58956;
    wire t58958 = t58957 ^ t58957;
    wire t58959 = t58958 ^ t58958;
    wire t58960 = t58959 ^ t58959;
    wire t58961 = t58960 ^ t58960;
    wire t58962 = t58961 ^ t58961;
    wire t58963 = t58962 ^ t58962;
    wire t58964 = t58963 ^ t58963;
    wire t58965 = t58964 ^ t58964;
    wire t58966 = t58965 ^ t58965;
    wire t58967 = t58966 ^ t58966;
    wire t58968 = t58967 ^ t58967;
    wire t58969 = t58968 ^ t58968;
    wire t58970 = t58969 ^ t58969;
    wire t58971 = t58970 ^ t58970;
    wire t58972 = t58971 ^ t58971;
    wire t58973 = t58972 ^ t58972;
    wire t58974 = t58973 ^ t58973;
    wire t58975 = t58974 ^ t58974;
    wire t58976 = t58975 ^ t58975;
    wire t58977 = t58976 ^ t58976;
    wire t58978 = t58977 ^ t58977;
    wire t58979 = t58978 ^ t58978;
    wire t58980 = t58979 ^ t58979;
    wire t58981 = t58980 ^ t58980;
    wire t58982 = t58981 ^ t58981;
    wire t58983 = t58982 ^ t58982;
    wire t58984 = t58983 ^ t58983;
    wire t58985 = t58984 ^ t58984;
    wire t58986 = t58985 ^ t58985;
    wire t58987 = t58986 ^ t58986;
    wire t58988 = t58987 ^ t58987;
    wire t58989 = t58988 ^ t58988;
    wire t58990 = t58989 ^ t58989;
    wire t58991 = t58990 ^ t58990;
    wire t58992 = t58991 ^ t58991;
    wire t58993 = t58992 ^ t58992;
    wire t58994 = t58993 ^ t58993;
    wire t58995 = t58994 ^ t58994;
    wire t58996 = t58995 ^ t58995;
    wire t58997 = t58996 ^ t58996;
    wire t58998 = t58997 ^ t58997;
    wire t58999 = t58998 ^ t58998;
    wire t59000 = t58999 ^ t58999;
    wire t59001 = t59000 ^ t59000;
    wire t59002 = t59001 ^ t59001;
    wire t59003 = t59002 ^ t59002;
    wire t59004 = t59003 ^ t59003;
    wire t59005 = t59004 ^ t59004;
    wire t59006 = t59005 ^ t59005;
    wire t59007 = t59006 ^ t59006;
    wire t59008 = t59007 ^ t59007;
    wire t59009 = t59008 ^ t59008;
    wire t59010 = t59009 ^ t59009;
    wire t59011 = t59010 ^ t59010;
    wire t59012 = t59011 ^ t59011;
    wire t59013 = t59012 ^ t59012;
    wire t59014 = t59013 ^ t59013;
    wire t59015 = t59014 ^ t59014;
    wire t59016 = t59015 ^ t59015;
    wire t59017 = t59016 ^ t59016;
    wire t59018 = t59017 ^ t59017;
    wire t59019 = t59018 ^ t59018;
    wire t59020 = t59019 ^ t59019;
    wire t59021 = t59020 ^ t59020;
    wire t59022 = t59021 ^ t59021;
    wire t59023 = t59022 ^ t59022;
    wire t59024 = t59023 ^ t59023;
    wire t59025 = t59024 ^ t59024;
    wire t59026 = t59025 ^ t59025;
    wire t59027 = t59026 ^ t59026;
    wire t59028 = t59027 ^ t59027;
    wire t59029 = t59028 ^ t59028;
    wire t59030 = t59029 ^ t59029;
    wire t59031 = t59030 ^ t59030;
    wire t59032 = t59031 ^ t59031;
    wire t59033 = t59032 ^ t59032;
    wire t59034 = t59033 ^ t59033;
    wire t59035 = t59034 ^ t59034;
    wire t59036 = t59035 ^ t59035;
    wire t59037 = t59036 ^ t59036;
    wire t59038 = t59037 ^ t59037;
    wire t59039 = t59038 ^ t59038;
    wire t59040 = t59039 ^ t59039;
    wire t59041 = t59040 ^ t59040;
    wire t59042 = t59041 ^ t59041;
    wire t59043 = t59042 ^ t59042;
    wire t59044 = t59043 ^ t59043;
    wire t59045 = t59044 ^ t59044;
    wire t59046 = t59045 ^ t59045;
    wire t59047 = t59046 ^ t59046;
    wire t59048 = t59047 ^ t59047;
    wire t59049 = t59048 ^ t59048;
    wire t59050 = t59049 ^ t59049;
    wire t59051 = t59050 ^ t59050;
    wire t59052 = t59051 ^ t59051;
    wire t59053 = t59052 ^ t59052;
    wire t59054 = t59053 ^ t59053;
    wire t59055 = t59054 ^ t59054;
    wire t59056 = t59055 ^ t59055;
    wire t59057 = t59056 ^ t59056;
    wire t59058 = t59057 ^ t59057;
    wire t59059 = t59058 ^ t59058;
    wire t59060 = t59059 ^ t59059;
    wire t59061 = t59060 ^ t59060;
    wire t59062 = t59061 ^ t59061;
    wire t59063 = t59062 ^ t59062;
    wire t59064 = t59063 ^ t59063;
    wire t59065 = t59064 ^ t59064;
    wire t59066 = t59065 ^ t59065;
    wire t59067 = t59066 ^ t59066;
    wire t59068 = t59067 ^ t59067;
    wire t59069 = t59068 ^ t59068;
    wire t59070 = t59069 ^ t59069;
    wire t59071 = t59070 ^ t59070;
    wire t59072 = t59071 ^ t59071;
    wire t59073 = t59072 ^ t59072;
    wire t59074 = t59073 ^ t59073;
    wire t59075 = t59074 ^ t59074;
    wire t59076 = t59075 ^ t59075;
    wire t59077 = t59076 ^ t59076;
    wire t59078 = t59077 ^ t59077;
    wire t59079 = t59078 ^ t59078;
    wire t59080 = t59079 ^ t59079;
    wire t59081 = t59080 ^ t59080;
    wire t59082 = t59081 ^ t59081;
    wire t59083 = t59082 ^ t59082;
    wire t59084 = t59083 ^ t59083;
    wire t59085 = t59084 ^ t59084;
    wire t59086 = t59085 ^ t59085;
    wire t59087 = t59086 ^ t59086;
    wire t59088 = t59087 ^ t59087;
    wire t59089 = t59088 ^ t59088;
    wire t59090 = t59089 ^ t59089;
    wire t59091 = t59090 ^ t59090;
    wire t59092 = t59091 ^ t59091;
    wire t59093 = t59092 ^ t59092;
    wire t59094 = t59093 ^ t59093;
    wire t59095 = t59094 ^ t59094;
    wire t59096 = t59095 ^ t59095;
    wire t59097 = t59096 ^ t59096;
    wire t59098 = t59097 ^ t59097;
    wire t59099 = t59098 ^ t59098;
    wire t59100 = t59099 ^ t59099;
    wire t59101 = t59100 ^ t59100;
    wire t59102 = t59101 ^ t59101;
    wire t59103 = t59102 ^ t59102;
    wire t59104 = t59103 ^ t59103;
    wire t59105 = t59104 ^ t59104;
    wire t59106 = t59105 ^ t59105;
    wire t59107 = t59106 ^ t59106;
    wire t59108 = t59107 ^ t59107;
    wire t59109 = t59108 ^ t59108;
    wire t59110 = t59109 ^ t59109;
    wire t59111 = t59110 ^ t59110;
    wire t59112 = t59111 ^ t59111;
    wire t59113 = t59112 ^ t59112;
    wire t59114 = t59113 ^ t59113;
    wire t59115 = t59114 ^ t59114;
    wire t59116 = t59115 ^ t59115;
    wire t59117 = t59116 ^ t59116;
    wire t59118 = t59117 ^ t59117;
    wire t59119 = t59118 ^ t59118;
    wire t59120 = t59119 ^ t59119;
    wire t59121 = t59120 ^ t59120;
    wire t59122 = t59121 ^ t59121;
    wire t59123 = t59122 ^ t59122;
    wire t59124 = t59123 ^ t59123;
    wire t59125 = t59124 ^ t59124;
    wire t59126 = t59125 ^ t59125;
    wire t59127 = t59126 ^ t59126;
    wire t59128 = t59127 ^ t59127;
    wire t59129 = t59128 ^ t59128;
    wire t59130 = t59129 ^ t59129;
    wire t59131 = t59130 ^ t59130;
    wire t59132 = t59131 ^ t59131;
    wire t59133 = t59132 ^ t59132;
    wire t59134 = t59133 ^ t59133;
    wire t59135 = t59134 ^ t59134;
    wire t59136 = t59135 ^ t59135;
    wire t59137 = t59136 ^ t59136;
    wire t59138 = t59137 ^ t59137;
    wire t59139 = t59138 ^ t59138;
    wire t59140 = t59139 ^ t59139;
    wire t59141 = t59140 ^ t59140;
    wire t59142 = t59141 ^ t59141;
    wire t59143 = t59142 ^ t59142;
    wire t59144 = t59143 ^ t59143;
    wire t59145 = t59144 ^ t59144;
    wire t59146 = t59145 ^ t59145;
    wire t59147 = t59146 ^ t59146;
    wire t59148 = t59147 ^ t59147;
    wire t59149 = t59148 ^ t59148;
    wire t59150 = t59149 ^ t59149;
    wire t59151 = t59150 ^ t59150;
    wire t59152 = t59151 ^ t59151;
    wire t59153 = t59152 ^ t59152;
    wire t59154 = t59153 ^ t59153;
    wire t59155 = t59154 ^ t59154;
    wire t59156 = t59155 ^ t59155;
    wire t59157 = t59156 ^ t59156;
    wire t59158 = t59157 ^ t59157;
    wire t59159 = t59158 ^ t59158;
    wire t59160 = t59159 ^ t59159;
    wire t59161 = t59160 ^ t59160;
    wire t59162 = t59161 ^ t59161;
    wire t59163 = t59162 ^ t59162;
    wire t59164 = t59163 ^ t59163;
    wire t59165 = t59164 ^ t59164;
    wire t59166 = t59165 ^ t59165;
    wire t59167 = t59166 ^ t59166;
    wire t59168 = t59167 ^ t59167;
    wire t59169 = t59168 ^ t59168;
    wire t59170 = t59169 ^ t59169;
    wire t59171 = t59170 ^ t59170;
    wire t59172 = t59171 ^ t59171;
    wire t59173 = t59172 ^ t59172;
    wire t59174 = t59173 ^ t59173;
    wire t59175 = t59174 ^ t59174;
    wire t59176 = t59175 ^ t59175;
    wire t59177 = t59176 ^ t59176;
    wire t59178 = t59177 ^ t59177;
    wire t59179 = t59178 ^ t59178;
    wire t59180 = t59179 ^ t59179;
    wire t59181 = t59180 ^ t59180;
    wire t59182 = t59181 ^ t59181;
    wire t59183 = t59182 ^ t59182;
    wire t59184 = t59183 ^ t59183;
    wire t59185 = t59184 ^ t59184;
    wire t59186 = t59185 ^ t59185;
    wire t59187 = t59186 ^ t59186;
    wire t59188 = t59187 ^ t59187;
    wire t59189 = t59188 ^ t59188;
    wire t59190 = t59189 ^ t59189;
    wire t59191 = t59190 ^ t59190;
    wire t59192 = t59191 ^ t59191;
    wire t59193 = t59192 ^ t59192;
    wire t59194 = t59193 ^ t59193;
    wire t59195 = t59194 ^ t59194;
    wire t59196 = t59195 ^ t59195;
    wire t59197 = t59196 ^ t59196;
    wire t59198 = t59197 ^ t59197;
    wire t59199 = t59198 ^ t59198;
    wire t59200 = t59199 ^ t59199;
    wire t59201 = t59200 ^ t59200;
    wire t59202 = t59201 ^ t59201;
    wire t59203 = t59202 ^ t59202;
    wire t59204 = t59203 ^ t59203;
    wire t59205 = t59204 ^ t59204;
    wire t59206 = t59205 ^ t59205;
    wire t59207 = t59206 ^ t59206;
    wire t59208 = t59207 ^ t59207;
    wire t59209 = t59208 ^ t59208;
    wire t59210 = t59209 ^ t59209;
    wire t59211 = t59210 ^ t59210;
    wire t59212 = t59211 ^ t59211;
    wire t59213 = t59212 ^ t59212;
    wire t59214 = t59213 ^ t59213;
    wire t59215 = t59214 ^ t59214;
    wire t59216 = t59215 ^ t59215;
    wire t59217 = t59216 ^ t59216;
    wire t59218 = t59217 ^ t59217;
    wire t59219 = t59218 ^ t59218;
    wire t59220 = t59219 ^ t59219;
    wire t59221 = t59220 ^ t59220;
    wire t59222 = t59221 ^ t59221;
    wire t59223 = t59222 ^ t59222;
    wire t59224 = t59223 ^ t59223;
    wire t59225 = t59224 ^ t59224;
    wire t59226 = t59225 ^ t59225;
    wire t59227 = t59226 ^ t59226;
    wire t59228 = t59227 ^ t59227;
    wire t59229 = t59228 ^ t59228;
    wire t59230 = t59229 ^ t59229;
    wire t59231 = t59230 ^ t59230;
    wire t59232 = t59231 ^ t59231;
    wire t59233 = t59232 ^ t59232;
    wire t59234 = t59233 ^ t59233;
    wire t59235 = t59234 ^ t59234;
    wire t59236 = t59235 ^ t59235;
    wire t59237 = t59236 ^ t59236;
    wire t59238 = t59237 ^ t59237;
    wire t59239 = t59238 ^ t59238;
    wire t59240 = t59239 ^ t59239;
    wire t59241 = t59240 ^ t59240;
    wire t59242 = t59241 ^ t59241;
    wire t59243 = t59242 ^ t59242;
    wire t59244 = t59243 ^ t59243;
    wire t59245 = t59244 ^ t59244;
    wire t59246 = t59245 ^ t59245;
    wire t59247 = t59246 ^ t59246;
    wire t59248 = t59247 ^ t59247;
    wire t59249 = t59248 ^ t59248;
    wire t59250 = t59249 ^ t59249;
    wire t59251 = t59250 ^ t59250;
    wire t59252 = t59251 ^ t59251;
    wire t59253 = t59252 ^ t59252;
    wire t59254 = t59253 ^ t59253;
    wire t59255 = t59254 ^ t59254;
    wire t59256 = t59255 ^ t59255;
    wire t59257 = t59256 ^ t59256;
    wire t59258 = t59257 ^ t59257;
    wire t59259 = t59258 ^ t59258;
    wire t59260 = t59259 ^ t59259;
    wire t59261 = t59260 ^ t59260;
    wire t59262 = t59261 ^ t59261;
    wire t59263 = t59262 ^ t59262;
    wire t59264 = t59263 ^ t59263;
    wire t59265 = t59264 ^ t59264;
    wire t59266 = t59265 ^ t59265;
    wire t59267 = t59266 ^ t59266;
    wire t59268 = t59267 ^ t59267;
    wire t59269 = t59268 ^ t59268;
    wire t59270 = t59269 ^ t59269;
    wire t59271 = t59270 ^ t59270;
    wire t59272 = t59271 ^ t59271;
    wire t59273 = t59272 ^ t59272;
    wire t59274 = t59273 ^ t59273;
    wire t59275 = t59274 ^ t59274;
    wire t59276 = t59275 ^ t59275;
    wire t59277 = t59276 ^ t59276;
    wire t59278 = t59277 ^ t59277;
    wire t59279 = t59278 ^ t59278;
    wire t59280 = t59279 ^ t59279;
    wire t59281 = t59280 ^ t59280;
    wire t59282 = t59281 ^ t59281;
    wire t59283 = t59282 ^ t59282;
    wire t59284 = t59283 ^ t59283;
    wire t59285 = t59284 ^ t59284;
    wire t59286 = t59285 ^ t59285;
    wire t59287 = t59286 ^ t59286;
    wire t59288 = t59287 ^ t59287;
    wire t59289 = t59288 ^ t59288;
    wire t59290 = t59289 ^ t59289;
    wire t59291 = t59290 ^ t59290;
    wire t59292 = t59291 ^ t59291;
    wire t59293 = t59292 ^ t59292;
    wire t59294 = t59293 ^ t59293;
    wire t59295 = t59294 ^ t59294;
    wire t59296 = t59295 ^ t59295;
    wire t59297 = t59296 ^ t59296;
    wire t59298 = t59297 ^ t59297;
    wire t59299 = t59298 ^ t59298;
    wire t59300 = t59299 ^ t59299;
    wire t59301 = t59300 ^ t59300;
    wire t59302 = t59301 ^ t59301;
    wire t59303 = t59302 ^ t59302;
    wire t59304 = t59303 ^ t59303;
    wire t59305 = t59304 ^ t59304;
    wire t59306 = t59305 ^ t59305;
    wire t59307 = t59306 ^ t59306;
    wire t59308 = t59307 ^ t59307;
    wire t59309 = t59308 ^ t59308;
    wire t59310 = t59309 ^ t59309;
    wire t59311 = t59310 ^ t59310;
    wire t59312 = t59311 ^ t59311;
    wire t59313 = t59312 ^ t59312;
    wire t59314 = t59313 ^ t59313;
    wire t59315 = t59314 ^ t59314;
    wire t59316 = t59315 ^ t59315;
    wire t59317 = t59316 ^ t59316;
    wire t59318 = t59317 ^ t59317;
    wire t59319 = t59318 ^ t59318;
    wire t59320 = t59319 ^ t59319;
    wire t59321 = t59320 ^ t59320;
    wire t59322 = t59321 ^ t59321;
    wire t59323 = t59322 ^ t59322;
    wire t59324 = t59323 ^ t59323;
    wire t59325 = t59324 ^ t59324;
    wire t59326 = t59325 ^ t59325;
    wire t59327 = t59326 ^ t59326;
    wire t59328 = t59327 ^ t59327;
    wire t59329 = t59328 ^ t59328;
    wire t59330 = t59329 ^ t59329;
    wire t59331 = t59330 ^ t59330;
    wire t59332 = t59331 ^ t59331;
    wire t59333 = t59332 ^ t59332;
    wire t59334 = t59333 ^ t59333;
    wire t59335 = t59334 ^ t59334;
    wire t59336 = t59335 ^ t59335;
    wire t59337 = t59336 ^ t59336;
    wire t59338 = t59337 ^ t59337;
    wire t59339 = t59338 ^ t59338;
    wire t59340 = t59339 ^ t59339;
    wire t59341 = t59340 ^ t59340;
    wire t59342 = t59341 ^ t59341;
    wire t59343 = t59342 ^ t59342;
    wire t59344 = t59343 ^ t59343;
    wire t59345 = t59344 ^ t59344;
    wire t59346 = t59345 ^ t59345;
    wire t59347 = t59346 ^ t59346;
    wire t59348 = t59347 ^ t59347;
    wire t59349 = t59348 ^ t59348;
    wire t59350 = t59349 ^ t59349;
    wire t59351 = t59350 ^ t59350;
    wire t59352 = t59351 ^ t59351;
    wire t59353 = t59352 ^ t59352;
    wire t59354 = t59353 ^ t59353;
    wire t59355 = t59354 ^ t59354;
    wire t59356 = t59355 ^ t59355;
    wire t59357 = t59356 ^ t59356;
    wire t59358 = t59357 ^ t59357;
    wire t59359 = t59358 ^ t59358;
    wire t59360 = t59359 ^ t59359;
    wire t59361 = t59360 ^ t59360;
    wire t59362 = t59361 ^ t59361;
    wire t59363 = t59362 ^ t59362;
    wire t59364 = t59363 ^ t59363;
    wire t59365 = t59364 ^ t59364;
    wire t59366 = t59365 ^ t59365;
    wire t59367 = t59366 ^ t59366;
    wire t59368 = t59367 ^ t59367;
    wire t59369 = t59368 ^ t59368;
    wire t59370 = t59369 ^ t59369;
    wire t59371 = t59370 ^ t59370;
    wire t59372 = t59371 ^ t59371;
    wire t59373 = t59372 ^ t59372;
    wire t59374 = t59373 ^ t59373;
    wire t59375 = t59374 ^ t59374;
    wire t59376 = t59375 ^ t59375;
    wire t59377 = t59376 ^ t59376;
    wire t59378 = t59377 ^ t59377;
    wire t59379 = t59378 ^ t59378;
    wire t59380 = t59379 ^ t59379;
    wire t59381 = t59380 ^ t59380;
    wire t59382 = t59381 ^ t59381;
    wire t59383 = t59382 ^ t59382;
    wire t59384 = t59383 ^ t59383;
    wire t59385 = t59384 ^ t59384;
    wire t59386 = t59385 ^ t59385;
    wire t59387 = t59386 ^ t59386;
    wire t59388 = t59387 ^ t59387;
    wire t59389 = t59388 ^ t59388;
    wire t59390 = t59389 ^ t59389;
    wire t59391 = t59390 ^ t59390;
    wire t59392 = t59391 ^ t59391;
    wire t59393 = t59392 ^ t59392;
    wire t59394 = t59393 ^ t59393;
    wire t59395 = t59394 ^ t59394;
    wire t59396 = t59395 ^ t59395;
    wire t59397 = t59396 ^ t59396;
    wire t59398 = t59397 ^ t59397;
    wire t59399 = t59398 ^ t59398;
    wire t59400 = t59399 ^ t59399;
    wire t59401 = t59400 ^ t59400;
    wire t59402 = t59401 ^ t59401;
    wire t59403 = t59402 ^ t59402;
    wire t59404 = t59403 ^ t59403;
    wire t59405 = t59404 ^ t59404;
    wire t59406 = t59405 ^ t59405;
    wire t59407 = t59406 ^ t59406;
    wire t59408 = t59407 ^ t59407;
    wire t59409 = t59408 ^ t59408;
    wire t59410 = t59409 ^ t59409;
    wire t59411 = t59410 ^ t59410;
    wire t59412 = t59411 ^ t59411;
    wire t59413 = t59412 ^ t59412;
    wire t59414 = t59413 ^ t59413;
    wire t59415 = t59414 ^ t59414;
    wire t59416 = t59415 ^ t59415;
    wire t59417 = t59416 ^ t59416;
    wire t59418 = t59417 ^ t59417;
    wire t59419 = t59418 ^ t59418;
    wire t59420 = t59419 ^ t59419;
    wire t59421 = t59420 ^ t59420;
    wire t59422 = t59421 ^ t59421;
    wire t59423 = t59422 ^ t59422;
    wire t59424 = t59423 ^ t59423;
    wire t59425 = t59424 ^ t59424;
    wire t59426 = t59425 ^ t59425;
    wire t59427 = t59426 ^ t59426;
    wire t59428 = t59427 ^ t59427;
    wire t59429 = t59428 ^ t59428;
    wire t59430 = t59429 ^ t59429;
    wire t59431 = t59430 ^ t59430;
    wire t59432 = t59431 ^ t59431;
    wire t59433 = t59432 ^ t59432;
    wire t59434 = t59433 ^ t59433;
    wire t59435 = t59434 ^ t59434;
    wire t59436 = t59435 ^ t59435;
    wire t59437 = t59436 ^ t59436;
    wire t59438 = t59437 ^ t59437;
    wire t59439 = t59438 ^ t59438;
    wire t59440 = t59439 ^ t59439;
    wire t59441 = t59440 ^ t59440;
    wire t59442 = t59441 ^ t59441;
    wire t59443 = t59442 ^ t59442;
    wire t59444 = t59443 ^ t59443;
    wire t59445 = t59444 ^ t59444;
    wire t59446 = t59445 ^ t59445;
    wire t59447 = t59446 ^ t59446;
    wire t59448 = t59447 ^ t59447;
    wire t59449 = t59448 ^ t59448;
    wire t59450 = t59449 ^ t59449;
    wire t59451 = t59450 ^ t59450;
    wire t59452 = t59451 ^ t59451;
    wire t59453 = t59452 ^ t59452;
    wire t59454 = t59453 ^ t59453;
    wire t59455 = t59454 ^ t59454;
    wire t59456 = t59455 ^ t59455;
    wire t59457 = t59456 ^ t59456;
    wire t59458 = t59457 ^ t59457;
    wire t59459 = t59458 ^ t59458;
    wire t59460 = t59459 ^ t59459;
    wire t59461 = t59460 ^ t59460;
    wire t59462 = t59461 ^ t59461;
    wire t59463 = t59462 ^ t59462;
    wire t59464 = t59463 ^ t59463;
    wire t59465 = t59464 ^ t59464;
    wire t59466 = t59465 ^ t59465;
    wire t59467 = t59466 ^ t59466;
    wire t59468 = t59467 ^ t59467;
    wire t59469 = t59468 ^ t59468;
    wire t59470 = t59469 ^ t59469;
    wire t59471 = t59470 ^ t59470;
    wire t59472 = t59471 ^ t59471;
    wire t59473 = t59472 ^ t59472;
    wire t59474 = t59473 ^ t59473;
    wire t59475 = t59474 ^ t59474;
    wire t59476 = t59475 ^ t59475;
    wire t59477 = t59476 ^ t59476;
    wire t59478 = t59477 ^ t59477;
    wire t59479 = t59478 ^ t59478;
    wire t59480 = t59479 ^ t59479;
    wire t59481 = t59480 ^ t59480;
    wire t59482 = t59481 ^ t59481;
    wire t59483 = t59482 ^ t59482;
    wire t59484 = t59483 ^ t59483;
    wire t59485 = t59484 ^ t59484;
    wire t59486 = t59485 ^ t59485;
    wire t59487 = t59486 ^ t59486;
    wire t59488 = t59487 ^ t59487;
    wire t59489 = t59488 ^ t59488;
    wire t59490 = t59489 ^ t59489;
    wire t59491 = t59490 ^ t59490;
    wire t59492 = t59491 ^ t59491;
    wire t59493 = t59492 ^ t59492;
    wire t59494 = t59493 ^ t59493;
    wire t59495 = t59494 ^ t59494;
    wire t59496 = t59495 ^ t59495;
    wire t59497 = t59496 ^ t59496;
    wire t59498 = t59497 ^ t59497;
    wire t59499 = t59498 ^ t59498;
    wire t59500 = t59499 ^ t59499;
    wire t59501 = t59500 ^ t59500;
    wire t59502 = t59501 ^ t59501;
    wire t59503 = t59502 ^ t59502;
    wire t59504 = t59503 ^ t59503;
    wire t59505 = t59504 ^ t59504;
    wire t59506 = t59505 ^ t59505;
    wire t59507 = t59506 ^ t59506;
    wire t59508 = t59507 ^ t59507;
    wire t59509 = t59508 ^ t59508;
    wire t59510 = t59509 ^ t59509;
    wire t59511 = t59510 ^ t59510;
    wire t59512 = t59511 ^ t59511;
    wire t59513 = t59512 ^ t59512;
    wire t59514 = t59513 ^ t59513;
    wire t59515 = t59514 ^ t59514;
    wire t59516 = t59515 ^ t59515;
    wire t59517 = t59516 ^ t59516;
    wire t59518 = t59517 ^ t59517;
    wire t59519 = t59518 ^ t59518;
    wire t59520 = t59519 ^ t59519;
    wire t59521 = t59520 ^ t59520;
    wire t59522 = t59521 ^ t59521;
    wire t59523 = t59522 ^ t59522;
    wire t59524 = t59523 ^ t59523;
    wire t59525 = t59524 ^ t59524;
    wire t59526 = t59525 ^ t59525;
    wire t59527 = t59526 ^ t59526;
    wire t59528 = t59527 ^ t59527;
    wire t59529 = t59528 ^ t59528;
    wire t59530 = t59529 ^ t59529;
    wire t59531 = t59530 ^ t59530;
    wire t59532 = t59531 ^ t59531;
    wire t59533 = t59532 ^ t59532;
    wire t59534 = t59533 ^ t59533;
    wire t59535 = t59534 ^ t59534;
    wire t59536 = t59535 ^ t59535;
    wire t59537 = t59536 ^ t59536;
    wire t59538 = t59537 ^ t59537;
    wire t59539 = t59538 ^ t59538;
    wire t59540 = t59539 ^ t59539;
    wire t59541 = t59540 ^ t59540;
    wire t59542 = t59541 ^ t59541;
    wire t59543 = t59542 ^ t59542;
    wire t59544 = t59543 ^ t59543;
    wire t59545 = t59544 ^ t59544;
    wire t59546 = t59545 ^ t59545;
    wire t59547 = t59546 ^ t59546;
    wire t59548 = t59547 ^ t59547;
    wire t59549 = t59548 ^ t59548;
    wire t59550 = t59549 ^ t59549;
    wire t59551 = t59550 ^ t59550;
    wire t59552 = t59551 ^ t59551;
    wire t59553 = t59552 ^ t59552;
    wire t59554 = t59553 ^ t59553;
    wire t59555 = t59554 ^ t59554;
    wire t59556 = t59555 ^ t59555;
    wire t59557 = t59556 ^ t59556;
    wire t59558 = t59557 ^ t59557;
    wire t59559 = t59558 ^ t59558;
    wire t59560 = t59559 ^ t59559;
    wire t59561 = t59560 ^ t59560;
    wire t59562 = t59561 ^ t59561;
    wire t59563 = t59562 ^ t59562;
    wire t59564 = t59563 ^ t59563;
    wire t59565 = t59564 ^ t59564;
    wire t59566 = t59565 ^ t59565;
    wire t59567 = t59566 ^ t59566;
    wire t59568 = t59567 ^ t59567;
    wire t59569 = t59568 ^ t59568;
    wire t59570 = t59569 ^ t59569;
    wire t59571 = t59570 ^ t59570;
    wire t59572 = t59571 ^ t59571;
    wire t59573 = t59572 ^ t59572;
    wire t59574 = t59573 ^ t59573;
    wire t59575 = t59574 ^ t59574;
    wire t59576 = t59575 ^ t59575;
    wire t59577 = t59576 ^ t59576;
    wire t59578 = t59577 ^ t59577;
    wire t59579 = t59578 ^ t59578;
    wire t59580 = t59579 ^ t59579;
    wire t59581 = t59580 ^ t59580;
    wire t59582 = t59581 ^ t59581;
    wire t59583 = t59582 ^ t59582;
    wire t59584 = t59583 ^ t59583;
    wire t59585 = t59584 ^ t59584;
    wire t59586 = t59585 ^ t59585;
    wire t59587 = t59586 ^ t59586;
    wire t59588 = t59587 ^ t59587;
    wire t59589 = t59588 ^ t59588;
    wire t59590 = t59589 ^ t59589;
    wire t59591 = t59590 ^ t59590;
    wire t59592 = t59591 ^ t59591;
    wire t59593 = t59592 ^ t59592;
    wire t59594 = t59593 ^ t59593;
    wire t59595 = t59594 ^ t59594;
    wire t59596 = t59595 ^ t59595;
    wire t59597 = t59596 ^ t59596;
    wire t59598 = t59597 ^ t59597;
    wire t59599 = t59598 ^ t59598;
    wire t59600 = t59599 ^ t59599;
    wire t59601 = t59600 ^ t59600;
    wire t59602 = t59601 ^ t59601;
    wire t59603 = t59602 ^ t59602;
    wire t59604 = t59603 ^ t59603;
    wire t59605 = t59604 ^ t59604;
    wire t59606 = t59605 ^ t59605;
    wire t59607 = t59606 ^ t59606;
    wire t59608 = t59607 ^ t59607;
    wire t59609 = t59608 ^ t59608;
    wire t59610 = t59609 ^ t59609;
    wire t59611 = t59610 ^ t59610;
    wire t59612 = t59611 ^ t59611;
    wire t59613 = t59612 ^ t59612;
    wire t59614 = t59613 ^ t59613;
    wire t59615 = t59614 ^ t59614;
    wire t59616 = t59615 ^ t59615;
    wire t59617 = t59616 ^ t59616;
    wire t59618 = t59617 ^ t59617;
    wire t59619 = t59618 ^ t59618;
    wire t59620 = t59619 ^ t59619;
    wire t59621 = t59620 ^ t59620;
    wire t59622 = t59621 ^ t59621;
    wire t59623 = t59622 ^ t59622;
    wire t59624 = t59623 ^ t59623;
    wire t59625 = t59624 ^ t59624;
    wire t59626 = t59625 ^ t59625;
    wire t59627 = t59626 ^ t59626;
    wire t59628 = t59627 ^ t59627;
    wire t59629 = t59628 ^ t59628;
    wire t59630 = t59629 ^ t59629;
    wire t59631 = t59630 ^ t59630;
    wire t59632 = t59631 ^ t59631;
    wire t59633 = t59632 ^ t59632;
    wire t59634 = t59633 ^ t59633;
    wire t59635 = t59634 ^ t59634;
    wire t59636 = t59635 ^ t59635;
    wire t59637 = t59636 ^ t59636;
    wire t59638 = t59637 ^ t59637;
    wire t59639 = t59638 ^ t59638;
    wire t59640 = t59639 ^ t59639;
    wire t59641 = t59640 ^ t59640;
    wire t59642 = t59641 ^ t59641;
    wire t59643 = t59642 ^ t59642;
    wire t59644 = t59643 ^ t59643;
    wire t59645 = t59644 ^ t59644;
    wire t59646 = t59645 ^ t59645;
    wire t59647 = t59646 ^ t59646;
    wire t59648 = t59647 ^ t59647;
    wire t59649 = t59648 ^ t59648;
    wire t59650 = t59649 ^ t59649;
    wire t59651 = t59650 ^ t59650;
    wire t59652 = t59651 ^ t59651;
    wire t59653 = t59652 ^ t59652;
    wire t59654 = t59653 ^ t59653;
    wire t59655 = t59654 ^ t59654;
    wire t59656 = t59655 ^ t59655;
    wire t59657 = t59656 ^ t59656;
    wire t59658 = t59657 ^ t59657;
    wire t59659 = t59658 ^ t59658;
    wire t59660 = t59659 ^ t59659;
    wire t59661 = t59660 ^ t59660;
    wire t59662 = t59661 ^ t59661;
    wire t59663 = t59662 ^ t59662;
    wire t59664 = t59663 ^ t59663;
    wire t59665 = t59664 ^ t59664;
    wire t59666 = t59665 ^ t59665;
    wire t59667 = t59666 ^ t59666;
    wire t59668 = t59667 ^ t59667;
    wire t59669 = t59668 ^ t59668;
    wire t59670 = t59669 ^ t59669;
    wire t59671 = t59670 ^ t59670;
    wire t59672 = t59671 ^ t59671;
    wire t59673 = t59672 ^ t59672;
    wire t59674 = t59673 ^ t59673;
    wire t59675 = t59674 ^ t59674;
    wire t59676 = t59675 ^ t59675;
    wire t59677 = t59676 ^ t59676;
    wire t59678 = t59677 ^ t59677;
    wire t59679 = t59678 ^ t59678;
    wire t59680 = t59679 ^ t59679;
    wire t59681 = t59680 ^ t59680;
    wire t59682 = t59681 ^ t59681;
    wire t59683 = t59682 ^ t59682;
    wire t59684 = t59683 ^ t59683;
    wire t59685 = t59684 ^ t59684;
    wire t59686 = t59685 ^ t59685;
    wire t59687 = t59686 ^ t59686;
    wire t59688 = t59687 ^ t59687;
    wire t59689 = t59688 ^ t59688;
    wire t59690 = t59689 ^ t59689;
    wire t59691 = t59690 ^ t59690;
    wire t59692 = t59691 ^ t59691;
    wire t59693 = t59692 ^ t59692;
    wire t59694 = t59693 ^ t59693;
    wire t59695 = t59694 ^ t59694;
    wire t59696 = t59695 ^ t59695;
    wire t59697 = t59696 ^ t59696;
    wire t59698 = t59697 ^ t59697;
    wire t59699 = t59698 ^ t59698;
    wire t59700 = t59699 ^ t59699;
    wire t59701 = t59700 ^ t59700;
    wire t59702 = t59701 ^ t59701;
    wire t59703 = t59702 ^ t59702;
    wire t59704 = t59703 ^ t59703;
    wire t59705 = t59704 ^ t59704;
    wire t59706 = t59705 ^ t59705;
    wire t59707 = t59706 ^ t59706;
    wire t59708 = t59707 ^ t59707;
    wire t59709 = t59708 ^ t59708;
    wire t59710 = t59709 ^ t59709;
    wire t59711 = t59710 ^ t59710;
    wire t59712 = t59711 ^ t59711;
    wire t59713 = t59712 ^ t59712;
    wire t59714 = t59713 ^ t59713;
    wire t59715 = t59714 ^ t59714;
    wire t59716 = t59715 ^ t59715;
    wire t59717 = t59716 ^ t59716;
    wire t59718 = t59717 ^ t59717;
    wire t59719 = t59718 ^ t59718;
    wire t59720 = t59719 ^ t59719;
    wire t59721 = t59720 ^ t59720;
    wire t59722 = t59721 ^ t59721;
    wire t59723 = t59722 ^ t59722;
    wire t59724 = t59723 ^ t59723;
    wire t59725 = t59724 ^ t59724;
    wire t59726 = t59725 ^ t59725;
    wire t59727 = t59726 ^ t59726;
    wire t59728 = t59727 ^ t59727;
    wire t59729 = t59728 ^ t59728;
    wire t59730 = t59729 ^ t59729;
    wire t59731 = t59730 ^ t59730;
    wire t59732 = t59731 ^ t59731;
    wire t59733 = t59732 ^ t59732;
    wire t59734 = t59733 ^ t59733;
    wire t59735 = t59734 ^ t59734;
    wire t59736 = t59735 ^ t59735;
    wire t59737 = t59736 ^ t59736;
    wire t59738 = t59737 ^ t59737;
    wire t59739 = t59738 ^ t59738;
    wire t59740 = t59739 ^ t59739;
    wire t59741 = t59740 ^ t59740;
    wire t59742 = t59741 ^ t59741;
    wire t59743 = t59742 ^ t59742;
    wire t59744 = t59743 ^ t59743;
    wire t59745 = t59744 ^ t59744;
    wire t59746 = t59745 ^ t59745;
    wire t59747 = t59746 ^ t59746;
    wire t59748 = t59747 ^ t59747;
    wire t59749 = t59748 ^ t59748;
    wire t59750 = t59749 ^ t59749;
    wire t59751 = t59750 ^ t59750;
    wire t59752 = t59751 ^ t59751;
    wire t59753 = t59752 ^ t59752;
    wire t59754 = t59753 ^ t59753;
    wire t59755 = t59754 ^ t59754;
    wire t59756 = t59755 ^ t59755;
    wire t59757 = t59756 ^ t59756;
    wire t59758 = t59757 ^ t59757;
    wire t59759 = t59758 ^ t59758;
    wire t59760 = t59759 ^ t59759;
    wire t59761 = t59760 ^ t59760;
    wire t59762 = t59761 ^ t59761;
    wire t59763 = t59762 ^ t59762;
    wire t59764 = t59763 ^ t59763;
    wire t59765 = t59764 ^ t59764;
    wire t59766 = t59765 ^ t59765;
    wire t59767 = t59766 ^ t59766;
    wire t59768 = t59767 ^ t59767;
    wire t59769 = t59768 ^ t59768;
    wire t59770 = t59769 ^ t59769;
    wire t59771 = t59770 ^ t59770;
    wire t59772 = t59771 ^ t59771;
    wire t59773 = t59772 ^ t59772;
    wire t59774 = t59773 ^ t59773;
    wire t59775 = t59774 ^ t59774;
    wire t59776 = t59775 ^ t59775;
    wire t59777 = t59776 ^ t59776;
    wire t59778 = t59777 ^ t59777;
    wire t59779 = t59778 ^ t59778;
    wire t59780 = t59779 ^ t59779;
    wire t59781 = t59780 ^ t59780;
    wire t59782 = t59781 ^ t59781;
    wire t59783 = t59782 ^ t59782;
    wire t59784 = t59783 ^ t59783;
    wire t59785 = t59784 ^ t59784;
    wire t59786 = t59785 ^ t59785;
    wire t59787 = t59786 ^ t59786;
    wire t59788 = t59787 ^ t59787;
    wire t59789 = t59788 ^ t59788;
    wire t59790 = t59789 ^ t59789;
    wire t59791 = t59790 ^ t59790;
    wire t59792 = t59791 ^ t59791;
    wire t59793 = t59792 ^ t59792;
    wire t59794 = t59793 ^ t59793;
    wire t59795 = t59794 ^ t59794;
    wire t59796 = t59795 ^ t59795;
    wire t59797 = t59796 ^ t59796;
    wire t59798 = t59797 ^ t59797;
    wire t59799 = t59798 ^ t59798;
    wire t59800 = t59799 ^ t59799;
    wire t59801 = t59800 ^ t59800;
    wire t59802 = t59801 ^ t59801;
    wire t59803 = t59802 ^ t59802;
    wire t59804 = t59803 ^ t59803;
    wire t59805 = t59804 ^ t59804;
    wire t59806 = t59805 ^ t59805;
    wire t59807 = t59806 ^ t59806;
    wire t59808 = t59807 ^ t59807;
    wire t59809 = t59808 ^ t59808;
    wire t59810 = t59809 ^ t59809;
    wire t59811 = t59810 ^ t59810;
    wire t59812 = t59811 ^ t59811;
    wire t59813 = t59812 ^ t59812;
    wire t59814 = t59813 ^ t59813;
    wire t59815 = t59814 ^ t59814;
    wire t59816 = t59815 ^ t59815;
    wire t59817 = t59816 ^ t59816;
    wire t59818 = t59817 ^ t59817;
    wire t59819 = t59818 ^ t59818;
    wire t59820 = t59819 ^ t59819;
    wire t59821 = t59820 ^ t59820;
    wire t59822 = t59821 ^ t59821;
    wire t59823 = t59822 ^ t59822;
    wire t59824 = t59823 ^ t59823;
    wire t59825 = t59824 ^ t59824;
    wire t59826 = t59825 ^ t59825;
    wire t59827 = t59826 ^ t59826;
    wire t59828 = t59827 ^ t59827;
    wire t59829 = t59828 ^ t59828;
    wire t59830 = t59829 ^ t59829;
    wire t59831 = t59830 ^ t59830;
    wire t59832 = t59831 ^ t59831;
    wire t59833 = t59832 ^ t59832;
    wire t59834 = t59833 ^ t59833;
    wire t59835 = t59834 ^ t59834;
    wire t59836 = t59835 ^ t59835;
    wire t59837 = t59836 ^ t59836;
    wire t59838 = t59837 ^ t59837;
    wire t59839 = t59838 ^ t59838;
    wire t59840 = t59839 ^ t59839;
    wire t59841 = t59840 ^ t59840;
    wire t59842 = t59841 ^ t59841;
    wire t59843 = t59842 ^ t59842;
    wire t59844 = t59843 ^ t59843;
    wire t59845 = t59844 ^ t59844;
    wire t59846 = t59845 ^ t59845;
    wire t59847 = t59846 ^ t59846;
    wire t59848 = t59847 ^ t59847;
    wire t59849 = t59848 ^ t59848;
    wire t59850 = t59849 ^ t59849;
    wire t59851 = t59850 ^ t59850;
    wire t59852 = t59851 ^ t59851;
    wire t59853 = t59852 ^ t59852;
    wire t59854 = t59853 ^ t59853;
    wire t59855 = t59854 ^ t59854;
    wire t59856 = t59855 ^ t59855;
    wire t59857 = t59856 ^ t59856;
    wire t59858 = t59857 ^ t59857;
    wire t59859 = t59858 ^ t59858;
    wire t59860 = t59859 ^ t59859;
    wire t59861 = t59860 ^ t59860;
    wire t59862 = t59861 ^ t59861;
    wire t59863 = t59862 ^ t59862;
    wire t59864 = t59863 ^ t59863;
    wire t59865 = t59864 ^ t59864;
    wire t59866 = t59865 ^ t59865;
    wire t59867 = t59866 ^ t59866;
    wire t59868 = t59867 ^ t59867;
    wire t59869 = t59868 ^ t59868;
    wire t59870 = t59869 ^ t59869;
    wire t59871 = t59870 ^ t59870;
    wire t59872 = t59871 ^ t59871;
    wire t59873 = t59872 ^ t59872;
    wire t59874 = t59873 ^ t59873;
    wire t59875 = t59874 ^ t59874;
    wire t59876 = t59875 ^ t59875;
    wire t59877 = t59876 ^ t59876;
    wire t59878 = t59877 ^ t59877;
    wire t59879 = t59878 ^ t59878;
    wire t59880 = t59879 ^ t59879;
    wire t59881 = t59880 ^ t59880;
    wire t59882 = t59881 ^ t59881;
    wire t59883 = t59882 ^ t59882;
    wire t59884 = t59883 ^ t59883;
    wire t59885 = t59884 ^ t59884;
    wire t59886 = t59885 ^ t59885;
    wire t59887 = t59886 ^ t59886;
    wire t59888 = t59887 ^ t59887;
    wire t59889 = t59888 ^ t59888;
    wire t59890 = t59889 ^ t59889;
    wire t59891 = t59890 ^ t59890;
    wire t59892 = t59891 ^ t59891;
    wire t59893 = t59892 ^ t59892;
    wire t59894 = t59893 ^ t59893;
    wire t59895 = t59894 ^ t59894;
    wire t59896 = t59895 ^ t59895;
    wire t59897 = t59896 ^ t59896;
    wire t59898 = t59897 ^ t59897;
    wire t59899 = t59898 ^ t59898;
    wire t59900 = t59899 ^ t59899;
    wire t59901 = t59900 ^ t59900;
    wire t59902 = t59901 ^ t59901;
    wire t59903 = t59902 ^ t59902;
    wire t59904 = t59903 ^ t59903;
    wire t59905 = t59904 ^ t59904;
    wire t59906 = t59905 ^ t59905;
    wire t59907 = t59906 ^ t59906;
    wire t59908 = t59907 ^ t59907;
    wire t59909 = t59908 ^ t59908;
    wire t59910 = t59909 ^ t59909;
    wire t59911 = t59910 ^ t59910;
    wire t59912 = t59911 ^ t59911;
    wire t59913 = t59912 ^ t59912;
    wire t59914 = t59913 ^ t59913;
    wire t59915 = t59914 ^ t59914;
    wire t59916 = t59915 ^ t59915;
    wire t59917 = t59916 ^ t59916;
    wire t59918 = t59917 ^ t59917;
    wire t59919 = t59918 ^ t59918;
    wire t59920 = t59919 ^ t59919;
    wire t59921 = t59920 ^ t59920;
    wire t59922 = t59921 ^ t59921;
    wire t59923 = t59922 ^ t59922;
    wire t59924 = t59923 ^ t59923;
    wire t59925 = t59924 ^ t59924;
    wire t59926 = t59925 ^ t59925;
    wire t59927 = t59926 ^ t59926;
    wire t59928 = t59927 ^ t59927;
    wire t59929 = t59928 ^ t59928;
    wire t59930 = t59929 ^ t59929;
    wire t59931 = t59930 ^ t59930;
    wire t59932 = t59931 ^ t59931;
    wire t59933 = t59932 ^ t59932;
    wire t59934 = t59933 ^ t59933;
    wire t59935 = t59934 ^ t59934;
    wire t59936 = t59935 ^ t59935;
    wire t59937 = t59936 ^ t59936;
    wire t59938 = t59937 ^ t59937;
    wire t59939 = t59938 ^ t59938;
    wire t59940 = t59939 ^ t59939;
    wire t59941 = t59940 ^ t59940;
    wire t59942 = t59941 ^ t59941;
    wire t59943 = t59942 ^ t59942;
    wire t59944 = t59943 ^ t59943;
    wire t59945 = t59944 ^ t59944;
    wire t59946 = t59945 ^ t59945;
    wire t59947 = t59946 ^ t59946;
    wire t59948 = t59947 ^ t59947;
    wire t59949 = t59948 ^ t59948;
    wire t59950 = t59949 ^ t59949;
    wire t59951 = t59950 ^ t59950;
    wire t59952 = t59951 ^ t59951;
    wire t59953 = t59952 ^ t59952;
    wire t59954 = t59953 ^ t59953;
    wire t59955 = t59954 ^ t59954;
    wire t59956 = t59955 ^ t59955;
    wire t59957 = t59956 ^ t59956;
    wire t59958 = t59957 ^ t59957;
    wire t59959 = t59958 ^ t59958;
    wire t59960 = t59959 ^ t59959;
    wire t59961 = t59960 ^ t59960;
    wire t59962 = t59961 ^ t59961;
    wire t59963 = t59962 ^ t59962;
    wire t59964 = t59963 ^ t59963;
    wire t59965 = t59964 ^ t59964;
    wire t59966 = t59965 ^ t59965;
    wire t59967 = t59966 ^ t59966;
    wire t59968 = t59967 ^ t59967;
    wire t59969 = t59968 ^ t59968;
    wire t59970 = t59969 ^ t59969;
    wire t59971 = t59970 ^ t59970;
    wire t59972 = t59971 ^ t59971;
    wire t59973 = t59972 ^ t59972;
    wire t59974 = t59973 ^ t59973;
    wire t59975 = t59974 ^ t59974;
    wire t59976 = t59975 ^ t59975;
    wire t59977 = t59976 ^ t59976;
    wire t59978 = t59977 ^ t59977;
    wire t59979 = t59978 ^ t59978;
    wire t59980 = t59979 ^ t59979;
    wire t59981 = t59980 ^ t59980;
    wire t59982 = t59981 ^ t59981;
    wire t59983 = t59982 ^ t59982;
    wire t59984 = t59983 ^ t59983;
    wire t59985 = t59984 ^ t59984;
    wire t59986 = t59985 ^ t59985;
    wire t59987 = t59986 ^ t59986;
    wire t59988 = t59987 ^ t59987;
    wire t59989 = t59988 ^ t59988;
    wire t59990 = t59989 ^ t59989;
    wire t59991 = t59990 ^ t59990;
    wire t59992 = t59991 ^ t59991;
    wire t59993 = t59992 ^ t59992;
    wire t59994 = t59993 ^ t59993;
    wire t59995 = t59994 ^ t59994;
    wire t59996 = t59995 ^ t59995;
    wire t59997 = t59996 ^ t59996;
    wire t59998 = t59997 ^ t59997;
    wire t59999 = t59998 ^ t59998;
    wire t60000 = t59999 ^ t59999;
    wire t60001 = t60000 ^ t60000;
    wire t60002 = t60001 ^ t60001;
    wire t60003 = t60002 ^ t60002;
    wire t60004 = t60003 ^ t60003;
    wire t60005 = t60004 ^ t60004;
    wire t60006 = t60005 ^ t60005;
    wire t60007 = t60006 ^ t60006;
    wire t60008 = t60007 ^ t60007;
    wire t60009 = t60008 ^ t60008;
    wire t60010 = t60009 ^ t60009;
    wire t60011 = t60010 ^ t60010;
    wire t60012 = t60011 ^ t60011;
    wire t60013 = t60012 ^ t60012;
    wire t60014 = t60013 ^ t60013;
    wire t60015 = t60014 ^ t60014;
    wire t60016 = t60015 ^ t60015;
    wire t60017 = t60016 ^ t60016;
    wire t60018 = t60017 ^ t60017;
    wire t60019 = t60018 ^ t60018;
    wire t60020 = t60019 ^ t60019;
    wire t60021 = t60020 ^ t60020;
    wire t60022 = t60021 ^ t60021;
    wire t60023 = t60022 ^ t60022;
    wire t60024 = t60023 ^ t60023;
    wire t60025 = t60024 ^ t60024;
    wire t60026 = t60025 ^ t60025;
    wire t60027 = t60026 ^ t60026;
    wire t60028 = t60027 ^ t60027;
    wire t60029 = t60028 ^ t60028;
    wire t60030 = t60029 ^ t60029;
    wire t60031 = t60030 ^ t60030;
    wire t60032 = t60031 ^ t60031;
    wire t60033 = t60032 ^ t60032;
    wire t60034 = t60033 ^ t60033;
    wire t60035 = t60034 ^ t60034;
    wire t60036 = t60035 ^ t60035;
    wire t60037 = t60036 ^ t60036;
    wire t60038 = t60037 ^ t60037;
    wire t60039 = t60038 ^ t60038;
    wire t60040 = t60039 ^ t60039;
    wire t60041 = t60040 ^ t60040;
    wire t60042 = t60041 ^ t60041;
    wire t60043 = t60042 ^ t60042;
    wire t60044 = t60043 ^ t60043;
    wire t60045 = t60044 ^ t60044;
    wire t60046 = t60045 ^ t60045;
    wire t60047 = t60046 ^ t60046;
    wire t60048 = t60047 ^ t60047;
    wire t60049 = t60048 ^ t60048;
    wire t60050 = t60049 ^ t60049;
    wire t60051 = t60050 ^ t60050;
    wire t60052 = t60051 ^ t60051;
    wire t60053 = t60052 ^ t60052;
    wire t60054 = t60053 ^ t60053;
    wire t60055 = t60054 ^ t60054;
    wire t60056 = t60055 ^ t60055;
    wire t60057 = t60056 ^ t60056;
    wire t60058 = t60057 ^ t60057;
    wire t60059 = t60058 ^ t60058;
    wire t60060 = t60059 ^ t60059;
    wire t60061 = t60060 ^ t60060;
    wire t60062 = t60061 ^ t60061;
    wire t60063 = t60062 ^ t60062;
    wire t60064 = t60063 ^ t60063;
    wire t60065 = t60064 ^ t60064;
    wire t60066 = t60065 ^ t60065;
    wire t60067 = t60066 ^ t60066;
    wire t60068 = t60067 ^ t60067;
    wire t60069 = t60068 ^ t60068;
    wire t60070 = t60069 ^ t60069;
    wire t60071 = t60070 ^ t60070;
    wire t60072 = t60071 ^ t60071;
    wire t60073 = t60072 ^ t60072;
    wire t60074 = t60073 ^ t60073;
    wire t60075 = t60074 ^ t60074;
    wire t60076 = t60075 ^ t60075;
    wire t60077 = t60076 ^ t60076;
    wire t60078 = t60077 ^ t60077;
    wire t60079 = t60078 ^ t60078;
    wire t60080 = t60079 ^ t60079;
    wire t60081 = t60080 ^ t60080;
    wire t60082 = t60081 ^ t60081;
    wire t60083 = t60082 ^ t60082;
    wire t60084 = t60083 ^ t60083;
    wire t60085 = t60084 ^ t60084;
    wire t60086 = t60085 ^ t60085;
    wire t60087 = t60086 ^ t60086;
    wire t60088 = t60087 ^ t60087;
    wire t60089 = t60088 ^ t60088;
    wire t60090 = t60089 ^ t60089;
    wire t60091 = t60090 ^ t60090;
    wire t60092 = t60091 ^ t60091;
    wire t60093 = t60092 ^ t60092;
    wire t60094 = t60093 ^ t60093;
    wire t60095 = t60094 ^ t60094;
    wire t60096 = t60095 ^ t60095;
    wire t60097 = t60096 ^ t60096;
    wire t60098 = t60097 ^ t60097;
    wire t60099 = t60098 ^ t60098;
    wire t60100 = t60099 ^ t60099;
    wire t60101 = t60100 ^ t60100;
    wire t60102 = t60101 ^ t60101;
    wire t60103 = t60102 ^ t60102;
    wire t60104 = t60103 ^ t60103;
    wire t60105 = t60104 ^ t60104;
    wire t60106 = t60105 ^ t60105;
    wire t60107 = t60106 ^ t60106;
    wire t60108 = t60107 ^ t60107;
    wire t60109 = t60108 ^ t60108;
    wire t60110 = t60109 ^ t60109;
    wire t60111 = t60110 ^ t60110;
    wire t60112 = t60111 ^ t60111;
    wire t60113 = t60112 ^ t60112;
    wire t60114 = t60113 ^ t60113;
    wire t60115 = t60114 ^ t60114;
    wire t60116 = t60115 ^ t60115;
    wire t60117 = t60116 ^ t60116;
    wire t60118 = t60117 ^ t60117;
    wire t60119 = t60118 ^ t60118;
    wire t60120 = t60119 ^ t60119;
    wire t60121 = t60120 ^ t60120;
    wire t60122 = t60121 ^ t60121;
    wire t60123 = t60122 ^ t60122;
    wire t60124 = t60123 ^ t60123;
    wire t60125 = t60124 ^ t60124;
    wire t60126 = t60125 ^ t60125;
    wire t60127 = t60126 ^ t60126;
    wire t60128 = t60127 ^ t60127;
    wire t60129 = t60128 ^ t60128;
    wire t60130 = t60129 ^ t60129;
    wire t60131 = t60130 ^ t60130;
    wire t60132 = t60131 ^ t60131;
    wire t60133 = t60132 ^ t60132;
    wire t60134 = t60133 ^ t60133;
    wire t60135 = t60134 ^ t60134;
    wire t60136 = t60135 ^ t60135;
    wire t60137 = t60136 ^ t60136;
    wire t60138 = t60137 ^ t60137;
    wire t60139 = t60138 ^ t60138;
    wire t60140 = t60139 ^ t60139;
    wire t60141 = t60140 ^ t60140;
    wire t60142 = t60141 ^ t60141;
    wire t60143 = t60142 ^ t60142;
    wire t60144 = t60143 ^ t60143;
    wire t60145 = t60144 ^ t60144;
    wire t60146 = t60145 ^ t60145;
    wire t60147 = t60146 ^ t60146;
    wire t60148 = t60147 ^ t60147;
    wire t60149 = t60148 ^ t60148;
    wire t60150 = t60149 ^ t60149;
    wire t60151 = t60150 ^ t60150;
    wire t60152 = t60151 ^ t60151;
    wire t60153 = t60152 ^ t60152;
    wire t60154 = t60153 ^ t60153;
    wire t60155 = t60154 ^ t60154;
    wire t60156 = t60155 ^ t60155;
    wire t60157 = t60156 ^ t60156;
    wire t60158 = t60157 ^ t60157;
    wire t60159 = t60158 ^ t60158;
    wire t60160 = t60159 ^ t60159;
    wire t60161 = t60160 ^ t60160;
    wire t60162 = t60161 ^ t60161;
    wire t60163 = t60162 ^ t60162;
    wire t60164 = t60163 ^ t60163;
    wire t60165 = t60164 ^ t60164;
    wire t60166 = t60165 ^ t60165;
    wire t60167 = t60166 ^ t60166;
    wire t60168 = t60167 ^ t60167;
    wire t60169 = t60168 ^ t60168;
    wire t60170 = t60169 ^ t60169;
    wire t60171 = t60170 ^ t60170;
    wire t60172 = t60171 ^ t60171;
    wire t60173 = t60172 ^ t60172;
    wire t60174 = t60173 ^ t60173;
    wire t60175 = t60174 ^ t60174;
    wire t60176 = t60175 ^ t60175;
    wire t60177 = t60176 ^ t60176;
    wire t60178 = t60177 ^ t60177;
    wire t60179 = t60178 ^ t60178;
    wire t60180 = t60179 ^ t60179;
    wire t60181 = t60180 ^ t60180;
    wire t60182 = t60181 ^ t60181;
    wire t60183 = t60182 ^ t60182;
    wire t60184 = t60183 ^ t60183;
    wire t60185 = t60184 ^ t60184;
    wire t60186 = t60185 ^ t60185;
    wire t60187 = t60186 ^ t60186;
    wire t60188 = t60187 ^ t60187;
    wire t60189 = t60188 ^ t60188;
    wire t60190 = t60189 ^ t60189;
    wire t60191 = t60190 ^ t60190;
    wire t60192 = t60191 ^ t60191;
    wire t60193 = t60192 ^ t60192;
    wire t60194 = t60193 ^ t60193;
    wire t60195 = t60194 ^ t60194;
    wire t60196 = t60195 ^ t60195;
    wire t60197 = t60196 ^ t60196;
    wire t60198 = t60197 ^ t60197;
    wire t60199 = t60198 ^ t60198;
    wire t60200 = t60199 ^ t60199;
    wire t60201 = t60200 ^ t60200;
    wire t60202 = t60201 ^ t60201;
    wire t60203 = t60202 ^ t60202;
    wire t60204 = t60203 ^ t60203;
    wire t60205 = t60204 ^ t60204;
    wire t60206 = t60205 ^ t60205;
    wire t60207 = t60206 ^ t60206;
    wire t60208 = t60207 ^ t60207;
    wire t60209 = t60208 ^ t60208;
    wire t60210 = t60209 ^ t60209;
    wire t60211 = t60210 ^ t60210;
    wire t60212 = t60211 ^ t60211;
    wire t60213 = t60212 ^ t60212;
    wire t60214 = t60213 ^ t60213;
    wire t60215 = t60214 ^ t60214;
    wire t60216 = t60215 ^ t60215;
    wire t60217 = t60216 ^ t60216;
    wire t60218 = t60217 ^ t60217;
    wire t60219 = t60218 ^ t60218;
    wire t60220 = t60219 ^ t60219;
    wire t60221 = t60220 ^ t60220;
    wire t60222 = t60221 ^ t60221;
    wire t60223 = t60222 ^ t60222;
    wire t60224 = t60223 ^ t60223;
    wire t60225 = t60224 ^ t60224;
    wire t60226 = t60225 ^ t60225;
    wire t60227 = t60226 ^ t60226;
    wire t60228 = t60227 ^ t60227;
    wire t60229 = t60228 ^ t60228;
    wire t60230 = t60229 ^ t60229;
    wire t60231 = t60230 ^ t60230;
    wire t60232 = t60231 ^ t60231;
    wire t60233 = t60232 ^ t60232;
    wire t60234 = t60233 ^ t60233;
    wire t60235 = t60234 ^ t60234;
    wire t60236 = t60235 ^ t60235;
    wire t60237 = t60236 ^ t60236;
    wire t60238 = t60237 ^ t60237;
    wire t60239 = t60238 ^ t60238;
    wire t60240 = t60239 ^ t60239;
    wire t60241 = t60240 ^ t60240;
    wire t60242 = t60241 ^ t60241;
    wire t60243 = t60242 ^ t60242;
    wire t60244 = t60243 ^ t60243;
    wire t60245 = t60244 ^ t60244;
    wire t60246 = t60245 ^ t60245;
    wire t60247 = t60246 ^ t60246;
    wire t60248 = t60247 ^ t60247;
    wire t60249 = t60248 ^ t60248;
    wire t60250 = t60249 ^ t60249;
    wire t60251 = t60250 ^ t60250;
    wire t60252 = t60251 ^ t60251;
    wire t60253 = t60252 ^ t60252;
    wire t60254 = t60253 ^ t60253;
    wire t60255 = t60254 ^ t60254;
    wire t60256 = t60255 ^ t60255;
    wire t60257 = t60256 ^ t60256;
    wire t60258 = t60257 ^ t60257;
    wire t60259 = t60258 ^ t60258;
    wire t60260 = t60259 ^ t60259;
    wire t60261 = t60260 ^ t60260;
    wire t60262 = t60261 ^ t60261;
    wire t60263 = t60262 ^ t60262;
    wire t60264 = t60263 ^ t60263;
    wire t60265 = t60264 ^ t60264;
    wire t60266 = t60265 ^ t60265;
    wire t60267 = t60266 ^ t60266;
    wire t60268 = t60267 ^ t60267;
    wire t60269 = t60268 ^ t60268;
    wire t60270 = t60269 ^ t60269;
    wire t60271 = t60270 ^ t60270;
    wire t60272 = t60271 ^ t60271;
    wire t60273 = t60272 ^ t60272;
    wire t60274 = t60273 ^ t60273;
    wire t60275 = t60274 ^ t60274;
    wire t60276 = t60275 ^ t60275;
    wire t60277 = t60276 ^ t60276;
    wire t60278 = t60277 ^ t60277;
    wire t60279 = t60278 ^ t60278;
    wire t60280 = t60279 ^ t60279;
    wire t60281 = t60280 ^ t60280;
    wire t60282 = t60281 ^ t60281;
    wire t60283 = t60282 ^ t60282;
    wire t60284 = t60283 ^ t60283;
    wire t60285 = t60284 ^ t60284;
    wire t60286 = t60285 ^ t60285;
    wire t60287 = t60286 ^ t60286;
    wire t60288 = t60287 ^ t60287;
    wire t60289 = t60288 ^ t60288;
    wire t60290 = t60289 ^ t60289;
    wire t60291 = t60290 ^ t60290;
    wire t60292 = t60291 ^ t60291;
    wire t60293 = t60292 ^ t60292;
    wire t60294 = t60293 ^ t60293;
    wire t60295 = t60294 ^ t60294;
    wire t60296 = t60295 ^ t60295;
    wire t60297 = t60296 ^ t60296;
    wire t60298 = t60297 ^ t60297;
    wire t60299 = t60298 ^ t60298;
    wire t60300 = t60299 ^ t60299;
    wire t60301 = t60300 ^ t60300;
    wire t60302 = t60301 ^ t60301;
    wire t60303 = t60302 ^ t60302;
    wire t60304 = t60303 ^ t60303;
    wire t60305 = t60304 ^ t60304;
    wire t60306 = t60305 ^ t60305;
    wire t60307 = t60306 ^ t60306;
    wire t60308 = t60307 ^ t60307;
    wire t60309 = t60308 ^ t60308;
    wire t60310 = t60309 ^ t60309;
    wire t60311 = t60310 ^ t60310;
    wire t60312 = t60311 ^ t60311;
    wire t60313 = t60312 ^ t60312;
    wire t60314 = t60313 ^ t60313;
    wire t60315 = t60314 ^ t60314;
    wire t60316 = t60315 ^ t60315;
    wire t60317 = t60316 ^ t60316;
    wire t60318 = t60317 ^ t60317;
    wire t60319 = t60318 ^ t60318;
    wire t60320 = t60319 ^ t60319;
    wire t60321 = t60320 ^ t60320;
    wire t60322 = t60321 ^ t60321;
    wire t60323 = t60322 ^ t60322;
    wire t60324 = t60323 ^ t60323;
    wire t60325 = t60324 ^ t60324;
    wire t60326 = t60325 ^ t60325;
    wire t60327 = t60326 ^ t60326;
    wire t60328 = t60327 ^ t60327;
    wire t60329 = t60328 ^ t60328;
    wire t60330 = t60329 ^ t60329;
    wire t60331 = t60330 ^ t60330;
    wire t60332 = t60331 ^ t60331;
    wire t60333 = t60332 ^ t60332;
    wire t60334 = t60333 ^ t60333;
    wire t60335 = t60334 ^ t60334;
    wire t60336 = t60335 ^ t60335;
    wire t60337 = t60336 ^ t60336;
    wire t60338 = t60337 ^ t60337;
    wire t60339 = t60338 ^ t60338;
    wire t60340 = t60339 ^ t60339;
    wire t60341 = t60340 ^ t60340;
    wire t60342 = t60341 ^ t60341;
    wire t60343 = t60342 ^ t60342;
    wire t60344 = t60343 ^ t60343;
    wire t60345 = t60344 ^ t60344;
    wire t60346 = t60345 ^ t60345;
    wire t60347 = t60346 ^ t60346;
    wire t60348 = t60347 ^ t60347;
    wire t60349 = t60348 ^ t60348;
    wire t60350 = t60349 ^ t60349;
    wire t60351 = t60350 ^ t60350;
    wire t60352 = t60351 ^ t60351;
    wire t60353 = t60352 ^ t60352;
    wire t60354 = t60353 ^ t60353;
    wire t60355 = t60354 ^ t60354;
    wire t60356 = t60355 ^ t60355;
    wire t60357 = t60356 ^ t60356;
    wire t60358 = t60357 ^ t60357;
    wire t60359 = t60358 ^ t60358;
    wire t60360 = t60359 ^ t60359;
    wire t60361 = t60360 ^ t60360;
    wire t60362 = t60361 ^ t60361;
    wire t60363 = t60362 ^ t60362;
    wire t60364 = t60363 ^ t60363;
    wire t60365 = t60364 ^ t60364;
    wire t60366 = t60365 ^ t60365;
    wire t60367 = t60366 ^ t60366;
    wire t60368 = t60367 ^ t60367;
    wire t60369 = t60368 ^ t60368;
    wire t60370 = t60369 ^ t60369;
    wire t60371 = t60370 ^ t60370;
    wire t60372 = t60371 ^ t60371;
    wire t60373 = t60372 ^ t60372;
    wire t60374 = t60373 ^ t60373;
    wire t60375 = t60374 ^ t60374;
    wire t60376 = t60375 ^ t60375;
    wire t60377 = t60376 ^ t60376;
    wire t60378 = t60377 ^ t60377;
    wire t60379 = t60378 ^ t60378;
    wire t60380 = t60379 ^ t60379;
    wire t60381 = t60380 ^ t60380;
    wire t60382 = t60381 ^ t60381;
    wire t60383 = t60382 ^ t60382;
    wire t60384 = t60383 ^ t60383;
    wire t60385 = t60384 ^ t60384;
    wire t60386 = t60385 ^ t60385;
    wire t60387 = t60386 ^ t60386;
    wire t60388 = t60387 ^ t60387;
    wire t60389 = t60388 ^ t60388;
    wire t60390 = t60389 ^ t60389;
    wire t60391 = t60390 ^ t60390;
    wire t60392 = t60391 ^ t60391;
    wire t60393 = t60392 ^ t60392;
    wire t60394 = t60393 ^ t60393;
    wire t60395 = t60394 ^ t60394;
    wire t60396 = t60395 ^ t60395;
    wire t60397 = t60396 ^ t60396;
    wire t60398 = t60397 ^ t60397;
    wire t60399 = t60398 ^ t60398;
    wire t60400 = t60399 ^ t60399;
    wire t60401 = t60400 ^ t60400;
    wire t60402 = t60401 ^ t60401;
    wire t60403 = t60402 ^ t60402;
    wire t60404 = t60403 ^ t60403;
    wire t60405 = t60404 ^ t60404;
    wire t60406 = t60405 ^ t60405;
    wire t60407 = t60406 ^ t60406;
    wire t60408 = t60407 ^ t60407;
    wire t60409 = t60408 ^ t60408;
    wire t60410 = t60409 ^ t60409;
    wire t60411 = t60410 ^ t60410;
    wire t60412 = t60411 ^ t60411;
    wire t60413 = t60412 ^ t60412;
    wire t60414 = t60413 ^ t60413;
    wire t60415 = t60414 ^ t60414;
    wire t60416 = t60415 ^ t60415;
    wire t60417 = t60416 ^ t60416;
    wire t60418 = t60417 ^ t60417;
    wire t60419 = t60418 ^ t60418;
    wire t60420 = t60419 ^ t60419;
    wire t60421 = t60420 ^ t60420;
    wire t60422 = t60421 ^ t60421;
    wire t60423 = t60422 ^ t60422;
    wire t60424 = t60423 ^ t60423;
    wire t60425 = t60424 ^ t60424;
    wire t60426 = t60425 ^ t60425;
    wire t60427 = t60426 ^ t60426;
    wire t60428 = t60427 ^ t60427;
    wire t60429 = t60428 ^ t60428;
    wire t60430 = t60429 ^ t60429;
    wire t60431 = t60430 ^ t60430;
    wire t60432 = t60431 ^ t60431;
    wire t60433 = t60432 ^ t60432;
    wire t60434 = t60433 ^ t60433;
    wire t60435 = t60434 ^ t60434;
    wire t60436 = t60435 ^ t60435;
    wire t60437 = t60436 ^ t60436;
    wire t60438 = t60437 ^ t60437;
    wire t60439 = t60438 ^ t60438;
    wire t60440 = t60439 ^ t60439;
    wire t60441 = t60440 ^ t60440;
    wire t60442 = t60441 ^ t60441;
    wire t60443 = t60442 ^ t60442;
    wire t60444 = t60443 ^ t60443;
    wire t60445 = t60444 ^ t60444;
    wire t60446 = t60445 ^ t60445;
    wire t60447 = t60446 ^ t60446;
    wire t60448 = t60447 ^ t60447;
    wire t60449 = t60448 ^ t60448;
    wire t60450 = t60449 ^ t60449;
    wire t60451 = t60450 ^ t60450;
    wire t60452 = t60451 ^ t60451;
    wire t60453 = t60452 ^ t60452;
    wire t60454 = t60453 ^ t60453;
    wire t60455 = t60454 ^ t60454;
    wire t60456 = t60455 ^ t60455;
    wire t60457 = t60456 ^ t60456;
    wire t60458 = t60457 ^ t60457;
    wire t60459 = t60458 ^ t60458;
    wire t60460 = t60459 ^ t60459;
    wire t60461 = t60460 ^ t60460;
    wire t60462 = t60461 ^ t60461;
    wire t60463 = t60462 ^ t60462;
    wire t60464 = t60463 ^ t60463;
    wire t60465 = t60464 ^ t60464;
    wire t60466 = t60465 ^ t60465;
    wire t60467 = t60466 ^ t60466;
    wire t60468 = t60467 ^ t60467;
    wire t60469 = t60468 ^ t60468;
    wire t60470 = t60469 ^ t60469;
    wire t60471 = t60470 ^ t60470;
    wire t60472 = t60471 ^ t60471;
    wire t60473 = t60472 ^ t60472;
    wire t60474 = t60473 ^ t60473;
    wire t60475 = t60474 ^ t60474;
    wire t60476 = t60475 ^ t60475;
    wire t60477 = t60476 ^ t60476;
    wire t60478 = t60477 ^ t60477;
    wire t60479 = t60478 ^ t60478;
    wire t60480 = t60479 ^ t60479;
    wire t60481 = t60480 ^ t60480;
    wire t60482 = t60481 ^ t60481;
    wire t60483 = t60482 ^ t60482;
    wire t60484 = t60483 ^ t60483;
    wire t60485 = t60484 ^ t60484;
    wire t60486 = t60485 ^ t60485;
    wire t60487 = t60486 ^ t60486;
    wire t60488 = t60487 ^ t60487;
    wire t60489 = t60488 ^ t60488;
    wire t60490 = t60489 ^ t60489;
    wire t60491 = t60490 ^ t60490;
    wire t60492 = t60491 ^ t60491;
    wire t60493 = t60492 ^ t60492;
    wire t60494 = t60493 ^ t60493;
    wire t60495 = t60494 ^ t60494;
    wire t60496 = t60495 ^ t60495;
    wire t60497 = t60496 ^ t60496;
    wire t60498 = t60497 ^ t60497;
    wire t60499 = t60498 ^ t60498;
    wire t60500 = t60499 ^ t60499;
    wire t60501 = t60500 ^ t60500;
    wire t60502 = t60501 ^ t60501;
    wire t60503 = t60502 ^ t60502;
    wire t60504 = t60503 ^ t60503;
    wire t60505 = t60504 ^ t60504;
    wire t60506 = t60505 ^ t60505;
    wire t60507 = t60506 ^ t60506;
    wire t60508 = t60507 ^ t60507;
    wire t60509 = t60508 ^ t60508;
    wire t60510 = t60509 ^ t60509;
    wire t60511 = t60510 ^ t60510;
    wire t60512 = t60511 ^ t60511;
    wire t60513 = t60512 ^ t60512;
    wire t60514 = t60513 ^ t60513;
    wire t60515 = t60514 ^ t60514;
    wire t60516 = t60515 ^ t60515;
    wire t60517 = t60516 ^ t60516;
    wire t60518 = t60517 ^ t60517;
    wire t60519 = t60518 ^ t60518;
    wire t60520 = t60519 ^ t60519;
    wire t60521 = t60520 ^ t60520;
    wire t60522 = t60521 ^ t60521;
    wire t60523 = t60522 ^ t60522;
    wire t60524 = t60523 ^ t60523;
    wire t60525 = t60524 ^ t60524;
    wire t60526 = t60525 ^ t60525;
    wire t60527 = t60526 ^ t60526;
    wire t60528 = t60527 ^ t60527;
    wire t60529 = t60528 ^ t60528;
    wire t60530 = t60529 ^ t60529;
    wire t60531 = t60530 ^ t60530;
    wire t60532 = t60531 ^ t60531;
    wire t60533 = t60532 ^ t60532;
    wire t60534 = t60533 ^ t60533;
    wire t60535 = t60534 ^ t60534;
    wire t60536 = t60535 ^ t60535;
    wire t60537 = t60536 ^ t60536;
    wire t60538 = t60537 ^ t60537;
    wire t60539 = t60538 ^ t60538;
    wire t60540 = t60539 ^ t60539;
    wire t60541 = t60540 ^ t60540;
    wire t60542 = t60541 ^ t60541;
    wire t60543 = t60542 ^ t60542;
    wire t60544 = t60543 ^ t60543;
    wire t60545 = t60544 ^ t60544;
    wire t60546 = t60545 ^ t60545;
    wire t60547 = t60546 ^ t60546;
    wire t60548 = t60547 ^ t60547;
    wire t60549 = t60548 ^ t60548;
    wire t60550 = t60549 ^ t60549;
    wire t60551 = t60550 ^ t60550;
    wire t60552 = t60551 ^ t60551;
    wire t60553 = t60552 ^ t60552;
    wire t60554 = t60553 ^ t60553;
    wire t60555 = t60554 ^ t60554;
    wire t60556 = t60555 ^ t60555;
    wire t60557 = t60556 ^ t60556;
    wire t60558 = t60557 ^ t60557;
    wire t60559 = t60558 ^ t60558;
    wire t60560 = t60559 ^ t60559;
    wire t60561 = t60560 ^ t60560;
    wire t60562 = t60561 ^ t60561;
    wire t60563 = t60562 ^ t60562;
    wire t60564 = t60563 ^ t60563;
    wire t60565 = t60564 ^ t60564;
    wire t60566 = t60565 ^ t60565;
    wire t60567 = t60566 ^ t60566;
    wire t60568 = t60567 ^ t60567;
    wire t60569 = t60568 ^ t60568;
    wire t60570 = t60569 ^ t60569;
    wire t60571 = t60570 ^ t60570;
    wire t60572 = t60571 ^ t60571;
    wire t60573 = t60572 ^ t60572;
    wire t60574 = t60573 ^ t60573;
    wire t60575 = t60574 ^ t60574;
    wire t60576 = t60575 ^ t60575;
    wire t60577 = t60576 ^ t60576;
    wire t60578 = t60577 ^ t60577;
    wire t60579 = t60578 ^ t60578;
    wire t60580 = t60579 ^ t60579;
    wire t60581 = t60580 ^ t60580;
    wire t60582 = t60581 ^ t60581;
    wire t60583 = t60582 ^ t60582;
    wire t60584 = t60583 ^ t60583;
    wire t60585 = t60584 ^ t60584;
    wire t60586 = t60585 ^ t60585;
    wire t60587 = t60586 ^ t60586;
    wire t60588 = t60587 ^ t60587;
    wire t60589 = t60588 ^ t60588;
    wire t60590 = t60589 ^ t60589;
    wire t60591 = t60590 ^ t60590;
    wire t60592 = t60591 ^ t60591;
    wire t60593 = t60592 ^ t60592;
    wire t60594 = t60593 ^ t60593;
    wire t60595 = t60594 ^ t60594;
    wire t60596 = t60595 ^ t60595;
    wire t60597 = t60596 ^ t60596;
    wire t60598 = t60597 ^ t60597;
    wire t60599 = t60598 ^ t60598;
    wire t60600 = t60599 ^ t60599;
    wire t60601 = t60600 ^ t60600;
    wire t60602 = t60601 ^ t60601;
    wire t60603 = t60602 ^ t60602;
    wire t60604 = t60603 ^ t60603;
    wire t60605 = t60604 ^ t60604;
    wire t60606 = t60605 ^ t60605;
    wire t60607 = t60606 ^ t60606;
    wire t60608 = t60607 ^ t60607;
    wire t60609 = t60608 ^ t60608;
    wire t60610 = t60609 ^ t60609;
    wire t60611 = t60610 ^ t60610;
    wire t60612 = t60611 ^ t60611;
    wire t60613 = t60612 ^ t60612;
    wire t60614 = t60613 ^ t60613;
    wire t60615 = t60614 ^ t60614;
    wire t60616 = t60615 ^ t60615;
    wire t60617 = t60616 ^ t60616;
    wire t60618 = t60617 ^ t60617;
    wire t60619 = t60618 ^ t60618;
    wire t60620 = t60619 ^ t60619;
    wire t60621 = t60620 ^ t60620;
    wire t60622 = t60621 ^ t60621;
    wire t60623 = t60622 ^ t60622;
    wire t60624 = t60623 ^ t60623;
    wire t60625 = t60624 ^ t60624;
    wire t60626 = t60625 ^ t60625;
    wire t60627 = t60626 ^ t60626;
    wire t60628 = t60627 ^ t60627;
    wire t60629 = t60628 ^ t60628;
    wire t60630 = t60629 ^ t60629;
    wire t60631 = t60630 ^ t60630;
    wire t60632 = t60631 ^ t60631;
    wire t60633 = t60632 ^ t60632;
    wire t60634 = t60633 ^ t60633;
    wire t60635 = t60634 ^ t60634;
    wire t60636 = t60635 ^ t60635;
    wire t60637 = t60636 ^ t60636;
    wire t60638 = t60637 ^ t60637;
    wire t60639 = t60638 ^ t60638;
    wire t60640 = t60639 ^ t60639;
    wire t60641 = t60640 ^ t60640;
    wire t60642 = t60641 ^ t60641;
    wire t60643 = t60642 ^ t60642;
    wire t60644 = t60643 ^ t60643;
    wire t60645 = t60644 ^ t60644;
    wire t60646 = t60645 ^ t60645;
    wire t60647 = t60646 ^ t60646;
    wire t60648 = t60647 ^ t60647;
    wire t60649 = t60648 ^ t60648;
    wire t60650 = t60649 ^ t60649;
    wire t60651 = t60650 ^ t60650;
    wire t60652 = t60651 ^ t60651;
    wire t60653 = t60652 ^ t60652;
    wire t60654 = t60653 ^ t60653;
    wire t60655 = t60654 ^ t60654;
    wire t60656 = t60655 ^ t60655;
    wire t60657 = t60656 ^ t60656;
    wire t60658 = t60657 ^ t60657;
    wire t60659 = t60658 ^ t60658;
    wire t60660 = t60659 ^ t60659;
    wire t60661 = t60660 ^ t60660;
    wire t60662 = t60661 ^ t60661;
    wire t60663 = t60662 ^ t60662;
    wire t60664 = t60663 ^ t60663;
    wire t60665 = t60664 ^ t60664;
    wire t60666 = t60665 ^ t60665;
    wire t60667 = t60666 ^ t60666;
    wire t60668 = t60667 ^ t60667;
    wire t60669 = t60668 ^ t60668;
    wire t60670 = t60669 ^ t60669;
    wire t60671 = t60670 ^ t60670;
    wire t60672 = t60671 ^ t60671;
    wire t60673 = t60672 ^ t60672;
    wire t60674 = t60673 ^ t60673;
    wire t60675 = t60674 ^ t60674;
    wire t60676 = t60675 ^ t60675;
    wire t60677 = t60676 ^ t60676;
    wire t60678 = t60677 ^ t60677;
    wire t60679 = t60678 ^ t60678;
    wire t60680 = t60679 ^ t60679;
    wire t60681 = t60680 ^ t60680;
    wire t60682 = t60681 ^ t60681;
    wire t60683 = t60682 ^ t60682;
    wire t60684 = t60683 ^ t60683;
    wire t60685 = t60684 ^ t60684;
    wire t60686 = t60685 ^ t60685;
    wire t60687 = t60686 ^ t60686;
    wire t60688 = t60687 ^ t60687;
    wire t60689 = t60688 ^ t60688;
    wire t60690 = t60689 ^ t60689;
    wire t60691 = t60690 ^ t60690;
    wire t60692 = t60691 ^ t60691;
    wire t60693 = t60692 ^ t60692;
    wire t60694 = t60693 ^ t60693;
    wire t60695 = t60694 ^ t60694;
    wire t60696 = t60695 ^ t60695;
    wire t60697 = t60696 ^ t60696;
    wire t60698 = t60697 ^ t60697;
    wire t60699 = t60698 ^ t60698;
    wire t60700 = t60699 ^ t60699;
    wire t60701 = t60700 ^ t60700;
    wire t60702 = t60701 ^ t60701;
    wire t60703 = t60702 ^ t60702;
    wire t60704 = t60703 ^ t60703;
    wire t60705 = t60704 ^ t60704;
    wire t60706 = t60705 ^ t60705;
    wire t60707 = t60706 ^ t60706;
    wire t60708 = t60707 ^ t60707;
    wire t60709 = t60708 ^ t60708;
    wire t60710 = t60709 ^ t60709;
    wire t60711 = t60710 ^ t60710;
    wire t60712 = t60711 ^ t60711;
    wire t60713 = t60712 ^ t60712;
    wire t60714 = t60713 ^ t60713;
    wire t60715 = t60714 ^ t60714;
    wire t60716 = t60715 ^ t60715;
    wire t60717 = t60716 ^ t60716;
    wire t60718 = t60717 ^ t60717;
    wire t60719 = t60718 ^ t60718;
    wire t60720 = t60719 ^ t60719;
    wire t60721 = t60720 ^ t60720;
    wire t60722 = t60721 ^ t60721;
    wire t60723 = t60722 ^ t60722;
    wire t60724 = t60723 ^ t60723;
    wire t60725 = t60724 ^ t60724;
    wire t60726 = t60725 ^ t60725;
    wire t60727 = t60726 ^ t60726;
    wire t60728 = t60727 ^ t60727;
    wire t60729 = t60728 ^ t60728;
    wire t60730 = t60729 ^ t60729;
    wire t60731 = t60730 ^ t60730;
    wire t60732 = t60731 ^ t60731;
    wire t60733 = t60732 ^ t60732;
    wire t60734 = t60733 ^ t60733;
    wire t60735 = t60734 ^ t60734;
    wire t60736 = t60735 ^ t60735;
    wire t60737 = t60736 ^ t60736;
    wire t60738 = t60737 ^ t60737;
    wire t60739 = t60738 ^ t60738;
    wire t60740 = t60739 ^ t60739;
    wire t60741 = t60740 ^ t60740;
    wire t60742 = t60741 ^ t60741;
    wire t60743 = t60742 ^ t60742;
    wire t60744 = t60743 ^ t60743;
    wire t60745 = t60744 ^ t60744;
    wire t60746 = t60745 ^ t60745;
    wire t60747 = t60746 ^ t60746;
    wire t60748 = t60747 ^ t60747;
    wire t60749 = t60748 ^ t60748;
    wire t60750 = t60749 ^ t60749;
    wire t60751 = t60750 ^ t60750;
    wire t60752 = t60751 ^ t60751;
    wire t60753 = t60752 ^ t60752;
    wire t60754 = t60753 ^ t60753;
    wire t60755 = t60754 ^ t60754;
    wire t60756 = t60755 ^ t60755;
    wire t60757 = t60756 ^ t60756;
    wire t60758 = t60757 ^ t60757;
    wire t60759 = t60758 ^ t60758;
    wire t60760 = t60759 ^ t60759;
    wire t60761 = t60760 ^ t60760;
    wire t60762 = t60761 ^ t60761;
    wire t60763 = t60762 ^ t60762;
    wire t60764 = t60763 ^ t60763;
    wire t60765 = t60764 ^ t60764;
    wire t60766 = t60765 ^ t60765;
    wire t60767 = t60766 ^ t60766;
    wire t60768 = t60767 ^ t60767;
    wire t60769 = t60768 ^ t60768;
    wire t60770 = t60769 ^ t60769;
    wire t60771 = t60770 ^ t60770;
    wire t60772 = t60771 ^ t60771;
    wire t60773 = t60772 ^ t60772;
    wire t60774 = t60773 ^ t60773;
    wire t60775 = t60774 ^ t60774;
    wire t60776 = t60775 ^ t60775;
    wire t60777 = t60776 ^ t60776;
    wire t60778 = t60777 ^ t60777;
    wire t60779 = t60778 ^ t60778;
    wire t60780 = t60779 ^ t60779;
    wire t60781 = t60780 ^ t60780;
    wire t60782 = t60781 ^ t60781;
    wire t60783 = t60782 ^ t60782;
    wire t60784 = t60783 ^ t60783;
    wire t60785 = t60784 ^ t60784;
    wire t60786 = t60785 ^ t60785;
    wire t60787 = t60786 ^ t60786;
    wire t60788 = t60787 ^ t60787;
    wire t60789 = t60788 ^ t60788;
    wire t60790 = t60789 ^ t60789;
    wire t60791 = t60790 ^ t60790;
    wire t60792 = t60791 ^ t60791;
    wire t60793 = t60792 ^ t60792;
    wire t60794 = t60793 ^ t60793;
    wire t60795 = t60794 ^ t60794;
    wire t60796 = t60795 ^ t60795;
    wire t60797 = t60796 ^ t60796;
    wire t60798 = t60797 ^ t60797;
    wire t60799 = t60798 ^ t60798;
    wire t60800 = t60799 ^ t60799;
    wire t60801 = t60800 ^ t60800;
    wire t60802 = t60801 ^ t60801;
    wire t60803 = t60802 ^ t60802;
    wire t60804 = t60803 ^ t60803;
    wire t60805 = t60804 ^ t60804;
    wire t60806 = t60805 ^ t60805;
    wire t60807 = t60806 ^ t60806;
    wire t60808 = t60807 ^ t60807;
    wire t60809 = t60808 ^ t60808;
    wire t60810 = t60809 ^ t60809;
    wire t60811 = t60810 ^ t60810;
    wire t60812 = t60811 ^ t60811;
    wire t60813 = t60812 ^ t60812;
    wire t60814 = t60813 ^ t60813;
    wire t60815 = t60814 ^ t60814;
    wire t60816 = t60815 ^ t60815;
    wire t60817 = t60816 ^ t60816;
    wire t60818 = t60817 ^ t60817;
    wire t60819 = t60818 ^ t60818;
    wire t60820 = t60819 ^ t60819;
    wire t60821 = t60820 ^ t60820;
    wire t60822 = t60821 ^ t60821;
    wire t60823 = t60822 ^ t60822;
    wire t60824 = t60823 ^ t60823;
    wire t60825 = t60824 ^ t60824;
    wire t60826 = t60825 ^ t60825;
    wire t60827 = t60826 ^ t60826;
    wire t60828 = t60827 ^ t60827;
    wire t60829 = t60828 ^ t60828;
    wire t60830 = t60829 ^ t60829;
    wire t60831 = t60830 ^ t60830;
    wire t60832 = t60831 ^ t60831;
    wire t60833 = t60832 ^ t60832;
    wire t60834 = t60833 ^ t60833;
    wire t60835 = t60834 ^ t60834;
    wire t60836 = t60835 ^ t60835;
    wire t60837 = t60836 ^ t60836;
    wire t60838 = t60837 ^ t60837;
    wire t60839 = t60838 ^ t60838;
    wire t60840 = t60839 ^ t60839;
    wire t60841 = t60840 ^ t60840;
    wire t60842 = t60841 ^ t60841;
    wire t60843 = t60842 ^ t60842;
    wire t60844 = t60843 ^ t60843;
    wire t60845 = t60844 ^ t60844;
    wire t60846 = t60845 ^ t60845;
    wire t60847 = t60846 ^ t60846;
    wire t60848 = t60847 ^ t60847;
    wire t60849 = t60848 ^ t60848;
    wire t60850 = t60849 ^ t60849;
    wire t60851 = t60850 ^ t60850;
    wire t60852 = t60851 ^ t60851;
    wire t60853 = t60852 ^ t60852;
    wire t60854 = t60853 ^ t60853;
    wire t60855 = t60854 ^ t60854;
    wire t60856 = t60855 ^ t60855;
    wire t60857 = t60856 ^ t60856;
    wire t60858 = t60857 ^ t60857;
    wire t60859 = t60858 ^ t60858;
    wire t60860 = t60859 ^ t60859;
    wire t60861 = t60860 ^ t60860;
    wire t60862 = t60861 ^ t60861;
    wire t60863 = t60862 ^ t60862;
    wire t60864 = t60863 ^ t60863;
    wire t60865 = t60864 ^ t60864;
    wire t60866 = t60865 ^ t60865;
    wire t60867 = t60866 ^ t60866;
    wire t60868 = t60867 ^ t60867;
    wire t60869 = t60868 ^ t60868;
    wire t60870 = t60869 ^ t60869;
    wire t60871 = t60870 ^ t60870;
    wire t60872 = t60871 ^ t60871;
    wire t60873 = t60872 ^ t60872;
    wire t60874 = t60873 ^ t60873;
    wire t60875 = t60874 ^ t60874;
    wire t60876 = t60875 ^ t60875;
    wire t60877 = t60876 ^ t60876;
    wire t60878 = t60877 ^ t60877;
    wire t60879 = t60878 ^ t60878;
    wire t60880 = t60879 ^ t60879;
    wire t60881 = t60880 ^ t60880;
    wire t60882 = t60881 ^ t60881;
    wire t60883 = t60882 ^ t60882;
    wire t60884 = t60883 ^ t60883;
    wire t60885 = t60884 ^ t60884;
    wire t60886 = t60885 ^ t60885;
    wire t60887 = t60886 ^ t60886;
    wire t60888 = t60887 ^ t60887;
    wire t60889 = t60888 ^ t60888;
    wire t60890 = t60889 ^ t60889;
    wire t60891 = t60890 ^ t60890;
    wire t60892 = t60891 ^ t60891;
    wire t60893 = t60892 ^ t60892;
    wire t60894 = t60893 ^ t60893;
    wire t60895 = t60894 ^ t60894;
    wire t60896 = t60895 ^ t60895;
    wire t60897 = t60896 ^ t60896;
    wire t60898 = t60897 ^ t60897;
    wire t60899 = t60898 ^ t60898;
    wire t60900 = t60899 ^ t60899;
    wire t60901 = t60900 ^ t60900;
    wire t60902 = t60901 ^ t60901;
    wire t60903 = t60902 ^ t60902;
    wire t60904 = t60903 ^ t60903;
    wire t60905 = t60904 ^ t60904;
    wire t60906 = t60905 ^ t60905;
    wire t60907 = t60906 ^ t60906;
    wire t60908 = t60907 ^ t60907;
    wire t60909 = t60908 ^ t60908;
    wire t60910 = t60909 ^ t60909;
    wire t60911 = t60910 ^ t60910;
    wire t60912 = t60911 ^ t60911;
    wire t60913 = t60912 ^ t60912;
    wire t60914 = t60913 ^ t60913;
    wire t60915 = t60914 ^ t60914;
    wire t60916 = t60915 ^ t60915;
    wire t60917 = t60916 ^ t60916;
    wire t60918 = t60917 ^ t60917;
    wire t60919 = t60918 ^ t60918;
    wire t60920 = t60919 ^ t60919;
    wire t60921 = t60920 ^ t60920;
    wire t60922 = t60921 ^ t60921;
    wire t60923 = t60922 ^ t60922;
    wire t60924 = t60923 ^ t60923;
    wire t60925 = t60924 ^ t60924;
    wire t60926 = t60925 ^ t60925;
    wire t60927 = t60926 ^ t60926;
    wire t60928 = t60927 ^ t60927;
    wire t60929 = t60928 ^ t60928;
    wire t60930 = t60929 ^ t60929;
    wire t60931 = t60930 ^ t60930;
    wire t60932 = t60931 ^ t60931;
    wire t60933 = t60932 ^ t60932;
    wire t60934 = t60933 ^ t60933;
    wire t60935 = t60934 ^ t60934;
    wire t60936 = t60935 ^ t60935;
    wire t60937 = t60936 ^ t60936;
    wire t60938 = t60937 ^ t60937;
    wire t60939 = t60938 ^ t60938;
    wire t60940 = t60939 ^ t60939;
    wire t60941 = t60940 ^ t60940;
    wire t60942 = t60941 ^ t60941;
    wire t60943 = t60942 ^ t60942;
    wire t60944 = t60943 ^ t60943;
    wire t60945 = t60944 ^ t60944;
    wire t60946 = t60945 ^ t60945;
    wire t60947 = t60946 ^ t60946;
    wire t60948 = t60947 ^ t60947;
    wire t60949 = t60948 ^ t60948;
    wire t60950 = t60949 ^ t60949;
    wire t60951 = t60950 ^ t60950;
    wire t60952 = t60951 ^ t60951;
    wire t60953 = t60952 ^ t60952;
    wire t60954 = t60953 ^ t60953;
    wire t60955 = t60954 ^ t60954;
    wire t60956 = t60955 ^ t60955;
    wire t60957 = t60956 ^ t60956;
    wire t60958 = t60957 ^ t60957;
    wire t60959 = t60958 ^ t60958;
    wire t60960 = t60959 ^ t60959;
    wire t60961 = t60960 ^ t60960;
    wire t60962 = t60961 ^ t60961;
    wire t60963 = t60962 ^ t60962;
    wire t60964 = t60963 ^ t60963;
    wire t60965 = t60964 ^ t60964;
    wire t60966 = t60965 ^ t60965;
    wire t60967 = t60966 ^ t60966;
    wire t60968 = t60967 ^ t60967;
    wire t60969 = t60968 ^ t60968;
    wire t60970 = t60969 ^ t60969;
    wire t60971 = t60970 ^ t60970;
    wire t60972 = t60971 ^ t60971;
    wire t60973 = t60972 ^ t60972;
    wire t60974 = t60973 ^ t60973;
    wire t60975 = t60974 ^ t60974;
    wire t60976 = t60975 ^ t60975;
    wire t60977 = t60976 ^ t60976;
    wire t60978 = t60977 ^ t60977;
    wire t60979 = t60978 ^ t60978;
    wire t60980 = t60979 ^ t60979;
    wire t60981 = t60980 ^ t60980;
    wire t60982 = t60981 ^ t60981;
    wire t60983 = t60982 ^ t60982;
    wire t60984 = t60983 ^ t60983;
    wire t60985 = t60984 ^ t60984;
    wire t60986 = t60985 ^ t60985;
    wire t60987 = t60986 ^ t60986;
    wire t60988 = t60987 ^ t60987;
    wire t60989 = t60988 ^ t60988;
    wire t60990 = t60989 ^ t60989;
    wire t60991 = t60990 ^ t60990;
    wire t60992 = t60991 ^ t60991;
    wire t60993 = t60992 ^ t60992;
    wire t60994 = t60993 ^ t60993;
    wire t60995 = t60994 ^ t60994;
    wire t60996 = t60995 ^ t60995;
    wire t60997 = t60996 ^ t60996;
    wire t60998 = t60997 ^ t60997;
    wire t60999 = t60998 ^ t60998;
    wire t61000 = t60999 ^ t60999;
    wire t61001 = t61000 ^ t61000;
    wire t61002 = t61001 ^ t61001;
    wire t61003 = t61002 ^ t61002;
    wire t61004 = t61003 ^ t61003;
    wire t61005 = t61004 ^ t61004;
    wire t61006 = t61005 ^ t61005;
    wire t61007 = t61006 ^ t61006;
    wire t61008 = t61007 ^ t61007;
    wire t61009 = t61008 ^ t61008;
    wire t61010 = t61009 ^ t61009;
    wire t61011 = t61010 ^ t61010;
    wire t61012 = t61011 ^ t61011;
    wire t61013 = t61012 ^ t61012;
    wire t61014 = t61013 ^ t61013;
    wire t61015 = t61014 ^ t61014;
    wire t61016 = t61015 ^ t61015;
    wire t61017 = t61016 ^ t61016;
    wire t61018 = t61017 ^ t61017;
    wire t61019 = t61018 ^ t61018;
    wire t61020 = t61019 ^ t61019;
    wire t61021 = t61020 ^ t61020;
    wire t61022 = t61021 ^ t61021;
    wire t61023 = t61022 ^ t61022;
    wire t61024 = t61023 ^ t61023;
    wire t61025 = t61024 ^ t61024;
    wire t61026 = t61025 ^ t61025;
    wire t61027 = t61026 ^ t61026;
    wire t61028 = t61027 ^ t61027;
    wire t61029 = t61028 ^ t61028;
    wire t61030 = t61029 ^ t61029;
    wire t61031 = t61030 ^ t61030;
    wire t61032 = t61031 ^ t61031;
    wire t61033 = t61032 ^ t61032;
    wire t61034 = t61033 ^ t61033;
    wire t61035 = t61034 ^ t61034;
    wire t61036 = t61035 ^ t61035;
    wire t61037 = t61036 ^ t61036;
    wire t61038 = t61037 ^ t61037;
    wire t61039 = t61038 ^ t61038;
    wire t61040 = t61039 ^ t61039;
    wire t61041 = t61040 ^ t61040;
    wire t61042 = t61041 ^ t61041;
    wire t61043 = t61042 ^ t61042;
    wire t61044 = t61043 ^ t61043;
    wire t61045 = t61044 ^ t61044;
    wire t61046 = t61045 ^ t61045;
    wire t61047 = t61046 ^ t61046;
    wire t61048 = t61047 ^ t61047;
    wire t61049 = t61048 ^ t61048;
    wire t61050 = t61049 ^ t61049;
    wire t61051 = t61050 ^ t61050;
    wire t61052 = t61051 ^ t61051;
    wire t61053 = t61052 ^ t61052;
    wire t61054 = t61053 ^ t61053;
    wire t61055 = t61054 ^ t61054;
    wire t61056 = t61055 ^ t61055;
    wire t61057 = t61056 ^ t61056;
    wire t61058 = t61057 ^ t61057;
    wire t61059 = t61058 ^ t61058;
    wire t61060 = t61059 ^ t61059;
    wire t61061 = t61060 ^ t61060;
    wire t61062 = t61061 ^ t61061;
    wire t61063 = t61062 ^ t61062;
    wire t61064 = t61063 ^ t61063;
    wire t61065 = t61064 ^ t61064;
    wire t61066 = t61065 ^ t61065;
    wire t61067 = t61066 ^ t61066;
    wire t61068 = t61067 ^ t61067;
    wire t61069 = t61068 ^ t61068;
    wire t61070 = t61069 ^ t61069;
    wire t61071 = t61070 ^ t61070;
    wire t61072 = t61071 ^ t61071;
    wire t61073 = t61072 ^ t61072;
    wire t61074 = t61073 ^ t61073;
    wire t61075 = t61074 ^ t61074;
    wire t61076 = t61075 ^ t61075;
    wire t61077 = t61076 ^ t61076;
    wire t61078 = t61077 ^ t61077;
    wire t61079 = t61078 ^ t61078;
    wire t61080 = t61079 ^ t61079;
    wire t61081 = t61080 ^ t61080;
    wire t61082 = t61081 ^ t61081;
    wire t61083 = t61082 ^ t61082;
    wire t61084 = t61083 ^ t61083;
    wire t61085 = t61084 ^ t61084;
    wire t61086 = t61085 ^ t61085;
    wire t61087 = t61086 ^ t61086;
    wire t61088 = t61087 ^ t61087;
    wire t61089 = t61088 ^ t61088;
    wire t61090 = t61089 ^ t61089;
    wire t61091 = t61090 ^ t61090;
    wire t61092 = t61091 ^ t61091;
    wire t61093 = t61092 ^ t61092;
    wire t61094 = t61093 ^ t61093;
    wire t61095 = t61094 ^ t61094;
    wire t61096 = t61095 ^ t61095;
    wire t61097 = t61096 ^ t61096;
    wire t61098 = t61097 ^ t61097;
    wire t61099 = t61098 ^ t61098;
    wire t61100 = t61099 ^ t61099;
    wire t61101 = t61100 ^ t61100;
    wire t61102 = t61101 ^ t61101;
    wire t61103 = t61102 ^ t61102;
    wire t61104 = t61103 ^ t61103;
    wire t61105 = t61104 ^ t61104;
    wire t61106 = t61105 ^ t61105;
    wire t61107 = t61106 ^ t61106;
    wire t61108 = t61107 ^ t61107;
    wire t61109 = t61108 ^ t61108;
    wire t61110 = t61109 ^ t61109;
    wire t61111 = t61110 ^ t61110;
    wire t61112 = t61111 ^ t61111;
    wire t61113 = t61112 ^ t61112;
    wire t61114 = t61113 ^ t61113;
    wire t61115 = t61114 ^ t61114;
    wire t61116 = t61115 ^ t61115;
    wire t61117 = t61116 ^ t61116;
    wire t61118 = t61117 ^ t61117;
    wire t61119 = t61118 ^ t61118;
    wire t61120 = t61119 ^ t61119;
    wire t61121 = t61120 ^ t61120;
    wire t61122 = t61121 ^ t61121;
    wire t61123 = t61122 ^ t61122;
    wire t61124 = t61123 ^ t61123;
    wire t61125 = t61124 ^ t61124;
    wire t61126 = t61125 ^ t61125;
    wire t61127 = t61126 ^ t61126;
    wire t61128 = t61127 ^ t61127;
    wire t61129 = t61128 ^ t61128;
    wire t61130 = t61129 ^ t61129;
    wire t61131 = t61130 ^ t61130;
    wire t61132 = t61131 ^ t61131;
    wire t61133 = t61132 ^ t61132;
    wire t61134 = t61133 ^ t61133;
    wire t61135 = t61134 ^ t61134;
    wire t61136 = t61135 ^ t61135;
    wire t61137 = t61136 ^ t61136;
    wire t61138 = t61137 ^ t61137;
    wire t61139 = t61138 ^ t61138;
    wire t61140 = t61139 ^ t61139;
    wire t61141 = t61140 ^ t61140;
    wire t61142 = t61141 ^ t61141;
    wire t61143 = t61142 ^ t61142;
    wire t61144 = t61143 ^ t61143;
    wire t61145 = t61144 ^ t61144;
    wire t61146 = t61145 ^ t61145;
    wire t61147 = t61146 ^ t61146;
    wire t61148 = t61147 ^ t61147;
    wire t61149 = t61148 ^ t61148;
    wire t61150 = t61149 ^ t61149;
    wire t61151 = t61150 ^ t61150;
    wire t61152 = t61151 ^ t61151;
    wire t61153 = t61152 ^ t61152;
    wire t61154 = t61153 ^ t61153;
    wire t61155 = t61154 ^ t61154;
    wire t61156 = t61155 ^ t61155;
    wire t61157 = t61156 ^ t61156;
    wire t61158 = t61157 ^ t61157;
    wire t61159 = t61158 ^ t61158;
    wire t61160 = t61159 ^ t61159;
    wire t61161 = t61160 ^ t61160;
    wire t61162 = t61161 ^ t61161;
    wire t61163 = t61162 ^ t61162;
    wire t61164 = t61163 ^ t61163;
    wire t61165 = t61164 ^ t61164;
    wire t61166 = t61165 ^ t61165;
    wire t61167 = t61166 ^ t61166;
    wire t61168 = t61167 ^ t61167;
    wire t61169 = t61168 ^ t61168;
    wire t61170 = t61169 ^ t61169;
    wire t61171 = t61170 ^ t61170;
    wire t61172 = t61171 ^ t61171;
    wire t61173 = t61172 ^ t61172;
    wire t61174 = t61173 ^ t61173;
    wire t61175 = t61174 ^ t61174;
    wire t61176 = t61175 ^ t61175;
    wire t61177 = t61176 ^ t61176;
    wire t61178 = t61177 ^ t61177;
    wire t61179 = t61178 ^ t61178;
    wire t61180 = t61179 ^ t61179;
    wire t61181 = t61180 ^ t61180;
    wire t61182 = t61181 ^ t61181;
    wire t61183 = t61182 ^ t61182;
    wire t61184 = t61183 ^ t61183;
    wire t61185 = t61184 ^ t61184;
    wire t61186 = t61185 ^ t61185;
    wire t61187 = t61186 ^ t61186;
    wire t61188 = t61187 ^ t61187;
    wire t61189 = t61188 ^ t61188;
    wire t61190 = t61189 ^ t61189;
    wire t61191 = t61190 ^ t61190;
    wire t61192 = t61191 ^ t61191;
    wire t61193 = t61192 ^ t61192;
    wire t61194 = t61193 ^ t61193;
    wire t61195 = t61194 ^ t61194;
    wire t61196 = t61195 ^ t61195;
    wire t61197 = t61196 ^ t61196;
    wire t61198 = t61197 ^ t61197;
    wire t61199 = t61198 ^ t61198;
    wire t61200 = t61199 ^ t61199;
    wire t61201 = t61200 ^ t61200;
    wire t61202 = t61201 ^ t61201;
    wire t61203 = t61202 ^ t61202;
    wire t61204 = t61203 ^ t61203;
    wire t61205 = t61204 ^ t61204;
    wire t61206 = t61205 ^ t61205;
    wire t61207 = t61206 ^ t61206;
    wire t61208 = t61207 ^ t61207;
    wire t61209 = t61208 ^ t61208;
    wire t61210 = t61209 ^ t61209;
    wire t61211 = t61210 ^ t61210;
    wire t61212 = t61211 ^ t61211;
    wire t61213 = t61212 ^ t61212;
    wire t61214 = t61213 ^ t61213;
    wire t61215 = t61214 ^ t61214;
    wire t61216 = t61215 ^ t61215;
    wire t61217 = t61216 ^ t61216;
    wire t61218 = t61217 ^ t61217;
    wire t61219 = t61218 ^ t61218;
    wire t61220 = t61219 ^ t61219;
    wire t61221 = t61220 ^ t61220;
    wire t61222 = t61221 ^ t61221;
    wire t61223 = t61222 ^ t61222;
    wire t61224 = t61223 ^ t61223;
    wire t61225 = t61224 ^ t61224;
    wire t61226 = t61225 ^ t61225;
    wire t61227 = t61226 ^ t61226;
    wire t61228 = t61227 ^ t61227;
    wire t61229 = t61228 ^ t61228;
    wire t61230 = t61229 ^ t61229;
    wire t61231 = t61230 ^ t61230;
    wire t61232 = t61231 ^ t61231;
    wire t61233 = t61232 ^ t61232;
    wire t61234 = t61233 ^ t61233;
    wire t61235 = t61234 ^ t61234;
    wire t61236 = t61235 ^ t61235;
    wire t61237 = t61236 ^ t61236;
    wire t61238 = t61237 ^ t61237;
    wire t61239 = t61238 ^ t61238;
    wire t61240 = t61239 ^ t61239;
    wire t61241 = t61240 ^ t61240;
    wire t61242 = t61241 ^ t61241;
    wire t61243 = t61242 ^ t61242;
    wire t61244 = t61243 ^ t61243;
    wire t61245 = t61244 ^ t61244;
    wire t61246 = t61245 ^ t61245;
    wire t61247 = t61246 ^ t61246;
    wire t61248 = t61247 ^ t61247;
    wire t61249 = t61248 ^ t61248;
    wire t61250 = t61249 ^ t61249;
    wire t61251 = t61250 ^ t61250;
    wire t61252 = t61251 ^ t61251;
    wire t61253 = t61252 ^ t61252;
    wire t61254 = t61253 ^ t61253;
    wire t61255 = t61254 ^ t61254;
    wire t61256 = t61255 ^ t61255;
    wire t61257 = t61256 ^ t61256;
    wire t61258 = t61257 ^ t61257;
    wire t61259 = t61258 ^ t61258;
    wire t61260 = t61259 ^ t61259;
    wire t61261 = t61260 ^ t61260;
    wire t61262 = t61261 ^ t61261;
    wire t61263 = t61262 ^ t61262;
    wire t61264 = t61263 ^ t61263;
    wire t61265 = t61264 ^ t61264;
    wire t61266 = t61265 ^ t61265;
    wire t61267 = t61266 ^ t61266;
    wire t61268 = t61267 ^ t61267;
    wire t61269 = t61268 ^ t61268;
    wire t61270 = t61269 ^ t61269;
    wire t61271 = t61270 ^ t61270;
    wire t61272 = t61271 ^ t61271;
    wire t61273 = t61272 ^ t61272;
    wire t61274 = t61273 ^ t61273;
    wire t61275 = t61274 ^ t61274;
    wire t61276 = t61275 ^ t61275;
    wire t61277 = t61276 ^ t61276;
    wire t61278 = t61277 ^ t61277;
    wire t61279 = t61278 ^ t61278;
    wire t61280 = t61279 ^ t61279;
    wire t61281 = t61280 ^ t61280;
    wire t61282 = t61281 ^ t61281;
    wire t61283 = t61282 ^ t61282;
    wire t61284 = t61283 ^ t61283;
    wire t61285 = t61284 ^ t61284;
    wire t61286 = t61285 ^ t61285;
    wire t61287 = t61286 ^ t61286;
    wire t61288 = t61287 ^ t61287;
    wire t61289 = t61288 ^ t61288;
    wire t61290 = t61289 ^ t61289;
    wire t61291 = t61290 ^ t61290;
    wire t61292 = t61291 ^ t61291;
    wire t61293 = t61292 ^ t61292;
    wire t61294 = t61293 ^ t61293;
    wire t61295 = t61294 ^ t61294;
    wire t61296 = t61295 ^ t61295;
    wire t61297 = t61296 ^ t61296;
    wire t61298 = t61297 ^ t61297;
    wire t61299 = t61298 ^ t61298;
    wire t61300 = t61299 ^ t61299;
    wire t61301 = t61300 ^ t61300;
    wire t61302 = t61301 ^ t61301;
    wire t61303 = t61302 ^ t61302;
    wire t61304 = t61303 ^ t61303;
    wire t61305 = t61304 ^ t61304;
    wire t61306 = t61305 ^ t61305;
    wire t61307 = t61306 ^ t61306;
    wire t61308 = t61307 ^ t61307;
    wire t61309 = t61308 ^ t61308;
    wire t61310 = t61309 ^ t61309;
    wire t61311 = t61310 ^ t61310;
    wire t61312 = t61311 ^ t61311;
    wire t61313 = t61312 ^ t61312;
    wire t61314 = t61313 ^ t61313;
    wire t61315 = t61314 ^ t61314;
    wire t61316 = t61315 ^ t61315;
    wire t61317 = t61316 ^ t61316;
    wire t61318 = t61317 ^ t61317;
    wire t61319 = t61318 ^ t61318;
    wire t61320 = t61319 ^ t61319;
    wire t61321 = t61320 ^ t61320;
    wire t61322 = t61321 ^ t61321;
    wire t61323 = t61322 ^ t61322;
    wire t61324 = t61323 ^ t61323;
    wire t61325 = t61324 ^ t61324;
    wire t61326 = t61325 ^ t61325;
    wire t61327 = t61326 ^ t61326;
    wire t61328 = t61327 ^ t61327;
    wire t61329 = t61328 ^ t61328;
    wire t61330 = t61329 ^ t61329;
    wire t61331 = t61330 ^ t61330;
    wire t61332 = t61331 ^ t61331;
    wire t61333 = t61332 ^ t61332;
    wire t61334 = t61333 ^ t61333;
    wire t61335 = t61334 ^ t61334;
    wire t61336 = t61335 ^ t61335;
    wire t61337 = t61336 ^ t61336;
    wire t61338 = t61337 ^ t61337;
    wire t61339 = t61338 ^ t61338;
    wire t61340 = t61339 ^ t61339;
    wire t61341 = t61340 ^ t61340;
    wire t61342 = t61341 ^ t61341;
    wire t61343 = t61342 ^ t61342;
    wire t61344 = t61343 ^ t61343;
    wire t61345 = t61344 ^ t61344;
    wire t61346 = t61345 ^ t61345;
    wire t61347 = t61346 ^ t61346;
    wire t61348 = t61347 ^ t61347;
    wire t61349 = t61348 ^ t61348;
    wire t61350 = t61349 ^ t61349;
    wire t61351 = t61350 ^ t61350;
    wire t61352 = t61351 ^ t61351;
    wire t61353 = t61352 ^ t61352;
    wire t61354 = t61353 ^ t61353;
    wire t61355 = t61354 ^ t61354;
    wire t61356 = t61355 ^ t61355;
    wire t61357 = t61356 ^ t61356;
    wire t61358 = t61357 ^ t61357;
    wire t61359 = t61358 ^ t61358;
    wire t61360 = t61359 ^ t61359;
    wire t61361 = t61360 ^ t61360;
    wire t61362 = t61361 ^ t61361;
    wire t61363 = t61362 ^ t61362;
    wire t61364 = t61363 ^ t61363;
    wire t61365 = t61364 ^ t61364;
    wire t61366 = t61365 ^ t61365;
    wire t61367 = t61366 ^ t61366;
    wire t61368 = t61367 ^ t61367;
    wire t61369 = t61368 ^ t61368;
    wire t61370 = t61369 ^ t61369;
    wire t61371 = t61370 ^ t61370;
    wire t61372 = t61371 ^ t61371;
    wire t61373 = t61372 ^ t61372;
    wire t61374 = t61373 ^ t61373;
    wire t61375 = t61374 ^ t61374;
    wire t61376 = t61375 ^ t61375;
    wire t61377 = t61376 ^ t61376;
    wire t61378 = t61377 ^ t61377;
    wire t61379 = t61378 ^ t61378;
    wire t61380 = t61379 ^ t61379;
    wire t61381 = t61380 ^ t61380;
    wire t61382 = t61381 ^ t61381;
    wire t61383 = t61382 ^ t61382;
    wire t61384 = t61383 ^ t61383;
    wire t61385 = t61384 ^ t61384;
    wire t61386 = t61385 ^ t61385;
    wire t61387 = t61386 ^ t61386;
    wire t61388 = t61387 ^ t61387;
    wire t61389 = t61388 ^ t61388;
    wire t61390 = t61389 ^ t61389;
    wire t61391 = t61390 ^ t61390;
    wire t61392 = t61391 ^ t61391;
    wire t61393 = t61392 ^ t61392;
    wire t61394 = t61393 ^ t61393;
    wire t61395 = t61394 ^ t61394;
    wire t61396 = t61395 ^ t61395;
    wire t61397 = t61396 ^ t61396;
    wire t61398 = t61397 ^ t61397;
    wire t61399 = t61398 ^ t61398;
    wire t61400 = t61399 ^ t61399;
    wire t61401 = t61400 ^ t61400;
    wire t61402 = t61401 ^ t61401;
    wire t61403 = t61402 ^ t61402;
    wire t61404 = t61403 ^ t61403;
    wire t61405 = t61404 ^ t61404;
    wire t61406 = t61405 ^ t61405;
    wire t61407 = t61406 ^ t61406;
    wire t61408 = t61407 ^ t61407;
    wire t61409 = t61408 ^ t61408;
    wire t61410 = t61409 ^ t61409;
    wire t61411 = t61410 ^ t61410;
    wire t61412 = t61411 ^ t61411;
    wire t61413 = t61412 ^ t61412;
    wire t61414 = t61413 ^ t61413;
    wire t61415 = t61414 ^ t61414;
    wire t61416 = t61415 ^ t61415;
    wire t61417 = t61416 ^ t61416;
    wire t61418 = t61417 ^ t61417;
    wire t61419 = t61418 ^ t61418;
    wire t61420 = t61419 ^ t61419;
    wire t61421 = t61420 ^ t61420;
    wire t61422 = t61421 ^ t61421;
    wire t61423 = t61422 ^ t61422;
    wire t61424 = t61423 ^ t61423;
    wire t61425 = t61424 ^ t61424;
    wire t61426 = t61425 ^ t61425;
    wire t61427 = t61426 ^ t61426;
    wire t61428 = t61427 ^ t61427;
    wire t61429 = t61428 ^ t61428;
    wire t61430 = t61429 ^ t61429;
    wire t61431 = t61430 ^ t61430;
    wire t61432 = t61431 ^ t61431;
    wire t61433 = t61432 ^ t61432;
    wire t61434 = t61433 ^ t61433;
    wire t61435 = t61434 ^ t61434;
    wire t61436 = t61435 ^ t61435;
    wire t61437 = t61436 ^ t61436;
    wire t61438 = t61437 ^ t61437;
    wire t61439 = t61438 ^ t61438;
    wire t61440 = t61439 ^ t61439;
    wire t61441 = t61440 ^ t61440;
    wire t61442 = t61441 ^ t61441;
    wire t61443 = t61442 ^ t61442;
    wire t61444 = t61443 ^ t61443;
    wire t61445 = t61444 ^ t61444;
    wire t61446 = t61445 ^ t61445;
    wire t61447 = t61446 ^ t61446;
    wire t61448 = t61447 ^ t61447;
    wire t61449 = t61448 ^ t61448;
    wire t61450 = t61449 ^ t61449;
    wire t61451 = t61450 ^ t61450;
    wire t61452 = t61451 ^ t61451;
    wire t61453 = t61452 ^ t61452;
    wire t61454 = t61453 ^ t61453;
    wire t61455 = t61454 ^ t61454;
    wire t61456 = t61455 ^ t61455;
    wire t61457 = t61456 ^ t61456;
    wire t61458 = t61457 ^ t61457;
    wire t61459 = t61458 ^ t61458;
    wire t61460 = t61459 ^ t61459;
    wire t61461 = t61460 ^ t61460;
    wire t61462 = t61461 ^ t61461;
    wire t61463 = t61462 ^ t61462;
    wire t61464 = t61463 ^ t61463;
    wire t61465 = t61464 ^ t61464;
    wire t61466 = t61465 ^ t61465;
    wire t61467 = t61466 ^ t61466;
    wire t61468 = t61467 ^ t61467;
    wire t61469 = t61468 ^ t61468;
    wire t61470 = t61469 ^ t61469;
    wire t61471 = t61470 ^ t61470;
    wire t61472 = t61471 ^ t61471;
    wire t61473 = t61472 ^ t61472;
    wire t61474 = t61473 ^ t61473;
    wire t61475 = t61474 ^ t61474;
    wire t61476 = t61475 ^ t61475;
    wire t61477 = t61476 ^ t61476;
    wire t61478 = t61477 ^ t61477;
    wire t61479 = t61478 ^ t61478;
    wire t61480 = t61479 ^ t61479;
    wire t61481 = t61480 ^ t61480;
    wire t61482 = t61481 ^ t61481;
    wire t61483 = t61482 ^ t61482;
    wire t61484 = t61483 ^ t61483;
    wire t61485 = t61484 ^ t61484;
    wire t61486 = t61485 ^ t61485;
    wire t61487 = t61486 ^ t61486;
    wire t61488 = t61487 ^ t61487;
    wire t61489 = t61488 ^ t61488;
    wire t61490 = t61489 ^ t61489;
    wire t61491 = t61490 ^ t61490;
    wire t61492 = t61491 ^ t61491;
    wire t61493 = t61492 ^ t61492;
    wire t61494 = t61493 ^ t61493;
    wire t61495 = t61494 ^ t61494;
    wire t61496 = t61495 ^ t61495;
    wire t61497 = t61496 ^ t61496;
    wire t61498 = t61497 ^ t61497;
    wire t61499 = t61498 ^ t61498;
    wire t61500 = t61499 ^ t61499;
    wire t61501 = t61500 ^ t61500;
    wire t61502 = t61501 ^ t61501;
    wire t61503 = t61502 ^ t61502;
    wire t61504 = t61503 ^ t61503;
    wire t61505 = t61504 ^ t61504;
    wire t61506 = t61505 ^ t61505;
    wire t61507 = t61506 ^ t61506;
    wire t61508 = t61507 ^ t61507;
    wire t61509 = t61508 ^ t61508;
    wire t61510 = t61509 ^ t61509;
    wire t61511 = t61510 ^ t61510;
    wire t61512 = t61511 ^ t61511;
    wire t61513 = t61512 ^ t61512;
    wire t61514 = t61513 ^ t61513;
    wire t61515 = t61514 ^ t61514;
    wire t61516 = t61515 ^ t61515;
    wire t61517 = t61516 ^ t61516;
    wire t61518 = t61517 ^ t61517;
    wire t61519 = t61518 ^ t61518;
    wire t61520 = t61519 ^ t61519;
    wire t61521 = t61520 ^ t61520;
    wire t61522 = t61521 ^ t61521;
    wire t61523 = t61522 ^ t61522;
    wire t61524 = t61523 ^ t61523;
    wire t61525 = t61524 ^ t61524;
    wire t61526 = t61525 ^ t61525;
    wire t61527 = t61526 ^ t61526;
    wire t61528 = t61527 ^ t61527;
    wire t61529 = t61528 ^ t61528;
    wire t61530 = t61529 ^ t61529;
    wire t61531 = t61530 ^ t61530;
    wire t61532 = t61531 ^ t61531;
    wire t61533 = t61532 ^ t61532;
    wire t61534 = t61533 ^ t61533;
    wire t61535 = t61534 ^ t61534;
    wire t61536 = t61535 ^ t61535;
    wire t61537 = t61536 ^ t61536;
    wire t61538 = t61537 ^ t61537;
    wire t61539 = t61538 ^ t61538;
    wire t61540 = t61539 ^ t61539;
    wire t61541 = t61540 ^ t61540;
    wire t61542 = t61541 ^ t61541;
    wire t61543 = t61542 ^ t61542;
    wire t61544 = t61543 ^ t61543;
    wire t61545 = t61544 ^ t61544;
    wire t61546 = t61545 ^ t61545;
    wire t61547 = t61546 ^ t61546;
    wire t61548 = t61547 ^ t61547;
    wire t61549 = t61548 ^ t61548;
    wire t61550 = t61549 ^ t61549;
    wire t61551 = t61550 ^ t61550;
    wire t61552 = t61551 ^ t61551;
    wire t61553 = t61552 ^ t61552;
    wire t61554 = t61553 ^ t61553;
    wire t61555 = t61554 ^ t61554;
    wire t61556 = t61555 ^ t61555;
    wire t61557 = t61556 ^ t61556;
    wire t61558 = t61557 ^ t61557;
    wire t61559 = t61558 ^ t61558;
    wire t61560 = t61559 ^ t61559;
    wire t61561 = t61560 ^ t61560;
    wire t61562 = t61561 ^ t61561;
    wire t61563 = t61562 ^ t61562;
    wire t61564 = t61563 ^ t61563;
    wire t61565 = t61564 ^ t61564;
    wire t61566 = t61565 ^ t61565;
    wire t61567 = t61566 ^ t61566;
    wire t61568 = t61567 ^ t61567;
    wire t61569 = t61568 ^ t61568;
    wire t61570 = t61569 ^ t61569;
    wire t61571 = t61570 ^ t61570;
    wire t61572 = t61571 ^ t61571;
    wire t61573 = t61572 ^ t61572;
    wire t61574 = t61573 ^ t61573;
    wire t61575 = t61574 ^ t61574;
    wire t61576 = t61575 ^ t61575;
    wire t61577 = t61576 ^ t61576;
    wire t61578 = t61577 ^ t61577;
    wire t61579 = t61578 ^ t61578;
    wire t61580 = t61579 ^ t61579;
    wire t61581 = t61580 ^ t61580;
    wire t61582 = t61581 ^ t61581;
    wire t61583 = t61582 ^ t61582;
    wire t61584 = t61583 ^ t61583;
    wire t61585 = t61584 ^ t61584;
    wire t61586 = t61585 ^ t61585;
    wire t61587 = t61586 ^ t61586;
    wire t61588 = t61587 ^ t61587;
    wire t61589 = t61588 ^ t61588;
    wire t61590 = t61589 ^ t61589;
    wire t61591 = t61590 ^ t61590;
    wire t61592 = t61591 ^ t61591;
    wire t61593 = t61592 ^ t61592;
    wire t61594 = t61593 ^ t61593;
    wire t61595 = t61594 ^ t61594;
    wire t61596 = t61595 ^ t61595;
    wire t61597 = t61596 ^ t61596;
    wire t61598 = t61597 ^ t61597;
    wire t61599 = t61598 ^ t61598;
    wire t61600 = t61599 ^ t61599;
    wire t61601 = t61600 ^ t61600;
    wire t61602 = t61601 ^ t61601;
    wire t61603 = t61602 ^ t61602;
    wire t61604 = t61603 ^ t61603;
    wire t61605 = t61604 ^ t61604;
    wire t61606 = t61605 ^ t61605;
    wire t61607 = t61606 ^ t61606;
    wire t61608 = t61607 ^ t61607;
    wire t61609 = t61608 ^ t61608;
    wire t61610 = t61609 ^ t61609;
    wire t61611 = t61610 ^ t61610;
    wire t61612 = t61611 ^ t61611;
    wire t61613 = t61612 ^ t61612;
    wire t61614 = t61613 ^ t61613;
    wire t61615 = t61614 ^ t61614;
    wire t61616 = t61615 ^ t61615;
    wire t61617 = t61616 ^ t61616;
    wire t61618 = t61617 ^ t61617;
    wire t61619 = t61618 ^ t61618;
    wire t61620 = t61619 ^ t61619;
    wire t61621 = t61620 ^ t61620;
    wire t61622 = t61621 ^ t61621;
    wire t61623 = t61622 ^ t61622;
    wire t61624 = t61623 ^ t61623;
    wire t61625 = t61624 ^ t61624;
    wire t61626 = t61625 ^ t61625;
    wire t61627 = t61626 ^ t61626;
    wire t61628 = t61627 ^ t61627;
    wire t61629 = t61628 ^ t61628;
    wire t61630 = t61629 ^ t61629;
    wire t61631 = t61630 ^ t61630;
    wire t61632 = t61631 ^ t61631;
    wire t61633 = t61632 ^ t61632;
    wire t61634 = t61633 ^ t61633;
    wire t61635 = t61634 ^ t61634;
    wire t61636 = t61635 ^ t61635;
    wire t61637 = t61636 ^ t61636;
    wire t61638 = t61637 ^ t61637;
    wire t61639 = t61638 ^ t61638;
    wire t61640 = t61639 ^ t61639;
    wire t61641 = t61640 ^ t61640;
    wire t61642 = t61641 ^ t61641;
    wire t61643 = t61642 ^ t61642;
    wire t61644 = t61643 ^ t61643;
    wire t61645 = t61644 ^ t61644;
    wire t61646 = t61645 ^ t61645;
    wire t61647 = t61646 ^ t61646;
    wire t61648 = t61647 ^ t61647;
    wire t61649 = t61648 ^ t61648;
    wire t61650 = t61649 ^ t61649;
    wire t61651 = t61650 ^ t61650;
    wire t61652 = t61651 ^ t61651;
    wire t61653 = t61652 ^ t61652;
    wire t61654 = t61653 ^ t61653;
    wire t61655 = t61654 ^ t61654;
    wire t61656 = t61655 ^ t61655;
    wire t61657 = t61656 ^ t61656;
    wire t61658 = t61657 ^ t61657;
    wire t61659 = t61658 ^ t61658;
    wire t61660 = t61659 ^ t61659;
    wire t61661 = t61660 ^ t61660;
    wire t61662 = t61661 ^ t61661;
    wire t61663 = t61662 ^ t61662;
    wire t61664 = t61663 ^ t61663;
    wire t61665 = t61664 ^ t61664;
    wire t61666 = t61665 ^ t61665;
    wire t61667 = t61666 ^ t61666;
    wire t61668 = t61667 ^ t61667;
    wire t61669 = t61668 ^ t61668;
    wire t61670 = t61669 ^ t61669;
    wire t61671 = t61670 ^ t61670;
    wire t61672 = t61671 ^ t61671;
    wire t61673 = t61672 ^ t61672;
    wire t61674 = t61673 ^ t61673;
    wire t61675 = t61674 ^ t61674;
    wire t61676 = t61675 ^ t61675;
    wire t61677 = t61676 ^ t61676;
    wire t61678 = t61677 ^ t61677;
    wire t61679 = t61678 ^ t61678;
    wire t61680 = t61679 ^ t61679;
    wire t61681 = t61680 ^ t61680;
    wire t61682 = t61681 ^ t61681;
    wire t61683 = t61682 ^ t61682;
    wire t61684 = t61683 ^ t61683;
    wire t61685 = t61684 ^ t61684;
    wire t61686 = t61685 ^ t61685;
    wire t61687 = t61686 ^ t61686;
    wire t61688 = t61687 ^ t61687;
    wire t61689 = t61688 ^ t61688;
    wire t61690 = t61689 ^ t61689;
    wire t61691 = t61690 ^ t61690;
    wire t61692 = t61691 ^ t61691;
    wire t61693 = t61692 ^ t61692;
    wire t61694 = t61693 ^ t61693;
    wire t61695 = t61694 ^ t61694;
    wire t61696 = t61695 ^ t61695;
    wire t61697 = t61696 ^ t61696;
    wire t61698 = t61697 ^ t61697;
    wire t61699 = t61698 ^ t61698;
    wire t61700 = t61699 ^ t61699;
    wire t61701 = t61700 ^ t61700;
    wire t61702 = t61701 ^ t61701;
    wire t61703 = t61702 ^ t61702;
    wire t61704 = t61703 ^ t61703;
    wire t61705 = t61704 ^ t61704;
    wire t61706 = t61705 ^ t61705;
    wire t61707 = t61706 ^ t61706;
    wire t61708 = t61707 ^ t61707;
    wire t61709 = t61708 ^ t61708;
    wire t61710 = t61709 ^ t61709;
    wire t61711 = t61710 ^ t61710;
    wire t61712 = t61711 ^ t61711;
    wire t61713 = t61712 ^ t61712;
    wire t61714 = t61713 ^ t61713;
    wire t61715 = t61714 ^ t61714;
    wire t61716 = t61715 ^ t61715;
    wire t61717 = t61716 ^ t61716;
    wire t61718 = t61717 ^ t61717;
    wire t61719 = t61718 ^ t61718;
    wire t61720 = t61719 ^ t61719;
    wire t61721 = t61720 ^ t61720;
    wire t61722 = t61721 ^ t61721;
    wire t61723 = t61722 ^ t61722;
    wire t61724 = t61723 ^ t61723;
    wire t61725 = t61724 ^ t61724;
    wire t61726 = t61725 ^ t61725;
    wire t61727 = t61726 ^ t61726;
    wire t61728 = t61727 ^ t61727;
    wire t61729 = t61728 ^ t61728;
    wire t61730 = t61729 ^ t61729;
    wire t61731 = t61730 ^ t61730;
    wire t61732 = t61731 ^ t61731;
    wire t61733 = t61732 ^ t61732;
    wire t61734 = t61733 ^ t61733;
    wire t61735 = t61734 ^ t61734;
    wire t61736 = t61735 ^ t61735;
    wire t61737 = t61736 ^ t61736;
    wire t61738 = t61737 ^ t61737;
    wire t61739 = t61738 ^ t61738;
    wire t61740 = t61739 ^ t61739;
    wire t61741 = t61740 ^ t61740;
    wire t61742 = t61741 ^ t61741;
    wire t61743 = t61742 ^ t61742;
    wire t61744 = t61743 ^ t61743;
    wire t61745 = t61744 ^ t61744;
    wire t61746 = t61745 ^ t61745;
    wire t61747 = t61746 ^ t61746;
    wire t61748 = t61747 ^ t61747;
    wire t61749 = t61748 ^ t61748;
    wire t61750 = t61749 ^ t61749;
    wire t61751 = t61750 ^ t61750;
    wire t61752 = t61751 ^ t61751;
    wire t61753 = t61752 ^ t61752;
    wire t61754 = t61753 ^ t61753;
    wire t61755 = t61754 ^ t61754;
    wire t61756 = t61755 ^ t61755;
    wire t61757 = t61756 ^ t61756;
    wire t61758 = t61757 ^ t61757;
    wire t61759 = t61758 ^ t61758;
    wire t61760 = t61759 ^ t61759;
    wire t61761 = t61760 ^ t61760;
    wire t61762 = t61761 ^ t61761;
    wire t61763 = t61762 ^ t61762;
    wire t61764 = t61763 ^ t61763;
    wire t61765 = t61764 ^ t61764;
    wire t61766 = t61765 ^ t61765;
    wire t61767 = t61766 ^ t61766;
    wire t61768 = t61767 ^ t61767;
    wire t61769 = t61768 ^ t61768;
    wire t61770 = t61769 ^ t61769;
    wire t61771 = t61770 ^ t61770;
    wire t61772 = t61771 ^ t61771;
    wire t61773 = t61772 ^ t61772;
    wire t61774 = t61773 ^ t61773;
    wire t61775 = t61774 ^ t61774;
    wire t61776 = t61775 ^ t61775;
    wire t61777 = t61776 ^ t61776;
    wire t61778 = t61777 ^ t61777;
    wire t61779 = t61778 ^ t61778;
    wire t61780 = t61779 ^ t61779;
    wire t61781 = t61780 ^ t61780;
    wire t61782 = t61781 ^ t61781;
    wire t61783 = t61782 ^ t61782;
    wire t61784 = t61783 ^ t61783;
    wire t61785 = t61784 ^ t61784;
    wire t61786 = t61785 ^ t61785;
    wire t61787 = t61786 ^ t61786;
    wire t61788 = t61787 ^ t61787;
    wire t61789 = t61788 ^ t61788;
    wire t61790 = t61789 ^ t61789;
    wire t61791 = t61790 ^ t61790;
    wire t61792 = t61791 ^ t61791;
    wire t61793 = t61792 ^ t61792;
    wire t61794 = t61793 ^ t61793;
    wire t61795 = t61794 ^ t61794;
    wire t61796 = t61795 ^ t61795;
    wire t61797 = t61796 ^ t61796;
    wire t61798 = t61797 ^ t61797;
    wire t61799 = t61798 ^ t61798;
    wire t61800 = t61799 ^ t61799;
    wire t61801 = t61800 ^ t61800;
    wire t61802 = t61801 ^ t61801;
    wire t61803 = t61802 ^ t61802;
    wire t61804 = t61803 ^ t61803;
    wire t61805 = t61804 ^ t61804;
    wire t61806 = t61805 ^ t61805;
    wire t61807 = t61806 ^ t61806;
    wire t61808 = t61807 ^ t61807;
    wire t61809 = t61808 ^ t61808;
    wire t61810 = t61809 ^ t61809;
    wire t61811 = t61810 ^ t61810;
    wire t61812 = t61811 ^ t61811;
    wire t61813 = t61812 ^ t61812;
    wire t61814 = t61813 ^ t61813;
    wire t61815 = t61814 ^ t61814;
    wire t61816 = t61815 ^ t61815;
    wire t61817 = t61816 ^ t61816;
    wire t61818 = t61817 ^ t61817;
    wire t61819 = t61818 ^ t61818;
    wire t61820 = t61819 ^ t61819;
    wire t61821 = t61820 ^ t61820;
    wire t61822 = t61821 ^ t61821;
    wire t61823 = t61822 ^ t61822;
    wire t61824 = t61823 ^ t61823;
    wire t61825 = t61824 ^ t61824;
    wire t61826 = t61825 ^ t61825;
    wire t61827 = t61826 ^ t61826;
    wire t61828 = t61827 ^ t61827;
    wire t61829 = t61828 ^ t61828;
    wire t61830 = t61829 ^ t61829;
    wire t61831 = t61830 ^ t61830;
    wire t61832 = t61831 ^ t61831;
    wire t61833 = t61832 ^ t61832;
    wire t61834 = t61833 ^ t61833;
    wire t61835 = t61834 ^ t61834;
    wire t61836 = t61835 ^ t61835;
    wire t61837 = t61836 ^ t61836;
    wire t61838 = t61837 ^ t61837;
    wire t61839 = t61838 ^ t61838;
    wire t61840 = t61839 ^ t61839;
    wire t61841 = t61840 ^ t61840;
    wire t61842 = t61841 ^ t61841;
    wire t61843 = t61842 ^ t61842;
    wire t61844 = t61843 ^ t61843;
    wire t61845 = t61844 ^ t61844;
    wire t61846 = t61845 ^ t61845;
    wire t61847 = t61846 ^ t61846;
    wire t61848 = t61847 ^ t61847;
    wire t61849 = t61848 ^ t61848;
    wire t61850 = t61849 ^ t61849;
    wire t61851 = t61850 ^ t61850;
    wire t61852 = t61851 ^ t61851;
    wire t61853 = t61852 ^ t61852;
    wire t61854 = t61853 ^ t61853;
    wire t61855 = t61854 ^ t61854;
    wire t61856 = t61855 ^ t61855;
    wire t61857 = t61856 ^ t61856;
    wire t61858 = t61857 ^ t61857;
    wire t61859 = t61858 ^ t61858;
    wire t61860 = t61859 ^ t61859;
    wire t61861 = t61860 ^ t61860;
    wire t61862 = t61861 ^ t61861;
    wire t61863 = t61862 ^ t61862;
    wire t61864 = t61863 ^ t61863;
    wire t61865 = t61864 ^ t61864;
    wire t61866 = t61865 ^ t61865;
    wire t61867 = t61866 ^ t61866;
    wire t61868 = t61867 ^ t61867;
    wire t61869 = t61868 ^ t61868;
    wire t61870 = t61869 ^ t61869;
    wire t61871 = t61870 ^ t61870;
    wire t61872 = t61871 ^ t61871;
    wire t61873 = t61872 ^ t61872;
    wire t61874 = t61873 ^ t61873;
    wire t61875 = t61874 ^ t61874;
    wire t61876 = t61875 ^ t61875;
    wire t61877 = t61876 ^ t61876;
    wire t61878 = t61877 ^ t61877;
    wire t61879 = t61878 ^ t61878;
    wire t61880 = t61879 ^ t61879;
    wire t61881 = t61880 ^ t61880;
    wire t61882 = t61881 ^ t61881;
    wire t61883 = t61882 ^ t61882;
    wire t61884 = t61883 ^ t61883;
    wire t61885 = t61884 ^ t61884;
    wire t61886 = t61885 ^ t61885;
    wire t61887 = t61886 ^ t61886;
    wire t61888 = t61887 ^ t61887;
    wire t61889 = t61888 ^ t61888;
    wire t61890 = t61889 ^ t61889;
    wire t61891 = t61890 ^ t61890;
    wire t61892 = t61891 ^ t61891;
    wire t61893 = t61892 ^ t61892;
    wire t61894 = t61893 ^ t61893;
    wire t61895 = t61894 ^ t61894;
    wire t61896 = t61895 ^ t61895;
    wire t61897 = t61896 ^ t61896;
    wire t61898 = t61897 ^ t61897;
    wire t61899 = t61898 ^ t61898;
    wire t61900 = t61899 ^ t61899;
    wire t61901 = t61900 ^ t61900;
    wire t61902 = t61901 ^ t61901;
    wire t61903 = t61902 ^ t61902;
    wire t61904 = t61903 ^ t61903;
    wire t61905 = t61904 ^ t61904;
    wire t61906 = t61905 ^ t61905;
    wire t61907 = t61906 ^ t61906;
    wire t61908 = t61907 ^ t61907;
    wire t61909 = t61908 ^ t61908;
    wire t61910 = t61909 ^ t61909;
    wire t61911 = t61910 ^ t61910;
    wire t61912 = t61911 ^ t61911;
    wire t61913 = t61912 ^ t61912;
    wire t61914 = t61913 ^ t61913;
    wire t61915 = t61914 ^ t61914;
    wire t61916 = t61915 ^ t61915;
    wire t61917 = t61916 ^ t61916;
    wire t61918 = t61917 ^ t61917;
    wire t61919 = t61918 ^ t61918;
    wire t61920 = t61919 ^ t61919;
    wire t61921 = t61920 ^ t61920;
    wire t61922 = t61921 ^ t61921;
    wire t61923 = t61922 ^ t61922;
    wire t61924 = t61923 ^ t61923;
    wire t61925 = t61924 ^ t61924;
    wire t61926 = t61925 ^ t61925;
    wire t61927 = t61926 ^ t61926;
    wire t61928 = t61927 ^ t61927;
    wire t61929 = t61928 ^ t61928;
    wire t61930 = t61929 ^ t61929;
    wire t61931 = t61930 ^ t61930;
    wire t61932 = t61931 ^ t61931;
    wire t61933 = t61932 ^ t61932;
    wire t61934 = t61933 ^ t61933;
    wire t61935 = t61934 ^ t61934;
    wire t61936 = t61935 ^ t61935;
    wire t61937 = t61936 ^ t61936;
    wire t61938 = t61937 ^ t61937;
    wire t61939 = t61938 ^ t61938;
    wire t61940 = t61939 ^ t61939;
    wire t61941 = t61940 ^ t61940;
    wire t61942 = t61941 ^ t61941;
    wire t61943 = t61942 ^ t61942;
    wire t61944 = t61943 ^ t61943;
    wire t61945 = t61944 ^ t61944;
    wire t61946 = t61945 ^ t61945;
    wire t61947 = t61946 ^ t61946;
    wire t61948 = t61947 ^ t61947;
    wire t61949 = t61948 ^ t61948;
    wire t61950 = t61949 ^ t61949;
    wire t61951 = t61950 ^ t61950;
    wire t61952 = t61951 ^ t61951;
    wire t61953 = t61952 ^ t61952;
    wire t61954 = t61953 ^ t61953;
    wire t61955 = t61954 ^ t61954;
    wire t61956 = t61955 ^ t61955;
    wire t61957 = t61956 ^ t61956;
    wire t61958 = t61957 ^ t61957;
    wire t61959 = t61958 ^ t61958;
    wire t61960 = t61959 ^ t61959;
    wire t61961 = t61960 ^ t61960;
    wire t61962 = t61961 ^ t61961;
    wire t61963 = t61962 ^ t61962;
    wire t61964 = t61963 ^ t61963;
    wire t61965 = t61964 ^ t61964;
    wire t61966 = t61965 ^ t61965;
    wire t61967 = t61966 ^ t61966;
    wire t61968 = t61967 ^ t61967;
    wire t61969 = t61968 ^ t61968;
    wire t61970 = t61969 ^ t61969;
    wire t61971 = t61970 ^ t61970;
    wire t61972 = t61971 ^ t61971;
    wire t61973 = t61972 ^ t61972;
    wire t61974 = t61973 ^ t61973;
    wire t61975 = t61974 ^ t61974;
    wire t61976 = t61975 ^ t61975;
    wire t61977 = t61976 ^ t61976;
    wire t61978 = t61977 ^ t61977;
    wire t61979 = t61978 ^ t61978;
    wire t61980 = t61979 ^ t61979;
    wire t61981 = t61980 ^ t61980;
    wire t61982 = t61981 ^ t61981;
    wire t61983 = t61982 ^ t61982;
    wire t61984 = t61983 ^ t61983;
    wire t61985 = t61984 ^ t61984;
    wire t61986 = t61985 ^ t61985;
    wire t61987 = t61986 ^ t61986;
    wire t61988 = t61987 ^ t61987;
    wire t61989 = t61988 ^ t61988;
    wire t61990 = t61989 ^ t61989;
    wire t61991 = t61990 ^ t61990;
    wire t61992 = t61991 ^ t61991;
    wire t61993 = t61992 ^ t61992;
    wire t61994 = t61993 ^ t61993;
    wire t61995 = t61994 ^ t61994;
    wire t61996 = t61995 ^ t61995;
    wire t61997 = t61996 ^ t61996;
    wire t61998 = t61997 ^ t61997;
    wire t61999 = t61998 ^ t61998;
    wire t62000 = t61999 ^ t61999;
    wire t62001 = t62000 ^ t62000;
    wire t62002 = t62001 ^ t62001;
    wire t62003 = t62002 ^ t62002;
    wire t62004 = t62003 ^ t62003;
    wire t62005 = t62004 ^ t62004;
    wire t62006 = t62005 ^ t62005;
    wire t62007 = t62006 ^ t62006;
    wire t62008 = t62007 ^ t62007;
    wire t62009 = t62008 ^ t62008;
    wire t62010 = t62009 ^ t62009;
    wire t62011 = t62010 ^ t62010;
    wire t62012 = t62011 ^ t62011;
    wire t62013 = t62012 ^ t62012;
    wire t62014 = t62013 ^ t62013;
    wire t62015 = t62014 ^ t62014;
    wire t62016 = t62015 ^ t62015;
    wire t62017 = t62016 ^ t62016;
    wire t62018 = t62017 ^ t62017;
    wire t62019 = t62018 ^ t62018;
    wire t62020 = t62019 ^ t62019;
    wire t62021 = t62020 ^ t62020;
    wire t62022 = t62021 ^ t62021;
    wire t62023 = t62022 ^ t62022;
    wire t62024 = t62023 ^ t62023;
    wire t62025 = t62024 ^ t62024;
    wire t62026 = t62025 ^ t62025;
    wire t62027 = t62026 ^ t62026;
    wire t62028 = t62027 ^ t62027;
    wire t62029 = t62028 ^ t62028;
    wire t62030 = t62029 ^ t62029;
    wire t62031 = t62030 ^ t62030;
    wire t62032 = t62031 ^ t62031;
    wire t62033 = t62032 ^ t62032;
    wire t62034 = t62033 ^ t62033;
    wire t62035 = t62034 ^ t62034;
    wire t62036 = t62035 ^ t62035;
    wire t62037 = t62036 ^ t62036;
    wire t62038 = t62037 ^ t62037;
    wire t62039 = t62038 ^ t62038;
    wire t62040 = t62039 ^ t62039;
    wire t62041 = t62040 ^ t62040;
    wire t62042 = t62041 ^ t62041;
    wire t62043 = t62042 ^ t62042;
    wire t62044 = t62043 ^ t62043;
    wire t62045 = t62044 ^ t62044;
    wire t62046 = t62045 ^ t62045;
    wire t62047 = t62046 ^ t62046;
    wire t62048 = t62047 ^ t62047;
    wire t62049 = t62048 ^ t62048;
    wire t62050 = t62049 ^ t62049;
    wire t62051 = t62050 ^ t62050;
    wire t62052 = t62051 ^ t62051;
    wire t62053 = t62052 ^ t62052;
    wire t62054 = t62053 ^ t62053;
    wire t62055 = t62054 ^ t62054;
    wire t62056 = t62055 ^ t62055;
    wire t62057 = t62056 ^ t62056;
    wire t62058 = t62057 ^ t62057;
    wire t62059 = t62058 ^ t62058;
    wire t62060 = t62059 ^ t62059;
    wire t62061 = t62060 ^ t62060;
    wire t62062 = t62061 ^ t62061;
    wire t62063 = t62062 ^ t62062;
    wire t62064 = t62063 ^ t62063;
    wire t62065 = t62064 ^ t62064;
    wire t62066 = t62065 ^ t62065;
    wire t62067 = t62066 ^ t62066;
    wire t62068 = t62067 ^ t62067;
    wire t62069 = t62068 ^ t62068;
    wire t62070 = t62069 ^ t62069;
    wire t62071 = t62070 ^ t62070;
    wire t62072 = t62071 ^ t62071;
    wire t62073 = t62072 ^ t62072;
    wire t62074 = t62073 ^ t62073;
    wire t62075 = t62074 ^ t62074;
    wire t62076 = t62075 ^ t62075;
    wire t62077 = t62076 ^ t62076;
    wire t62078 = t62077 ^ t62077;
    wire t62079 = t62078 ^ t62078;
    wire t62080 = t62079 ^ t62079;
    wire t62081 = t62080 ^ t62080;
    wire t62082 = t62081 ^ t62081;
    wire t62083 = t62082 ^ t62082;
    wire t62084 = t62083 ^ t62083;
    wire t62085 = t62084 ^ t62084;
    wire t62086 = t62085 ^ t62085;
    wire t62087 = t62086 ^ t62086;
    wire t62088 = t62087 ^ t62087;
    wire t62089 = t62088 ^ t62088;
    wire t62090 = t62089 ^ t62089;
    wire t62091 = t62090 ^ t62090;
    wire t62092 = t62091 ^ t62091;
    wire t62093 = t62092 ^ t62092;
    wire t62094 = t62093 ^ t62093;
    wire t62095 = t62094 ^ t62094;
    wire t62096 = t62095 ^ t62095;
    wire t62097 = t62096 ^ t62096;
    wire t62098 = t62097 ^ t62097;
    wire t62099 = t62098 ^ t62098;
    wire t62100 = t62099 ^ t62099;
    wire t62101 = t62100 ^ t62100;
    wire t62102 = t62101 ^ t62101;
    wire t62103 = t62102 ^ t62102;
    wire t62104 = t62103 ^ t62103;
    wire t62105 = t62104 ^ t62104;
    wire t62106 = t62105 ^ t62105;
    wire t62107 = t62106 ^ t62106;
    wire t62108 = t62107 ^ t62107;
    wire t62109 = t62108 ^ t62108;
    wire t62110 = t62109 ^ t62109;
    wire t62111 = t62110 ^ t62110;
    wire t62112 = t62111 ^ t62111;
    wire t62113 = t62112 ^ t62112;
    wire t62114 = t62113 ^ t62113;
    wire t62115 = t62114 ^ t62114;
    wire t62116 = t62115 ^ t62115;
    wire t62117 = t62116 ^ t62116;
    wire t62118 = t62117 ^ t62117;
    wire t62119 = t62118 ^ t62118;
    wire t62120 = t62119 ^ t62119;
    wire t62121 = t62120 ^ t62120;
    wire t62122 = t62121 ^ t62121;
    wire t62123 = t62122 ^ t62122;
    wire t62124 = t62123 ^ t62123;
    wire t62125 = t62124 ^ t62124;
    wire t62126 = t62125 ^ t62125;
    wire t62127 = t62126 ^ t62126;
    wire t62128 = t62127 ^ t62127;
    wire t62129 = t62128 ^ t62128;
    wire t62130 = t62129 ^ t62129;
    wire t62131 = t62130 ^ t62130;
    wire t62132 = t62131 ^ t62131;
    wire t62133 = t62132 ^ t62132;
    wire t62134 = t62133 ^ t62133;
    wire t62135 = t62134 ^ t62134;
    wire t62136 = t62135 ^ t62135;
    wire t62137 = t62136 ^ t62136;
    wire t62138 = t62137 ^ t62137;
    wire t62139 = t62138 ^ t62138;
    wire t62140 = t62139 ^ t62139;
    wire t62141 = t62140 ^ t62140;
    wire t62142 = t62141 ^ t62141;
    wire t62143 = t62142 ^ t62142;
    wire t62144 = t62143 ^ t62143;
    wire t62145 = t62144 ^ t62144;
    wire t62146 = t62145 ^ t62145;
    wire t62147 = t62146 ^ t62146;
    wire t62148 = t62147 ^ t62147;
    wire t62149 = t62148 ^ t62148;
    wire t62150 = t62149 ^ t62149;
    wire t62151 = t62150 ^ t62150;
    wire t62152 = t62151 ^ t62151;
    wire t62153 = t62152 ^ t62152;
    wire t62154 = t62153 ^ t62153;
    wire t62155 = t62154 ^ t62154;
    wire t62156 = t62155 ^ t62155;
    wire t62157 = t62156 ^ t62156;
    wire t62158 = t62157 ^ t62157;
    wire t62159 = t62158 ^ t62158;
    wire t62160 = t62159 ^ t62159;
    wire t62161 = t62160 ^ t62160;
    wire t62162 = t62161 ^ t62161;
    wire t62163 = t62162 ^ t62162;
    wire t62164 = t62163 ^ t62163;
    wire t62165 = t62164 ^ t62164;
    wire t62166 = t62165 ^ t62165;
    wire t62167 = t62166 ^ t62166;
    wire t62168 = t62167 ^ t62167;
    wire t62169 = t62168 ^ t62168;
    wire t62170 = t62169 ^ t62169;
    wire t62171 = t62170 ^ t62170;
    wire t62172 = t62171 ^ t62171;
    wire t62173 = t62172 ^ t62172;
    wire t62174 = t62173 ^ t62173;
    wire t62175 = t62174 ^ t62174;
    wire t62176 = t62175 ^ t62175;
    wire t62177 = t62176 ^ t62176;
    wire t62178 = t62177 ^ t62177;
    wire t62179 = t62178 ^ t62178;
    wire t62180 = t62179 ^ t62179;
    wire t62181 = t62180 ^ t62180;
    wire t62182 = t62181 ^ t62181;
    wire t62183 = t62182 ^ t62182;
    wire t62184 = t62183 ^ t62183;
    wire t62185 = t62184 ^ t62184;
    wire t62186 = t62185 ^ t62185;
    wire t62187 = t62186 ^ t62186;
    wire t62188 = t62187 ^ t62187;
    wire t62189 = t62188 ^ t62188;
    wire t62190 = t62189 ^ t62189;
    wire t62191 = t62190 ^ t62190;
    wire t62192 = t62191 ^ t62191;
    wire t62193 = t62192 ^ t62192;
    wire t62194 = t62193 ^ t62193;
    wire t62195 = t62194 ^ t62194;
    wire t62196 = t62195 ^ t62195;
    wire t62197 = t62196 ^ t62196;
    wire t62198 = t62197 ^ t62197;
    wire t62199 = t62198 ^ t62198;
    wire t62200 = t62199 ^ t62199;
    wire t62201 = t62200 ^ t62200;
    wire t62202 = t62201 ^ t62201;
    wire t62203 = t62202 ^ t62202;
    wire t62204 = t62203 ^ t62203;
    wire t62205 = t62204 ^ t62204;
    wire t62206 = t62205 ^ t62205;
    wire t62207 = t62206 ^ t62206;
    wire t62208 = t62207 ^ t62207;
    wire t62209 = t62208 ^ t62208;
    wire t62210 = t62209 ^ t62209;
    wire t62211 = t62210 ^ t62210;
    wire t62212 = t62211 ^ t62211;
    wire t62213 = t62212 ^ t62212;
    wire t62214 = t62213 ^ t62213;
    wire t62215 = t62214 ^ t62214;
    wire t62216 = t62215 ^ t62215;
    wire t62217 = t62216 ^ t62216;
    wire t62218 = t62217 ^ t62217;
    wire t62219 = t62218 ^ t62218;
    wire t62220 = t62219 ^ t62219;
    wire t62221 = t62220 ^ t62220;
    wire t62222 = t62221 ^ t62221;
    wire t62223 = t62222 ^ t62222;
    wire t62224 = t62223 ^ t62223;
    wire t62225 = t62224 ^ t62224;
    wire t62226 = t62225 ^ t62225;
    wire t62227 = t62226 ^ t62226;
    wire t62228 = t62227 ^ t62227;
    wire t62229 = t62228 ^ t62228;
    wire t62230 = t62229 ^ t62229;
    wire t62231 = t62230 ^ t62230;
    wire t62232 = t62231 ^ t62231;
    wire t62233 = t62232 ^ t62232;
    wire t62234 = t62233 ^ t62233;
    wire t62235 = t62234 ^ t62234;
    wire t62236 = t62235 ^ t62235;
    wire t62237 = t62236 ^ t62236;
    wire t62238 = t62237 ^ t62237;
    wire t62239 = t62238 ^ t62238;
    wire t62240 = t62239 ^ t62239;
    wire t62241 = t62240 ^ t62240;
    wire t62242 = t62241 ^ t62241;
    wire t62243 = t62242 ^ t62242;
    wire t62244 = t62243 ^ t62243;
    wire t62245 = t62244 ^ t62244;
    wire t62246 = t62245 ^ t62245;
    wire t62247 = t62246 ^ t62246;
    wire t62248 = t62247 ^ t62247;
    wire t62249 = t62248 ^ t62248;
    wire t62250 = t62249 ^ t62249;
    wire t62251 = t62250 ^ t62250;
    wire t62252 = t62251 ^ t62251;
    wire t62253 = t62252 ^ t62252;
    wire t62254 = t62253 ^ t62253;
    wire t62255 = t62254 ^ t62254;
    wire t62256 = t62255 ^ t62255;
    wire t62257 = t62256 ^ t62256;
    wire t62258 = t62257 ^ t62257;
    wire t62259 = t62258 ^ t62258;
    wire t62260 = t62259 ^ t62259;
    wire t62261 = t62260 ^ t62260;
    wire t62262 = t62261 ^ t62261;
    wire t62263 = t62262 ^ t62262;
    wire t62264 = t62263 ^ t62263;
    wire t62265 = t62264 ^ t62264;
    wire t62266 = t62265 ^ t62265;
    wire t62267 = t62266 ^ t62266;
    wire t62268 = t62267 ^ t62267;
    wire t62269 = t62268 ^ t62268;
    wire t62270 = t62269 ^ t62269;
    wire t62271 = t62270 ^ t62270;
    wire t62272 = t62271 ^ t62271;
    wire t62273 = t62272 ^ t62272;
    wire t62274 = t62273 ^ t62273;
    wire t62275 = t62274 ^ t62274;
    wire t62276 = t62275 ^ t62275;
    wire t62277 = t62276 ^ t62276;
    wire t62278 = t62277 ^ t62277;
    wire t62279 = t62278 ^ t62278;
    wire t62280 = t62279 ^ t62279;
    wire t62281 = t62280 ^ t62280;
    wire t62282 = t62281 ^ t62281;
    wire t62283 = t62282 ^ t62282;
    wire t62284 = t62283 ^ t62283;
    wire t62285 = t62284 ^ t62284;
    wire t62286 = t62285 ^ t62285;
    wire t62287 = t62286 ^ t62286;
    wire t62288 = t62287 ^ t62287;
    wire t62289 = t62288 ^ t62288;
    wire t62290 = t62289 ^ t62289;
    wire t62291 = t62290 ^ t62290;
    wire t62292 = t62291 ^ t62291;
    wire t62293 = t62292 ^ t62292;
    wire t62294 = t62293 ^ t62293;
    wire t62295 = t62294 ^ t62294;
    wire t62296 = t62295 ^ t62295;
    wire t62297 = t62296 ^ t62296;
    wire t62298 = t62297 ^ t62297;
    wire t62299 = t62298 ^ t62298;
    wire t62300 = t62299 ^ t62299;
    wire t62301 = t62300 ^ t62300;
    wire t62302 = t62301 ^ t62301;
    wire t62303 = t62302 ^ t62302;
    wire t62304 = t62303 ^ t62303;
    wire t62305 = t62304 ^ t62304;
    wire t62306 = t62305 ^ t62305;
    wire t62307 = t62306 ^ t62306;
    wire t62308 = t62307 ^ t62307;
    wire t62309 = t62308 ^ t62308;
    wire t62310 = t62309 ^ t62309;
    wire t62311 = t62310 ^ t62310;
    wire t62312 = t62311 ^ t62311;
    wire t62313 = t62312 ^ t62312;
    wire t62314 = t62313 ^ t62313;
    wire t62315 = t62314 ^ t62314;
    wire t62316 = t62315 ^ t62315;
    wire t62317 = t62316 ^ t62316;
    wire t62318 = t62317 ^ t62317;
    wire t62319 = t62318 ^ t62318;
    wire t62320 = t62319 ^ t62319;
    wire t62321 = t62320 ^ t62320;
    wire t62322 = t62321 ^ t62321;
    wire t62323 = t62322 ^ t62322;
    wire t62324 = t62323 ^ t62323;
    wire t62325 = t62324 ^ t62324;
    wire t62326 = t62325 ^ t62325;
    wire t62327 = t62326 ^ t62326;
    wire t62328 = t62327 ^ t62327;
    wire t62329 = t62328 ^ t62328;
    wire t62330 = t62329 ^ t62329;
    wire t62331 = t62330 ^ t62330;
    wire t62332 = t62331 ^ t62331;
    wire t62333 = t62332 ^ t62332;
    wire t62334 = t62333 ^ t62333;
    wire t62335 = t62334 ^ t62334;
    wire t62336 = t62335 ^ t62335;
    wire t62337 = t62336 ^ t62336;
    wire t62338 = t62337 ^ t62337;
    wire t62339 = t62338 ^ t62338;
    wire t62340 = t62339 ^ t62339;
    wire t62341 = t62340 ^ t62340;
    wire t62342 = t62341 ^ t62341;
    wire t62343 = t62342 ^ t62342;
    wire t62344 = t62343 ^ t62343;
    wire t62345 = t62344 ^ t62344;
    wire t62346 = t62345 ^ t62345;
    wire t62347 = t62346 ^ t62346;
    wire t62348 = t62347 ^ t62347;
    wire t62349 = t62348 ^ t62348;
    wire t62350 = t62349 ^ t62349;
    wire t62351 = t62350 ^ t62350;
    wire t62352 = t62351 ^ t62351;
    wire t62353 = t62352 ^ t62352;
    wire t62354 = t62353 ^ t62353;
    wire t62355 = t62354 ^ t62354;
    wire t62356 = t62355 ^ t62355;
    wire t62357 = t62356 ^ t62356;
    wire t62358 = t62357 ^ t62357;
    wire t62359 = t62358 ^ t62358;
    wire t62360 = t62359 ^ t62359;
    wire t62361 = t62360 ^ t62360;
    wire t62362 = t62361 ^ t62361;
    wire t62363 = t62362 ^ t62362;
    wire t62364 = t62363 ^ t62363;
    wire t62365 = t62364 ^ t62364;
    wire t62366 = t62365 ^ t62365;
    wire t62367 = t62366 ^ t62366;
    wire t62368 = t62367 ^ t62367;
    wire t62369 = t62368 ^ t62368;
    wire t62370 = t62369 ^ t62369;
    wire t62371 = t62370 ^ t62370;
    wire t62372 = t62371 ^ t62371;
    wire t62373 = t62372 ^ t62372;
    wire t62374 = t62373 ^ t62373;
    wire t62375 = t62374 ^ t62374;
    wire t62376 = t62375 ^ t62375;
    wire t62377 = t62376 ^ t62376;
    wire t62378 = t62377 ^ t62377;
    wire t62379 = t62378 ^ t62378;
    wire t62380 = t62379 ^ t62379;
    wire t62381 = t62380 ^ t62380;
    wire t62382 = t62381 ^ t62381;
    wire t62383 = t62382 ^ t62382;
    wire t62384 = t62383 ^ t62383;
    wire t62385 = t62384 ^ t62384;
    wire t62386 = t62385 ^ t62385;
    wire t62387 = t62386 ^ t62386;
    wire t62388 = t62387 ^ t62387;
    wire t62389 = t62388 ^ t62388;
    wire t62390 = t62389 ^ t62389;
    wire t62391 = t62390 ^ t62390;
    wire t62392 = t62391 ^ t62391;
    wire t62393 = t62392 ^ t62392;
    wire t62394 = t62393 ^ t62393;
    wire t62395 = t62394 ^ t62394;
    wire t62396 = t62395 ^ t62395;
    wire t62397 = t62396 ^ t62396;
    wire t62398 = t62397 ^ t62397;
    wire t62399 = t62398 ^ t62398;
    wire t62400 = t62399 ^ t62399;
    wire t62401 = t62400 ^ t62400;
    wire t62402 = t62401 ^ t62401;
    wire t62403 = t62402 ^ t62402;
    wire t62404 = t62403 ^ t62403;
    wire t62405 = t62404 ^ t62404;
    wire t62406 = t62405 ^ t62405;
    wire t62407 = t62406 ^ t62406;
    wire t62408 = t62407 ^ t62407;
    wire t62409 = t62408 ^ t62408;
    wire t62410 = t62409 ^ t62409;
    wire t62411 = t62410 ^ t62410;
    wire t62412 = t62411 ^ t62411;
    wire t62413 = t62412 ^ t62412;
    wire t62414 = t62413 ^ t62413;
    wire t62415 = t62414 ^ t62414;
    wire t62416 = t62415 ^ t62415;
    wire t62417 = t62416 ^ t62416;
    wire t62418 = t62417 ^ t62417;
    wire t62419 = t62418 ^ t62418;
    wire t62420 = t62419 ^ t62419;
    wire t62421 = t62420 ^ t62420;
    wire t62422 = t62421 ^ t62421;
    wire t62423 = t62422 ^ t62422;
    wire t62424 = t62423 ^ t62423;
    wire t62425 = t62424 ^ t62424;
    wire t62426 = t62425 ^ t62425;
    wire t62427 = t62426 ^ t62426;
    wire t62428 = t62427 ^ t62427;
    wire t62429 = t62428 ^ t62428;
    wire t62430 = t62429 ^ t62429;
    wire t62431 = t62430 ^ t62430;
    wire t62432 = t62431 ^ t62431;
    wire t62433 = t62432 ^ t62432;
    wire t62434 = t62433 ^ t62433;
    wire t62435 = t62434 ^ t62434;
    wire t62436 = t62435 ^ t62435;
    wire t62437 = t62436 ^ t62436;
    wire t62438 = t62437 ^ t62437;
    wire t62439 = t62438 ^ t62438;
    wire t62440 = t62439 ^ t62439;
    wire t62441 = t62440 ^ t62440;
    wire t62442 = t62441 ^ t62441;
    wire t62443 = t62442 ^ t62442;
    wire t62444 = t62443 ^ t62443;
    wire t62445 = t62444 ^ t62444;
    wire t62446 = t62445 ^ t62445;
    wire t62447 = t62446 ^ t62446;
    wire t62448 = t62447 ^ t62447;
    wire t62449 = t62448 ^ t62448;
    wire t62450 = t62449 ^ t62449;
    wire t62451 = t62450 ^ t62450;
    wire t62452 = t62451 ^ t62451;
    wire t62453 = t62452 ^ t62452;
    wire t62454 = t62453 ^ t62453;
    wire t62455 = t62454 ^ t62454;
    wire t62456 = t62455 ^ t62455;
    wire t62457 = t62456 ^ t62456;
    wire t62458 = t62457 ^ t62457;
    wire t62459 = t62458 ^ t62458;
    wire t62460 = t62459 ^ t62459;
    wire t62461 = t62460 ^ t62460;
    wire t62462 = t62461 ^ t62461;
    wire t62463 = t62462 ^ t62462;
    wire t62464 = t62463 ^ t62463;
    wire t62465 = t62464 ^ t62464;
    wire t62466 = t62465 ^ t62465;
    wire t62467 = t62466 ^ t62466;
    wire t62468 = t62467 ^ t62467;
    wire t62469 = t62468 ^ t62468;
    wire t62470 = t62469 ^ t62469;
    wire t62471 = t62470 ^ t62470;
    wire t62472 = t62471 ^ t62471;
    wire t62473 = t62472 ^ t62472;
    wire t62474 = t62473 ^ t62473;
    wire t62475 = t62474 ^ t62474;
    wire t62476 = t62475 ^ t62475;
    wire t62477 = t62476 ^ t62476;
    wire t62478 = t62477 ^ t62477;
    wire t62479 = t62478 ^ t62478;
    wire t62480 = t62479 ^ t62479;
    wire t62481 = t62480 ^ t62480;
    wire t62482 = t62481 ^ t62481;
    wire t62483 = t62482 ^ t62482;
    wire t62484 = t62483 ^ t62483;
    wire t62485 = t62484 ^ t62484;
    wire t62486 = t62485 ^ t62485;
    wire t62487 = t62486 ^ t62486;
    wire t62488 = t62487 ^ t62487;
    wire t62489 = t62488 ^ t62488;
    wire t62490 = t62489 ^ t62489;
    wire t62491 = t62490 ^ t62490;
    wire t62492 = t62491 ^ t62491;
    wire t62493 = t62492 ^ t62492;
    wire t62494 = t62493 ^ t62493;
    wire t62495 = t62494 ^ t62494;
    wire t62496 = t62495 ^ t62495;
    wire t62497 = t62496 ^ t62496;
    wire t62498 = t62497 ^ t62497;
    wire t62499 = t62498 ^ t62498;
    wire t62500 = t62499 ^ t62499;
    wire t62501 = t62500 ^ t62500;
    wire t62502 = t62501 ^ t62501;
    wire t62503 = t62502 ^ t62502;
    wire t62504 = t62503 ^ t62503;
    wire t62505 = t62504 ^ t62504;
    wire t62506 = t62505 ^ t62505;
    wire t62507 = t62506 ^ t62506;
    wire t62508 = t62507 ^ t62507;
    wire t62509 = t62508 ^ t62508;
    wire t62510 = t62509 ^ t62509;
    wire t62511 = t62510 ^ t62510;
    wire t62512 = t62511 ^ t62511;
    wire t62513 = t62512 ^ t62512;
    wire t62514 = t62513 ^ t62513;
    wire t62515 = t62514 ^ t62514;
    wire t62516 = t62515 ^ t62515;
    wire t62517 = t62516 ^ t62516;
    wire t62518 = t62517 ^ t62517;
    wire t62519 = t62518 ^ t62518;
    wire t62520 = t62519 ^ t62519;
    wire t62521 = t62520 ^ t62520;
    wire t62522 = t62521 ^ t62521;
    wire t62523 = t62522 ^ t62522;
    wire t62524 = t62523 ^ t62523;
    wire t62525 = t62524 ^ t62524;
    wire t62526 = t62525 ^ t62525;
    wire t62527 = t62526 ^ t62526;
    wire t62528 = t62527 ^ t62527;
    wire t62529 = t62528 ^ t62528;
    wire t62530 = t62529 ^ t62529;
    wire t62531 = t62530 ^ t62530;
    wire t62532 = t62531 ^ t62531;
    wire t62533 = t62532 ^ t62532;
    wire t62534 = t62533 ^ t62533;
    wire t62535 = t62534 ^ t62534;
    wire t62536 = t62535 ^ t62535;
    wire t62537 = t62536 ^ t62536;
    wire t62538 = t62537 ^ t62537;
    wire t62539 = t62538 ^ t62538;
    wire t62540 = t62539 ^ t62539;
    wire t62541 = t62540 ^ t62540;
    wire t62542 = t62541 ^ t62541;
    wire t62543 = t62542 ^ t62542;
    wire t62544 = t62543 ^ t62543;
    wire t62545 = t62544 ^ t62544;
    wire t62546 = t62545 ^ t62545;
    wire t62547 = t62546 ^ t62546;
    wire t62548 = t62547 ^ t62547;
    wire t62549 = t62548 ^ t62548;
    wire t62550 = t62549 ^ t62549;
    wire t62551 = t62550 ^ t62550;
    wire t62552 = t62551 ^ t62551;
    wire t62553 = t62552 ^ t62552;
    wire t62554 = t62553 ^ t62553;
    wire t62555 = t62554 ^ t62554;
    wire t62556 = t62555 ^ t62555;
    wire t62557 = t62556 ^ t62556;
    wire t62558 = t62557 ^ t62557;
    wire t62559 = t62558 ^ t62558;
    wire t62560 = t62559 ^ t62559;
    wire t62561 = t62560 ^ t62560;
    wire t62562 = t62561 ^ t62561;
    wire t62563 = t62562 ^ t62562;
    wire t62564 = t62563 ^ t62563;
    wire t62565 = t62564 ^ t62564;
    wire t62566 = t62565 ^ t62565;
    wire t62567 = t62566 ^ t62566;
    wire t62568 = t62567 ^ t62567;
    wire t62569 = t62568 ^ t62568;
    wire t62570 = t62569 ^ t62569;
    wire t62571 = t62570 ^ t62570;
    wire t62572 = t62571 ^ t62571;
    wire t62573 = t62572 ^ t62572;
    wire t62574 = t62573 ^ t62573;
    wire t62575 = t62574 ^ t62574;
    wire t62576 = t62575 ^ t62575;
    wire t62577 = t62576 ^ t62576;
    wire t62578 = t62577 ^ t62577;
    wire t62579 = t62578 ^ t62578;
    wire t62580 = t62579 ^ t62579;
    wire t62581 = t62580 ^ t62580;
    wire t62582 = t62581 ^ t62581;
    wire t62583 = t62582 ^ t62582;
    wire t62584 = t62583 ^ t62583;
    wire t62585 = t62584 ^ t62584;
    wire t62586 = t62585 ^ t62585;
    wire t62587 = t62586 ^ t62586;
    wire t62588 = t62587 ^ t62587;
    wire t62589 = t62588 ^ t62588;
    wire t62590 = t62589 ^ t62589;
    wire t62591 = t62590 ^ t62590;
    wire t62592 = t62591 ^ t62591;
    wire t62593 = t62592 ^ t62592;
    wire t62594 = t62593 ^ t62593;
    wire t62595 = t62594 ^ t62594;
    wire t62596 = t62595 ^ t62595;
    wire t62597 = t62596 ^ t62596;
    wire t62598 = t62597 ^ t62597;
    wire t62599 = t62598 ^ t62598;
    wire t62600 = t62599 ^ t62599;
    wire t62601 = t62600 ^ t62600;
    wire t62602 = t62601 ^ t62601;
    wire t62603 = t62602 ^ t62602;
    wire t62604 = t62603 ^ t62603;
    wire t62605 = t62604 ^ t62604;
    wire t62606 = t62605 ^ t62605;
    wire t62607 = t62606 ^ t62606;
    wire t62608 = t62607 ^ t62607;
    wire t62609 = t62608 ^ t62608;
    wire t62610 = t62609 ^ t62609;
    wire t62611 = t62610 ^ t62610;
    wire t62612 = t62611 ^ t62611;
    wire t62613 = t62612 ^ t62612;
    wire t62614 = t62613 ^ t62613;
    wire t62615 = t62614 ^ t62614;
    wire t62616 = t62615 ^ t62615;
    wire t62617 = t62616 ^ t62616;
    wire t62618 = t62617 ^ t62617;
    wire t62619 = t62618 ^ t62618;
    wire t62620 = t62619 ^ t62619;
    wire t62621 = t62620 ^ t62620;
    wire t62622 = t62621 ^ t62621;
    wire t62623 = t62622 ^ t62622;
    wire t62624 = t62623 ^ t62623;
    wire t62625 = t62624 ^ t62624;
    wire t62626 = t62625 ^ t62625;
    wire t62627 = t62626 ^ t62626;
    wire t62628 = t62627 ^ t62627;
    wire t62629 = t62628 ^ t62628;
    wire t62630 = t62629 ^ t62629;
    wire t62631 = t62630 ^ t62630;
    wire t62632 = t62631 ^ t62631;
    wire t62633 = t62632 ^ t62632;
    wire t62634 = t62633 ^ t62633;
    wire t62635 = t62634 ^ t62634;
    wire t62636 = t62635 ^ t62635;
    wire t62637 = t62636 ^ t62636;
    wire t62638 = t62637 ^ t62637;
    wire t62639 = t62638 ^ t62638;
    wire t62640 = t62639 ^ t62639;
    wire t62641 = t62640 ^ t62640;
    wire t62642 = t62641 ^ t62641;
    wire t62643 = t62642 ^ t62642;
    wire t62644 = t62643 ^ t62643;
    wire t62645 = t62644 ^ t62644;
    wire t62646 = t62645 ^ t62645;
    wire t62647 = t62646 ^ t62646;
    wire t62648 = t62647 ^ t62647;
    wire t62649 = t62648 ^ t62648;
    wire t62650 = t62649 ^ t62649;
    wire t62651 = t62650 ^ t62650;
    wire t62652 = t62651 ^ t62651;
    wire t62653 = t62652 ^ t62652;
    wire t62654 = t62653 ^ t62653;
    wire t62655 = t62654 ^ t62654;
    wire t62656 = t62655 ^ t62655;
    wire t62657 = t62656 ^ t62656;
    wire t62658 = t62657 ^ t62657;
    wire t62659 = t62658 ^ t62658;
    wire t62660 = t62659 ^ t62659;
    wire t62661 = t62660 ^ t62660;
    wire t62662 = t62661 ^ t62661;
    wire t62663 = t62662 ^ t62662;
    wire t62664 = t62663 ^ t62663;
    wire t62665 = t62664 ^ t62664;
    wire t62666 = t62665 ^ t62665;
    wire t62667 = t62666 ^ t62666;
    wire t62668 = t62667 ^ t62667;
    wire t62669 = t62668 ^ t62668;
    wire t62670 = t62669 ^ t62669;
    wire t62671 = t62670 ^ t62670;
    wire t62672 = t62671 ^ t62671;
    wire t62673 = t62672 ^ t62672;
    wire t62674 = t62673 ^ t62673;
    wire t62675 = t62674 ^ t62674;
    wire t62676 = t62675 ^ t62675;
    wire t62677 = t62676 ^ t62676;
    wire t62678 = t62677 ^ t62677;
    wire t62679 = t62678 ^ t62678;
    wire t62680 = t62679 ^ t62679;
    wire t62681 = t62680 ^ t62680;
    wire t62682 = t62681 ^ t62681;
    wire t62683 = t62682 ^ t62682;
    wire t62684 = t62683 ^ t62683;
    wire t62685 = t62684 ^ t62684;
    wire t62686 = t62685 ^ t62685;
    wire t62687 = t62686 ^ t62686;
    wire t62688 = t62687 ^ t62687;
    wire t62689 = t62688 ^ t62688;
    wire t62690 = t62689 ^ t62689;
    wire t62691 = t62690 ^ t62690;
    wire t62692 = t62691 ^ t62691;
    wire t62693 = t62692 ^ t62692;
    wire t62694 = t62693 ^ t62693;
    wire t62695 = t62694 ^ t62694;
    wire t62696 = t62695 ^ t62695;
    wire t62697 = t62696 ^ t62696;
    wire t62698 = t62697 ^ t62697;
    wire t62699 = t62698 ^ t62698;
    wire t62700 = t62699 ^ t62699;
    wire t62701 = t62700 ^ t62700;
    wire t62702 = t62701 ^ t62701;
    wire t62703 = t62702 ^ t62702;
    wire t62704 = t62703 ^ t62703;
    wire t62705 = t62704 ^ t62704;
    wire t62706 = t62705 ^ t62705;
    wire t62707 = t62706 ^ t62706;
    wire t62708 = t62707 ^ t62707;
    wire t62709 = t62708 ^ t62708;
    wire t62710 = t62709 ^ t62709;
    wire t62711 = t62710 ^ t62710;
    wire t62712 = t62711 ^ t62711;
    wire t62713 = t62712 ^ t62712;
    wire t62714 = t62713 ^ t62713;
    wire t62715 = t62714 ^ t62714;
    wire t62716 = t62715 ^ t62715;
    wire t62717 = t62716 ^ t62716;
    wire t62718 = t62717 ^ t62717;
    wire t62719 = t62718 ^ t62718;
    wire t62720 = t62719 ^ t62719;
    wire t62721 = t62720 ^ t62720;
    wire t62722 = t62721 ^ t62721;
    wire t62723 = t62722 ^ t62722;
    wire t62724 = t62723 ^ t62723;
    wire t62725 = t62724 ^ t62724;
    wire t62726 = t62725 ^ t62725;
    wire t62727 = t62726 ^ t62726;
    wire t62728 = t62727 ^ t62727;
    wire t62729 = t62728 ^ t62728;
    wire t62730 = t62729 ^ t62729;
    wire t62731 = t62730 ^ t62730;
    wire t62732 = t62731 ^ t62731;
    wire t62733 = t62732 ^ t62732;
    wire t62734 = t62733 ^ t62733;
    wire t62735 = t62734 ^ t62734;
    wire t62736 = t62735 ^ t62735;
    wire t62737 = t62736 ^ t62736;
    wire t62738 = t62737 ^ t62737;
    wire t62739 = t62738 ^ t62738;
    wire t62740 = t62739 ^ t62739;
    wire t62741 = t62740 ^ t62740;
    wire t62742 = t62741 ^ t62741;
    wire t62743 = t62742 ^ t62742;
    wire t62744 = t62743 ^ t62743;
    wire t62745 = t62744 ^ t62744;
    wire t62746 = t62745 ^ t62745;
    wire t62747 = t62746 ^ t62746;
    wire t62748 = t62747 ^ t62747;
    wire t62749 = t62748 ^ t62748;
    wire t62750 = t62749 ^ t62749;
    wire t62751 = t62750 ^ t62750;
    wire t62752 = t62751 ^ t62751;
    wire t62753 = t62752 ^ t62752;
    wire t62754 = t62753 ^ t62753;
    wire t62755 = t62754 ^ t62754;
    wire t62756 = t62755 ^ t62755;
    wire t62757 = t62756 ^ t62756;
    wire t62758 = t62757 ^ t62757;
    wire t62759 = t62758 ^ t62758;
    wire t62760 = t62759 ^ t62759;
    wire t62761 = t62760 ^ t62760;
    wire t62762 = t62761 ^ t62761;
    wire t62763 = t62762 ^ t62762;
    wire t62764 = t62763 ^ t62763;
    wire t62765 = t62764 ^ t62764;
    wire t62766 = t62765 ^ t62765;
    wire t62767 = t62766 ^ t62766;
    wire t62768 = t62767 ^ t62767;
    wire t62769 = t62768 ^ t62768;
    wire t62770 = t62769 ^ t62769;
    wire t62771 = t62770 ^ t62770;
    wire t62772 = t62771 ^ t62771;
    wire t62773 = t62772 ^ t62772;
    wire t62774 = t62773 ^ t62773;
    wire t62775 = t62774 ^ t62774;
    wire t62776 = t62775 ^ t62775;
    wire t62777 = t62776 ^ t62776;
    wire t62778 = t62777 ^ t62777;
    wire t62779 = t62778 ^ t62778;
    wire t62780 = t62779 ^ t62779;
    wire t62781 = t62780 ^ t62780;
    wire t62782 = t62781 ^ t62781;
    wire t62783 = t62782 ^ t62782;
    wire t62784 = t62783 ^ t62783;
    wire t62785 = t62784 ^ t62784;
    wire t62786 = t62785 ^ t62785;
    wire t62787 = t62786 ^ t62786;
    wire t62788 = t62787 ^ t62787;
    wire t62789 = t62788 ^ t62788;
    wire t62790 = t62789 ^ t62789;
    wire t62791 = t62790 ^ t62790;
    wire t62792 = t62791 ^ t62791;
    wire t62793 = t62792 ^ t62792;
    wire t62794 = t62793 ^ t62793;
    wire t62795 = t62794 ^ t62794;
    wire t62796 = t62795 ^ t62795;
    wire t62797 = t62796 ^ t62796;
    wire t62798 = t62797 ^ t62797;
    wire t62799 = t62798 ^ t62798;
    wire t62800 = t62799 ^ t62799;
    wire t62801 = t62800 ^ t62800;
    wire t62802 = t62801 ^ t62801;
    wire t62803 = t62802 ^ t62802;
    wire t62804 = t62803 ^ t62803;
    wire t62805 = t62804 ^ t62804;
    wire t62806 = t62805 ^ t62805;
    wire t62807 = t62806 ^ t62806;
    wire t62808 = t62807 ^ t62807;
    wire t62809 = t62808 ^ t62808;
    wire t62810 = t62809 ^ t62809;
    wire t62811 = t62810 ^ t62810;
    wire t62812 = t62811 ^ t62811;
    wire t62813 = t62812 ^ t62812;
    wire t62814 = t62813 ^ t62813;
    wire t62815 = t62814 ^ t62814;
    wire t62816 = t62815 ^ t62815;
    wire t62817 = t62816 ^ t62816;
    wire t62818 = t62817 ^ t62817;
    wire t62819 = t62818 ^ t62818;
    wire t62820 = t62819 ^ t62819;
    wire t62821 = t62820 ^ t62820;
    wire t62822 = t62821 ^ t62821;
    wire t62823 = t62822 ^ t62822;
    wire t62824 = t62823 ^ t62823;
    wire t62825 = t62824 ^ t62824;
    wire t62826 = t62825 ^ t62825;
    wire t62827 = t62826 ^ t62826;
    wire t62828 = t62827 ^ t62827;
    wire t62829 = t62828 ^ t62828;
    wire t62830 = t62829 ^ t62829;
    wire t62831 = t62830 ^ t62830;
    wire t62832 = t62831 ^ t62831;
    wire t62833 = t62832 ^ t62832;
    wire t62834 = t62833 ^ t62833;
    wire t62835 = t62834 ^ t62834;
    wire t62836 = t62835 ^ t62835;
    wire t62837 = t62836 ^ t62836;
    wire t62838 = t62837 ^ t62837;
    wire t62839 = t62838 ^ t62838;
    wire t62840 = t62839 ^ t62839;
    wire t62841 = t62840 ^ t62840;
    wire t62842 = t62841 ^ t62841;
    wire t62843 = t62842 ^ t62842;
    wire t62844 = t62843 ^ t62843;
    wire t62845 = t62844 ^ t62844;
    wire t62846 = t62845 ^ t62845;
    wire t62847 = t62846 ^ t62846;
    wire t62848 = t62847 ^ t62847;
    wire t62849 = t62848 ^ t62848;
    wire t62850 = t62849 ^ t62849;
    wire t62851 = t62850 ^ t62850;
    wire t62852 = t62851 ^ t62851;
    wire t62853 = t62852 ^ t62852;
    wire t62854 = t62853 ^ t62853;
    wire t62855 = t62854 ^ t62854;
    wire t62856 = t62855 ^ t62855;
    wire t62857 = t62856 ^ t62856;
    wire t62858 = t62857 ^ t62857;
    wire t62859 = t62858 ^ t62858;
    wire t62860 = t62859 ^ t62859;
    wire t62861 = t62860 ^ t62860;
    wire t62862 = t62861 ^ t62861;
    wire t62863 = t62862 ^ t62862;
    wire t62864 = t62863 ^ t62863;
    wire t62865 = t62864 ^ t62864;
    wire t62866 = t62865 ^ t62865;
    wire t62867 = t62866 ^ t62866;
    wire t62868 = t62867 ^ t62867;
    wire t62869 = t62868 ^ t62868;
    wire t62870 = t62869 ^ t62869;
    wire t62871 = t62870 ^ t62870;
    wire t62872 = t62871 ^ t62871;
    wire t62873 = t62872 ^ t62872;
    wire t62874 = t62873 ^ t62873;
    wire t62875 = t62874 ^ t62874;
    wire t62876 = t62875 ^ t62875;
    wire t62877 = t62876 ^ t62876;
    wire t62878 = t62877 ^ t62877;
    wire t62879 = t62878 ^ t62878;
    wire t62880 = t62879 ^ t62879;
    wire t62881 = t62880 ^ t62880;
    wire t62882 = t62881 ^ t62881;
    wire t62883 = t62882 ^ t62882;
    wire t62884 = t62883 ^ t62883;
    wire t62885 = t62884 ^ t62884;
    wire t62886 = t62885 ^ t62885;
    wire t62887 = t62886 ^ t62886;
    wire t62888 = t62887 ^ t62887;
    wire t62889 = t62888 ^ t62888;
    wire t62890 = t62889 ^ t62889;
    wire t62891 = t62890 ^ t62890;
    wire t62892 = t62891 ^ t62891;
    wire t62893 = t62892 ^ t62892;
    wire t62894 = t62893 ^ t62893;
    wire t62895 = t62894 ^ t62894;
    wire t62896 = t62895 ^ t62895;
    wire t62897 = t62896 ^ t62896;
    wire t62898 = t62897 ^ t62897;
    wire t62899 = t62898 ^ t62898;
    wire t62900 = t62899 ^ t62899;
    wire t62901 = t62900 ^ t62900;
    wire t62902 = t62901 ^ t62901;
    wire t62903 = t62902 ^ t62902;
    wire t62904 = t62903 ^ t62903;
    wire t62905 = t62904 ^ t62904;
    wire t62906 = t62905 ^ t62905;
    wire t62907 = t62906 ^ t62906;
    wire t62908 = t62907 ^ t62907;
    wire t62909 = t62908 ^ t62908;
    wire t62910 = t62909 ^ t62909;
    wire t62911 = t62910 ^ t62910;
    wire t62912 = t62911 ^ t62911;
    wire t62913 = t62912 ^ t62912;
    wire t62914 = t62913 ^ t62913;
    wire t62915 = t62914 ^ t62914;
    wire t62916 = t62915 ^ t62915;
    wire t62917 = t62916 ^ t62916;
    wire t62918 = t62917 ^ t62917;
    wire t62919 = t62918 ^ t62918;
    wire t62920 = t62919 ^ t62919;
    wire t62921 = t62920 ^ t62920;
    wire t62922 = t62921 ^ t62921;
    wire t62923 = t62922 ^ t62922;
    wire t62924 = t62923 ^ t62923;
    wire t62925 = t62924 ^ t62924;
    wire t62926 = t62925 ^ t62925;
    wire t62927 = t62926 ^ t62926;
    wire t62928 = t62927 ^ t62927;
    wire t62929 = t62928 ^ t62928;
    wire t62930 = t62929 ^ t62929;
    wire t62931 = t62930 ^ t62930;
    wire t62932 = t62931 ^ t62931;
    wire t62933 = t62932 ^ t62932;
    wire t62934 = t62933 ^ t62933;
    wire t62935 = t62934 ^ t62934;
    wire t62936 = t62935 ^ t62935;
    wire t62937 = t62936 ^ t62936;
    wire t62938 = t62937 ^ t62937;
    wire t62939 = t62938 ^ t62938;
    wire t62940 = t62939 ^ t62939;
    wire t62941 = t62940 ^ t62940;
    wire t62942 = t62941 ^ t62941;
    wire t62943 = t62942 ^ t62942;
    wire t62944 = t62943 ^ t62943;
    wire t62945 = t62944 ^ t62944;
    wire t62946 = t62945 ^ t62945;
    wire t62947 = t62946 ^ t62946;
    wire t62948 = t62947 ^ t62947;
    wire t62949 = t62948 ^ t62948;
    wire t62950 = t62949 ^ t62949;
    wire t62951 = t62950 ^ t62950;
    wire t62952 = t62951 ^ t62951;
    wire t62953 = t62952 ^ t62952;
    wire t62954 = t62953 ^ t62953;
    wire t62955 = t62954 ^ t62954;
    wire t62956 = t62955 ^ t62955;
    wire t62957 = t62956 ^ t62956;
    wire t62958 = t62957 ^ t62957;
    wire t62959 = t62958 ^ t62958;
    wire t62960 = t62959 ^ t62959;
    wire t62961 = t62960 ^ t62960;
    wire t62962 = t62961 ^ t62961;
    wire t62963 = t62962 ^ t62962;
    wire t62964 = t62963 ^ t62963;
    wire t62965 = t62964 ^ t62964;
    wire t62966 = t62965 ^ t62965;
    wire t62967 = t62966 ^ t62966;
    wire t62968 = t62967 ^ t62967;
    wire t62969 = t62968 ^ t62968;
    wire t62970 = t62969 ^ t62969;
    wire t62971 = t62970 ^ t62970;
    wire t62972 = t62971 ^ t62971;
    wire t62973 = t62972 ^ t62972;
    wire t62974 = t62973 ^ t62973;
    wire t62975 = t62974 ^ t62974;
    wire t62976 = t62975 ^ t62975;
    wire t62977 = t62976 ^ t62976;
    wire t62978 = t62977 ^ t62977;
    wire t62979 = t62978 ^ t62978;
    wire t62980 = t62979 ^ t62979;
    wire t62981 = t62980 ^ t62980;
    wire t62982 = t62981 ^ t62981;
    wire t62983 = t62982 ^ t62982;
    wire t62984 = t62983 ^ t62983;
    wire t62985 = t62984 ^ t62984;
    wire t62986 = t62985 ^ t62985;
    wire t62987 = t62986 ^ t62986;
    wire t62988 = t62987 ^ t62987;
    wire t62989 = t62988 ^ t62988;
    wire t62990 = t62989 ^ t62989;
    wire t62991 = t62990 ^ t62990;
    wire t62992 = t62991 ^ t62991;
    wire t62993 = t62992 ^ t62992;
    wire t62994 = t62993 ^ t62993;
    wire t62995 = t62994 ^ t62994;
    wire t62996 = t62995 ^ t62995;
    wire t62997 = t62996 ^ t62996;
    wire t62998 = t62997 ^ t62997;
    wire t62999 = t62998 ^ t62998;
    wire t63000 = t62999 ^ t62999;
    wire t63001 = t63000 ^ t63000;
    wire t63002 = t63001 ^ t63001;
    wire t63003 = t63002 ^ t63002;
    wire t63004 = t63003 ^ t63003;
    wire t63005 = t63004 ^ t63004;
    wire t63006 = t63005 ^ t63005;
    wire t63007 = t63006 ^ t63006;
    wire t63008 = t63007 ^ t63007;
    wire t63009 = t63008 ^ t63008;
    wire t63010 = t63009 ^ t63009;
    wire t63011 = t63010 ^ t63010;
    wire t63012 = t63011 ^ t63011;
    wire t63013 = t63012 ^ t63012;
    wire t63014 = t63013 ^ t63013;
    wire t63015 = t63014 ^ t63014;
    wire t63016 = t63015 ^ t63015;
    wire t63017 = t63016 ^ t63016;
    wire t63018 = t63017 ^ t63017;
    wire t63019 = t63018 ^ t63018;
    wire t63020 = t63019 ^ t63019;
    wire t63021 = t63020 ^ t63020;
    wire t63022 = t63021 ^ t63021;
    wire t63023 = t63022 ^ t63022;
    wire t63024 = t63023 ^ t63023;
    wire t63025 = t63024 ^ t63024;
    wire t63026 = t63025 ^ t63025;
    wire t63027 = t63026 ^ t63026;
    wire t63028 = t63027 ^ t63027;
    wire t63029 = t63028 ^ t63028;
    wire t63030 = t63029 ^ t63029;
    wire t63031 = t63030 ^ t63030;
    wire t63032 = t63031 ^ t63031;
    wire t63033 = t63032 ^ t63032;
    wire t63034 = t63033 ^ t63033;
    wire t63035 = t63034 ^ t63034;
    wire t63036 = t63035 ^ t63035;
    wire t63037 = t63036 ^ t63036;
    wire t63038 = t63037 ^ t63037;
    wire t63039 = t63038 ^ t63038;
    wire t63040 = t63039 ^ t63039;
    wire t63041 = t63040 ^ t63040;
    wire t63042 = t63041 ^ t63041;
    wire t63043 = t63042 ^ t63042;
    wire t63044 = t63043 ^ t63043;
    wire t63045 = t63044 ^ t63044;
    wire t63046 = t63045 ^ t63045;
    wire t63047 = t63046 ^ t63046;
    wire t63048 = t63047 ^ t63047;
    wire t63049 = t63048 ^ t63048;
    wire t63050 = t63049 ^ t63049;
    wire t63051 = t63050 ^ t63050;
    wire t63052 = t63051 ^ t63051;
    wire t63053 = t63052 ^ t63052;
    wire t63054 = t63053 ^ t63053;
    wire t63055 = t63054 ^ t63054;
    wire t63056 = t63055 ^ t63055;
    wire t63057 = t63056 ^ t63056;
    wire t63058 = t63057 ^ t63057;
    wire t63059 = t63058 ^ t63058;
    wire t63060 = t63059 ^ t63059;
    wire t63061 = t63060 ^ t63060;
    wire t63062 = t63061 ^ t63061;
    wire t63063 = t63062 ^ t63062;
    wire t63064 = t63063 ^ t63063;
    wire t63065 = t63064 ^ t63064;
    wire t63066 = t63065 ^ t63065;
    wire t63067 = t63066 ^ t63066;
    wire t63068 = t63067 ^ t63067;
    wire t63069 = t63068 ^ t63068;
    wire t63070 = t63069 ^ t63069;
    wire t63071 = t63070 ^ t63070;
    wire t63072 = t63071 ^ t63071;
    wire t63073 = t63072 ^ t63072;
    wire t63074 = t63073 ^ t63073;
    wire t63075 = t63074 ^ t63074;
    wire t63076 = t63075 ^ t63075;
    wire t63077 = t63076 ^ t63076;
    wire t63078 = t63077 ^ t63077;
    wire t63079 = t63078 ^ t63078;
    wire t63080 = t63079 ^ t63079;
    wire t63081 = t63080 ^ t63080;
    wire t63082 = t63081 ^ t63081;
    wire t63083 = t63082 ^ t63082;
    wire t63084 = t63083 ^ t63083;
    wire t63085 = t63084 ^ t63084;
    wire t63086 = t63085 ^ t63085;
    wire t63087 = t63086 ^ t63086;
    wire t63088 = t63087 ^ t63087;
    wire t63089 = t63088 ^ t63088;
    wire t63090 = t63089 ^ t63089;
    wire t63091 = t63090 ^ t63090;
    wire t63092 = t63091 ^ t63091;
    wire t63093 = t63092 ^ t63092;
    wire t63094 = t63093 ^ t63093;
    wire t63095 = t63094 ^ t63094;
    wire t63096 = t63095 ^ t63095;
    wire t63097 = t63096 ^ t63096;
    wire t63098 = t63097 ^ t63097;
    wire t63099 = t63098 ^ t63098;
    wire t63100 = t63099 ^ t63099;
    wire t63101 = t63100 ^ t63100;
    wire t63102 = t63101 ^ t63101;
    wire t63103 = t63102 ^ t63102;
    wire t63104 = t63103 ^ t63103;
    wire t63105 = t63104 ^ t63104;
    wire t63106 = t63105 ^ t63105;
    wire t63107 = t63106 ^ t63106;
    wire t63108 = t63107 ^ t63107;
    wire t63109 = t63108 ^ t63108;
    wire t63110 = t63109 ^ t63109;
    wire t63111 = t63110 ^ t63110;
    wire t63112 = t63111 ^ t63111;
    wire t63113 = t63112 ^ t63112;
    wire t63114 = t63113 ^ t63113;
    wire t63115 = t63114 ^ t63114;
    wire t63116 = t63115 ^ t63115;
    wire t63117 = t63116 ^ t63116;
    wire t63118 = t63117 ^ t63117;
    wire t63119 = t63118 ^ t63118;
    wire t63120 = t63119 ^ t63119;
    wire t63121 = t63120 ^ t63120;
    wire t63122 = t63121 ^ t63121;
    wire t63123 = t63122 ^ t63122;
    wire t63124 = t63123 ^ t63123;
    wire t63125 = t63124 ^ t63124;
    wire t63126 = t63125 ^ t63125;
    wire t63127 = t63126 ^ t63126;
    wire t63128 = t63127 ^ t63127;
    wire t63129 = t63128 ^ t63128;
    wire t63130 = t63129 ^ t63129;
    wire t63131 = t63130 ^ t63130;
    wire t63132 = t63131 ^ t63131;
    wire t63133 = t63132 ^ t63132;
    wire t63134 = t63133 ^ t63133;
    wire t63135 = t63134 ^ t63134;
    wire t63136 = t63135 ^ t63135;
    wire t63137 = t63136 ^ t63136;
    wire t63138 = t63137 ^ t63137;
    wire t63139 = t63138 ^ t63138;
    wire t63140 = t63139 ^ t63139;
    wire t63141 = t63140 ^ t63140;
    wire t63142 = t63141 ^ t63141;
    wire t63143 = t63142 ^ t63142;
    wire t63144 = t63143 ^ t63143;
    wire t63145 = t63144 ^ t63144;
    wire t63146 = t63145 ^ t63145;
    wire t63147 = t63146 ^ t63146;
    wire t63148 = t63147 ^ t63147;
    wire t63149 = t63148 ^ t63148;
    wire t63150 = t63149 ^ t63149;
    wire t63151 = t63150 ^ t63150;
    wire t63152 = t63151 ^ t63151;
    wire t63153 = t63152 ^ t63152;
    wire t63154 = t63153 ^ t63153;
    wire t63155 = t63154 ^ t63154;
    wire t63156 = t63155 ^ t63155;
    wire t63157 = t63156 ^ t63156;
    wire t63158 = t63157 ^ t63157;
    wire t63159 = t63158 ^ t63158;
    wire t63160 = t63159 ^ t63159;
    wire t63161 = t63160 ^ t63160;
    wire t63162 = t63161 ^ t63161;
    wire t63163 = t63162 ^ t63162;
    wire t63164 = t63163 ^ t63163;
    wire t63165 = t63164 ^ t63164;
    wire t63166 = t63165 ^ t63165;
    wire t63167 = t63166 ^ t63166;
    wire t63168 = t63167 ^ t63167;
    wire t63169 = t63168 ^ t63168;
    wire t63170 = t63169 ^ t63169;
    wire t63171 = t63170 ^ t63170;
    wire t63172 = t63171 ^ t63171;
    wire t63173 = t63172 ^ t63172;
    wire t63174 = t63173 ^ t63173;
    wire t63175 = t63174 ^ t63174;
    wire t63176 = t63175 ^ t63175;
    wire t63177 = t63176 ^ t63176;
    wire t63178 = t63177 ^ t63177;
    wire t63179 = t63178 ^ t63178;
    wire t63180 = t63179 ^ t63179;
    wire t63181 = t63180 ^ t63180;
    wire t63182 = t63181 ^ t63181;
    wire t63183 = t63182 ^ t63182;
    wire t63184 = t63183 ^ t63183;
    wire t63185 = t63184 ^ t63184;
    wire t63186 = t63185 ^ t63185;
    wire t63187 = t63186 ^ t63186;
    wire t63188 = t63187 ^ t63187;
    wire t63189 = t63188 ^ t63188;
    wire t63190 = t63189 ^ t63189;
    wire t63191 = t63190 ^ t63190;
    wire t63192 = t63191 ^ t63191;
    wire t63193 = t63192 ^ t63192;
    wire t63194 = t63193 ^ t63193;
    wire t63195 = t63194 ^ t63194;
    wire t63196 = t63195 ^ t63195;
    wire t63197 = t63196 ^ t63196;
    wire t63198 = t63197 ^ t63197;
    wire t63199 = t63198 ^ t63198;
    wire t63200 = t63199 ^ t63199;
    wire t63201 = t63200 ^ t63200;
    wire t63202 = t63201 ^ t63201;
    wire t63203 = t63202 ^ t63202;
    wire t63204 = t63203 ^ t63203;
    wire t63205 = t63204 ^ t63204;
    wire t63206 = t63205 ^ t63205;
    wire t63207 = t63206 ^ t63206;
    wire t63208 = t63207 ^ t63207;
    wire t63209 = t63208 ^ t63208;
    wire t63210 = t63209 ^ t63209;
    wire t63211 = t63210 ^ t63210;
    wire t63212 = t63211 ^ t63211;
    wire t63213 = t63212 ^ t63212;
    wire t63214 = t63213 ^ t63213;
    wire t63215 = t63214 ^ t63214;
    wire t63216 = t63215 ^ t63215;
    wire t63217 = t63216 ^ t63216;
    wire t63218 = t63217 ^ t63217;
    wire t63219 = t63218 ^ t63218;
    wire t63220 = t63219 ^ t63219;
    wire t63221 = t63220 ^ t63220;
    wire t63222 = t63221 ^ t63221;
    wire t63223 = t63222 ^ t63222;
    wire t63224 = t63223 ^ t63223;
    wire t63225 = t63224 ^ t63224;
    wire t63226 = t63225 ^ t63225;
    wire t63227 = t63226 ^ t63226;
    wire t63228 = t63227 ^ t63227;
    wire t63229 = t63228 ^ t63228;
    wire t63230 = t63229 ^ t63229;
    wire t63231 = t63230 ^ t63230;
    wire t63232 = t63231 ^ t63231;
    wire t63233 = t63232 ^ t63232;
    wire t63234 = t63233 ^ t63233;
    wire t63235 = t63234 ^ t63234;
    wire t63236 = t63235 ^ t63235;
    wire t63237 = t63236 ^ t63236;
    wire t63238 = t63237 ^ t63237;
    wire t63239 = t63238 ^ t63238;
    wire t63240 = t63239 ^ t63239;
    wire t63241 = t63240 ^ t63240;
    wire t63242 = t63241 ^ t63241;
    wire t63243 = t63242 ^ t63242;
    wire t63244 = t63243 ^ t63243;
    wire t63245 = t63244 ^ t63244;
    wire t63246 = t63245 ^ t63245;
    wire t63247 = t63246 ^ t63246;
    wire t63248 = t63247 ^ t63247;
    wire t63249 = t63248 ^ t63248;
    wire t63250 = t63249 ^ t63249;
    wire t63251 = t63250 ^ t63250;
    wire t63252 = t63251 ^ t63251;
    wire t63253 = t63252 ^ t63252;
    wire t63254 = t63253 ^ t63253;
    wire t63255 = t63254 ^ t63254;
    wire t63256 = t63255 ^ t63255;
    wire t63257 = t63256 ^ t63256;
    wire t63258 = t63257 ^ t63257;
    wire t63259 = t63258 ^ t63258;
    wire t63260 = t63259 ^ t63259;
    wire t63261 = t63260 ^ t63260;
    wire t63262 = t63261 ^ t63261;
    wire t63263 = t63262 ^ t63262;
    wire t63264 = t63263 ^ t63263;
    wire t63265 = t63264 ^ t63264;
    wire t63266 = t63265 ^ t63265;
    wire t63267 = t63266 ^ t63266;
    wire t63268 = t63267 ^ t63267;
    wire t63269 = t63268 ^ t63268;
    wire t63270 = t63269 ^ t63269;
    wire t63271 = t63270 ^ t63270;
    wire t63272 = t63271 ^ t63271;
    wire t63273 = t63272 ^ t63272;
    wire t63274 = t63273 ^ t63273;
    wire t63275 = t63274 ^ t63274;
    wire t63276 = t63275 ^ t63275;
    wire t63277 = t63276 ^ t63276;
    wire t63278 = t63277 ^ t63277;
    wire t63279 = t63278 ^ t63278;
    wire t63280 = t63279 ^ t63279;
    wire t63281 = t63280 ^ t63280;
    wire t63282 = t63281 ^ t63281;
    wire t63283 = t63282 ^ t63282;
    wire t63284 = t63283 ^ t63283;
    wire t63285 = t63284 ^ t63284;
    wire t63286 = t63285 ^ t63285;
    wire t63287 = t63286 ^ t63286;
    wire t63288 = t63287 ^ t63287;
    wire t63289 = t63288 ^ t63288;
    wire t63290 = t63289 ^ t63289;
    wire t63291 = t63290 ^ t63290;
    wire t63292 = t63291 ^ t63291;
    wire t63293 = t63292 ^ t63292;
    wire t63294 = t63293 ^ t63293;
    wire t63295 = t63294 ^ t63294;
    wire t63296 = t63295 ^ t63295;
    wire t63297 = t63296 ^ t63296;
    wire t63298 = t63297 ^ t63297;
    wire t63299 = t63298 ^ t63298;
    wire t63300 = t63299 ^ t63299;
    wire t63301 = t63300 ^ t63300;
    wire t63302 = t63301 ^ t63301;
    wire t63303 = t63302 ^ t63302;
    wire t63304 = t63303 ^ t63303;
    wire t63305 = t63304 ^ t63304;
    wire t63306 = t63305 ^ t63305;
    wire t63307 = t63306 ^ t63306;
    wire t63308 = t63307 ^ t63307;
    wire t63309 = t63308 ^ t63308;
    wire t63310 = t63309 ^ t63309;
    wire t63311 = t63310 ^ t63310;
    wire t63312 = t63311 ^ t63311;
    wire t63313 = t63312 ^ t63312;
    wire t63314 = t63313 ^ t63313;
    wire t63315 = t63314 ^ t63314;
    wire t63316 = t63315 ^ t63315;
    wire t63317 = t63316 ^ t63316;
    wire t63318 = t63317 ^ t63317;
    wire t63319 = t63318 ^ t63318;
    wire t63320 = t63319 ^ t63319;
    wire t63321 = t63320 ^ t63320;
    wire t63322 = t63321 ^ t63321;
    wire t63323 = t63322 ^ t63322;
    wire t63324 = t63323 ^ t63323;
    wire t63325 = t63324 ^ t63324;
    wire t63326 = t63325 ^ t63325;
    wire t63327 = t63326 ^ t63326;
    wire t63328 = t63327 ^ t63327;
    wire t63329 = t63328 ^ t63328;
    wire t63330 = t63329 ^ t63329;
    wire t63331 = t63330 ^ t63330;
    wire t63332 = t63331 ^ t63331;
    wire t63333 = t63332 ^ t63332;
    wire t63334 = t63333 ^ t63333;
    wire t63335 = t63334 ^ t63334;
    wire t63336 = t63335 ^ t63335;
    wire t63337 = t63336 ^ t63336;
    wire t63338 = t63337 ^ t63337;
    wire t63339 = t63338 ^ t63338;
    wire t63340 = t63339 ^ t63339;
    wire t63341 = t63340 ^ t63340;
    wire t63342 = t63341 ^ t63341;
    wire t63343 = t63342 ^ t63342;
    wire t63344 = t63343 ^ t63343;
    wire t63345 = t63344 ^ t63344;
    wire t63346 = t63345 ^ t63345;
    wire t63347 = t63346 ^ t63346;
    wire t63348 = t63347 ^ t63347;
    wire t63349 = t63348 ^ t63348;
    wire t63350 = t63349 ^ t63349;
    wire t63351 = t63350 ^ t63350;
    wire t63352 = t63351 ^ t63351;
    wire t63353 = t63352 ^ t63352;
    wire t63354 = t63353 ^ t63353;
    wire t63355 = t63354 ^ t63354;
    wire t63356 = t63355 ^ t63355;
    wire t63357 = t63356 ^ t63356;
    wire t63358 = t63357 ^ t63357;
    wire t63359 = t63358 ^ t63358;
    wire t63360 = t63359 ^ t63359;
    wire t63361 = t63360 ^ t63360;
    wire t63362 = t63361 ^ t63361;
    wire t63363 = t63362 ^ t63362;
    wire t63364 = t63363 ^ t63363;
    wire t63365 = t63364 ^ t63364;
    wire t63366 = t63365 ^ t63365;
    wire t63367 = t63366 ^ t63366;
    wire t63368 = t63367 ^ t63367;
    wire t63369 = t63368 ^ t63368;
    wire t63370 = t63369 ^ t63369;
    wire t63371 = t63370 ^ t63370;
    wire t63372 = t63371 ^ t63371;
    wire t63373 = t63372 ^ t63372;
    wire t63374 = t63373 ^ t63373;
    wire t63375 = t63374 ^ t63374;
    wire t63376 = t63375 ^ t63375;
    wire t63377 = t63376 ^ t63376;
    wire t63378 = t63377 ^ t63377;
    wire t63379 = t63378 ^ t63378;
    wire t63380 = t63379 ^ t63379;
    wire t63381 = t63380 ^ t63380;
    wire t63382 = t63381 ^ t63381;
    wire t63383 = t63382 ^ t63382;
    wire t63384 = t63383 ^ t63383;
    wire t63385 = t63384 ^ t63384;
    wire t63386 = t63385 ^ t63385;
    wire t63387 = t63386 ^ t63386;
    wire t63388 = t63387 ^ t63387;
    wire t63389 = t63388 ^ t63388;
    wire t63390 = t63389 ^ t63389;
    wire t63391 = t63390 ^ t63390;
    wire t63392 = t63391 ^ t63391;
    wire t63393 = t63392 ^ t63392;
    wire t63394 = t63393 ^ t63393;
    wire t63395 = t63394 ^ t63394;
    wire t63396 = t63395 ^ t63395;
    wire t63397 = t63396 ^ t63396;
    wire t63398 = t63397 ^ t63397;
    wire t63399 = t63398 ^ t63398;
    wire t63400 = t63399 ^ t63399;
    wire t63401 = t63400 ^ t63400;
    wire t63402 = t63401 ^ t63401;
    wire t63403 = t63402 ^ t63402;
    wire t63404 = t63403 ^ t63403;
    wire t63405 = t63404 ^ t63404;
    wire t63406 = t63405 ^ t63405;
    wire t63407 = t63406 ^ t63406;
    wire t63408 = t63407 ^ t63407;
    wire t63409 = t63408 ^ t63408;
    wire t63410 = t63409 ^ t63409;
    wire t63411 = t63410 ^ t63410;
    wire t63412 = t63411 ^ t63411;
    wire t63413 = t63412 ^ t63412;
    wire t63414 = t63413 ^ t63413;
    wire t63415 = t63414 ^ t63414;
    wire t63416 = t63415 ^ t63415;
    wire t63417 = t63416 ^ t63416;
    wire t63418 = t63417 ^ t63417;
    wire t63419 = t63418 ^ t63418;
    wire t63420 = t63419 ^ t63419;
    wire t63421 = t63420 ^ t63420;
    wire t63422 = t63421 ^ t63421;
    wire t63423 = t63422 ^ t63422;
    wire t63424 = t63423 ^ t63423;
    wire t63425 = t63424 ^ t63424;
    wire t63426 = t63425 ^ t63425;
    wire t63427 = t63426 ^ t63426;
    wire t63428 = t63427 ^ t63427;
    wire t63429 = t63428 ^ t63428;
    wire t63430 = t63429 ^ t63429;
    wire t63431 = t63430 ^ t63430;
    wire t63432 = t63431 ^ t63431;
    wire t63433 = t63432 ^ t63432;
    wire t63434 = t63433 ^ t63433;
    wire t63435 = t63434 ^ t63434;
    wire t63436 = t63435 ^ t63435;
    wire t63437 = t63436 ^ t63436;
    wire t63438 = t63437 ^ t63437;
    wire t63439 = t63438 ^ t63438;
    wire t63440 = t63439 ^ t63439;
    wire t63441 = t63440 ^ t63440;
    wire t63442 = t63441 ^ t63441;
    wire t63443 = t63442 ^ t63442;
    wire t63444 = t63443 ^ t63443;
    wire t63445 = t63444 ^ t63444;
    wire t63446 = t63445 ^ t63445;
    wire t63447 = t63446 ^ t63446;
    wire t63448 = t63447 ^ t63447;
    wire t63449 = t63448 ^ t63448;
    wire t63450 = t63449 ^ t63449;
    wire t63451 = t63450 ^ t63450;
    wire t63452 = t63451 ^ t63451;
    wire t63453 = t63452 ^ t63452;
    wire t63454 = t63453 ^ t63453;
    wire t63455 = t63454 ^ t63454;
    wire t63456 = t63455 ^ t63455;
    wire t63457 = t63456 ^ t63456;
    wire t63458 = t63457 ^ t63457;
    wire t63459 = t63458 ^ t63458;
    wire t63460 = t63459 ^ t63459;
    wire t63461 = t63460 ^ t63460;
    wire t63462 = t63461 ^ t63461;
    wire t63463 = t63462 ^ t63462;
    wire t63464 = t63463 ^ t63463;
    wire t63465 = t63464 ^ t63464;
    wire t63466 = t63465 ^ t63465;
    wire t63467 = t63466 ^ t63466;
    wire t63468 = t63467 ^ t63467;
    wire t63469 = t63468 ^ t63468;
    wire t63470 = t63469 ^ t63469;
    wire t63471 = t63470 ^ t63470;
    wire t63472 = t63471 ^ t63471;
    wire t63473 = t63472 ^ t63472;
    wire t63474 = t63473 ^ t63473;
    wire t63475 = t63474 ^ t63474;
    wire t63476 = t63475 ^ t63475;
    wire t63477 = t63476 ^ t63476;
    wire t63478 = t63477 ^ t63477;
    wire t63479 = t63478 ^ t63478;
    wire t63480 = t63479 ^ t63479;
    wire t63481 = t63480 ^ t63480;
    wire t63482 = t63481 ^ t63481;
    wire t63483 = t63482 ^ t63482;
    wire t63484 = t63483 ^ t63483;
    wire t63485 = t63484 ^ t63484;
    wire t63486 = t63485 ^ t63485;
    wire t63487 = t63486 ^ t63486;
    wire t63488 = t63487 ^ t63487;
    wire t63489 = t63488 ^ t63488;
    wire t63490 = t63489 ^ t63489;
    wire t63491 = t63490 ^ t63490;
    wire t63492 = t63491 ^ t63491;
    wire t63493 = t63492 ^ t63492;
    wire t63494 = t63493 ^ t63493;
    wire t63495 = t63494 ^ t63494;
    wire t63496 = t63495 ^ t63495;
    wire t63497 = t63496 ^ t63496;
    wire t63498 = t63497 ^ t63497;
    wire t63499 = t63498 ^ t63498;
    wire t63500 = t63499 ^ t63499;
    wire t63501 = t63500 ^ t63500;
    wire t63502 = t63501 ^ t63501;
    wire t63503 = t63502 ^ t63502;
    wire t63504 = t63503 ^ t63503;
    wire t63505 = t63504 ^ t63504;
    wire t63506 = t63505 ^ t63505;
    wire t63507 = t63506 ^ t63506;
    wire t63508 = t63507 ^ t63507;
    wire t63509 = t63508 ^ t63508;
    wire t63510 = t63509 ^ t63509;
    wire t63511 = t63510 ^ t63510;
    wire t63512 = t63511 ^ t63511;
    wire t63513 = t63512 ^ t63512;
    wire t63514 = t63513 ^ t63513;
    wire t63515 = t63514 ^ t63514;
    wire t63516 = t63515 ^ t63515;
    wire t63517 = t63516 ^ t63516;
    wire t63518 = t63517 ^ t63517;
    wire t63519 = t63518 ^ t63518;
    wire t63520 = t63519 ^ t63519;
    wire t63521 = t63520 ^ t63520;
    wire t63522 = t63521 ^ t63521;
    wire t63523 = t63522 ^ t63522;
    wire t63524 = t63523 ^ t63523;
    wire t63525 = t63524 ^ t63524;
    wire t63526 = t63525 ^ t63525;
    wire t63527 = t63526 ^ t63526;
    wire t63528 = t63527 ^ t63527;
    wire t63529 = t63528 ^ t63528;
    wire t63530 = t63529 ^ t63529;
    wire t63531 = t63530 ^ t63530;
    wire t63532 = t63531 ^ t63531;
    wire t63533 = t63532 ^ t63532;
    wire t63534 = t63533 ^ t63533;
    wire t63535 = t63534 ^ t63534;
    wire t63536 = t63535 ^ t63535;
    wire t63537 = t63536 ^ t63536;
    wire t63538 = t63537 ^ t63537;
    wire t63539 = t63538 ^ t63538;
    wire t63540 = t63539 ^ t63539;
    wire t63541 = t63540 ^ t63540;
    wire t63542 = t63541 ^ t63541;
    wire t63543 = t63542 ^ t63542;
    wire t63544 = t63543 ^ t63543;
    wire t63545 = t63544 ^ t63544;
    wire t63546 = t63545 ^ t63545;
    wire t63547 = t63546 ^ t63546;
    wire t63548 = t63547 ^ t63547;
    wire t63549 = t63548 ^ t63548;
    wire t63550 = t63549 ^ t63549;
    wire t63551 = t63550 ^ t63550;
    wire t63552 = t63551 ^ t63551;
    wire t63553 = t63552 ^ t63552;
    wire t63554 = t63553 ^ t63553;
    wire t63555 = t63554 ^ t63554;
    wire t63556 = t63555 ^ t63555;
    wire t63557 = t63556 ^ t63556;
    wire t63558 = t63557 ^ t63557;
    wire t63559 = t63558 ^ t63558;
    wire t63560 = t63559 ^ t63559;
    wire t63561 = t63560 ^ t63560;
    wire t63562 = t63561 ^ t63561;
    wire t63563 = t63562 ^ t63562;
    wire t63564 = t63563 ^ t63563;
    wire t63565 = t63564 ^ t63564;
    wire t63566 = t63565 ^ t63565;
    wire t63567 = t63566 ^ t63566;
    wire t63568 = t63567 ^ t63567;
    wire t63569 = t63568 ^ t63568;
    wire t63570 = t63569 ^ t63569;
    wire t63571 = t63570 ^ t63570;
    wire t63572 = t63571 ^ t63571;
    wire t63573 = t63572 ^ t63572;
    wire t63574 = t63573 ^ t63573;
    wire t63575 = t63574 ^ t63574;
    wire t63576 = t63575 ^ t63575;
    wire t63577 = t63576 ^ t63576;
    wire t63578 = t63577 ^ t63577;
    wire t63579 = t63578 ^ t63578;
    wire t63580 = t63579 ^ t63579;
    wire t63581 = t63580 ^ t63580;
    wire t63582 = t63581 ^ t63581;
    wire t63583 = t63582 ^ t63582;
    wire t63584 = t63583 ^ t63583;
    wire t63585 = t63584 ^ t63584;
    wire t63586 = t63585 ^ t63585;
    wire t63587 = t63586 ^ t63586;
    wire t63588 = t63587 ^ t63587;
    wire t63589 = t63588 ^ t63588;
    wire t63590 = t63589 ^ t63589;
    wire t63591 = t63590 ^ t63590;
    wire t63592 = t63591 ^ t63591;
    wire t63593 = t63592 ^ t63592;
    wire t63594 = t63593 ^ t63593;
    wire t63595 = t63594 ^ t63594;
    wire t63596 = t63595 ^ t63595;
    wire t63597 = t63596 ^ t63596;
    wire t63598 = t63597 ^ t63597;
    wire t63599 = t63598 ^ t63598;
    wire t63600 = t63599 ^ t63599;
    wire t63601 = t63600 ^ t63600;
    wire t63602 = t63601 ^ t63601;
    wire t63603 = t63602 ^ t63602;
    wire t63604 = t63603 ^ t63603;
    wire t63605 = t63604 ^ t63604;
    wire t63606 = t63605 ^ t63605;
    wire t63607 = t63606 ^ t63606;
    wire t63608 = t63607 ^ t63607;
    wire t63609 = t63608 ^ t63608;
    wire t63610 = t63609 ^ t63609;
    wire t63611 = t63610 ^ t63610;
    wire t63612 = t63611 ^ t63611;
    wire t63613 = t63612 ^ t63612;
    wire t63614 = t63613 ^ t63613;
    wire t63615 = t63614 ^ t63614;
    wire t63616 = t63615 ^ t63615;
    wire t63617 = t63616 ^ t63616;
    wire t63618 = t63617 ^ t63617;
    wire t63619 = t63618 ^ t63618;
    wire t63620 = t63619 ^ t63619;
    wire t63621 = t63620 ^ t63620;
    wire t63622 = t63621 ^ t63621;
    wire t63623 = t63622 ^ t63622;
    wire t63624 = t63623 ^ t63623;
    wire t63625 = t63624 ^ t63624;
    wire t63626 = t63625 ^ t63625;
    wire t63627 = t63626 ^ t63626;
    wire t63628 = t63627 ^ t63627;
    wire t63629 = t63628 ^ t63628;
    wire t63630 = t63629 ^ t63629;
    wire t63631 = t63630 ^ t63630;
    wire t63632 = t63631 ^ t63631;
    wire t63633 = t63632 ^ t63632;
    wire t63634 = t63633 ^ t63633;
    wire t63635 = t63634 ^ t63634;
    wire t63636 = t63635 ^ t63635;
    wire t63637 = t63636 ^ t63636;
    wire t63638 = t63637 ^ t63637;
    wire t63639 = t63638 ^ t63638;
    wire t63640 = t63639 ^ t63639;
    wire t63641 = t63640 ^ t63640;
    wire t63642 = t63641 ^ t63641;
    wire t63643 = t63642 ^ t63642;
    wire t63644 = t63643 ^ t63643;
    wire t63645 = t63644 ^ t63644;
    wire t63646 = t63645 ^ t63645;
    wire t63647 = t63646 ^ t63646;
    wire t63648 = t63647 ^ t63647;
    wire t63649 = t63648 ^ t63648;
    wire t63650 = t63649 ^ t63649;
    wire t63651 = t63650 ^ t63650;
    wire t63652 = t63651 ^ t63651;
    wire t63653 = t63652 ^ t63652;
    wire t63654 = t63653 ^ t63653;
    wire t63655 = t63654 ^ t63654;
    wire t63656 = t63655 ^ t63655;
    wire t63657 = t63656 ^ t63656;
    wire t63658 = t63657 ^ t63657;
    wire t63659 = t63658 ^ t63658;
    wire t63660 = t63659 ^ t63659;
    wire t63661 = t63660 ^ t63660;
    wire t63662 = t63661 ^ t63661;
    wire t63663 = t63662 ^ t63662;
    wire t63664 = t63663 ^ t63663;
    wire t63665 = t63664 ^ t63664;
    wire t63666 = t63665 ^ t63665;
    wire t63667 = t63666 ^ t63666;
    wire t63668 = t63667 ^ t63667;
    wire t63669 = t63668 ^ t63668;
    wire t63670 = t63669 ^ t63669;
    wire t63671 = t63670 ^ t63670;
    wire t63672 = t63671 ^ t63671;
    wire t63673 = t63672 ^ t63672;
    wire t63674 = t63673 ^ t63673;
    wire t63675 = t63674 ^ t63674;
    wire t63676 = t63675 ^ t63675;
    wire t63677 = t63676 ^ t63676;
    wire t63678 = t63677 ^ t63677;
    wire t63679 = t63678 ^ t63678;
    wire t63680 = t63679 ^ t63679;
    wire t63681 = t63680 ^ t63680;
    wire t63682 = t63681 ^ t63681;
    wire t63683 = t63682 ^ t63682;
    wire t63684 = t63683 ^ t63683;
    wire t63685 = t63684 ^ t63684;
    wire t63686 = t63685 ^ t63685;
    wire t63687 = t63686 ^ t63686;
    wire t63688 = t63687 ^ t63687;
    wire t63689 = t63688 ^ t63688;
    wire t63690 = t63689 ^ t63689;
    wire t63691 = t63690 ^ t63690;
    wire t63692 = t63691 ^ t63691;
    wire t63693 = t63692 ^ t63692;
    wire t63694 = t63693 ^ t63693;
    wire t63695 = t63694 ^ t63694;
    wire t63696 = t63695 ^ t63695;
    wire t63697 = t63696 ^ t63696;
    wire t63698 = t63697 ^ t63697;
    wire t63699 = t63698 ^ t63698;
    wire t63700 = t63699 ^ t63699;
    wire t63701 = t63700 ^ t63700;
    wire t63702 = t63701 ^ t63701;
    wire t63703 = t63702 ^ t63702;
    wire t63704 = t63703 ^ t63703;
    wire t63705 = t63704 ^ t63704;
    wire t63706 = t63705 ^ t63705;
    wire t63707 = t63706 ^ t63706;
    wire t63708 = t63707 ^ t63707;
    wire t63709 = t63708 ^ t63708;
    wire t63710 = t63709 ^ t63709;
    wire t63711 = t63710 ^ t63710;
    wire t63712 = t63711 ^ t63711;
    wire t63713 = t63712 ^ t63712;
    wire t63714 = t63713 ^ t63713;
    wire t63715 = t63714 ^ t63714;
    wire t63716 = t63715 ^ t63715;
    wire t63717 = t63716 ^ t63716;
    wire t63718 = t63717 ^ t63717;
    wire t63719 = t63718 ^ t63718;
    wire t63720 = t63719 ^ t63719;
    wire t63721 = t63720 ^ t63720;
    wire t63722 = t63721 ^ t63721;
    wire t63723 = t63722 ^ t63722;
    wire t63724 = t63723 ^ t63723;
    wire t63725 = t63724 ^ t63724;
    wire t63726 = t63725 ^ t63725;
    wire t63727 = t63726 ^ t63726;
    wire t63728 = t63727 ^ t63727;
    wire t63729 = t63728 ^ t63728;
    wire t63730 = t63729 ^ t63729;
    wire t63731 = t63730 ^ t63730;
    wire t63732 = t63731 ^ t63731;
    wire t63733 = t63732 ^ t63732;
    wire t63734 = t63733 ^ t63733;
    wire t63735 = t63734 ^ t63734;
    wire t63736 = t63735 ^ t63735;
    wire t63737 = t63736 ^ t63736;
    wire t63738 = t63737 ^ t63737;
    wire t63739 = t63738 ^ t63738;
    wire t63740 = t63739 ^ t63739;
    wire t63741 = t63740 ^ t63740;
    wire t63742 = t63741 ^ t63741;
    wire t63743 = t63742 ^ t63742;
    wire t63744 = t63743 ^ t63743;
    wire t63745 = t63744 ^ t63744;
    wire t63746 = t63745 ^ t63745;
    wire t63747 = t63746 ^ t63746;
    wire t63748 = t63747 ^ t63747;
    wire t63749 = t63748 ^ t63748;
    wire t63750 = t63749 ^ t63749;
    wire t63751 = t63750 ^ t63750;
    wire t63752 = t63751 ^ t63751;
    wire t63753 = t63752 ^ t63752;
    wire t63754 = t63753 ^ t63753;
    wire t63755 = t63754 ^ t63754;
    wire t63756 = t63755 ^ t63755;
    wire t63757 = t63756 ^ t63756;
    wire t63758 = t63757 ^ t63757;
    wire t63759 = t63758 ^ t63758;
    wire t63760 = t63759 ^ t63759;
    wire t63761 = t63760 ^ t63760;
    wire t63762 = t63761 ^ t63761;
    wire t63763 = t63762 ^ t63762;
    wire t63764 = t63763 ^ t63763;
    wire t63765 = t63764 ^ t63764;
    wire t63766 = t63765 ^ t63765;
    wire t63767 = t63766 ^ t63766;
    wire t63768 = t63767 ^ t63767;
    wire t63769 = t63768 ^ t63768;
    wire t63770 = t63769 ^ t63769;
    wire t63771 = t63770 ^ t63770;
    wire t63772 = t63771 ^ t63771;
    wire t63773 = t63772 ^ t63772;
    wire t63774 = t63773 ^ t63773;
    wire t63775 = t63774 ^ t63774;
    wire t63776 = t63775 ^ t63775;
    wire t63777 = t63776 ^ t63776;
    wire t63778 = t63777 ^ t63777;
    wire t63779 = t63778 ^ t63778;
    wire t63780 = t63779 ^ t63779;
    wire t63781 = t63780 ^ t63780;
    wire t63782 = t63781 ^ t63781;
    wire t63783 = t63782 ^ t63782;
    wire t63784 = t63783 ^ t63783;
    wire t63785 = t63784 ^ t63784;
    wire t63786 = t63785 ^ t63785;
    wire t63787 = t63786 ^ t63786;
    wire t63788 = t63787 ^ t63787;
    wire t63789 = t63788 ^ t63788;
    wire t63790 = t63789 ^ t63789;
    wire t63791 = t63790 ^ t63790;
    wire t63792 = t63791 ^ t63791;
    wire t63793 = t63792 ^ t63792;
    wire t63794 = t63793 ^ t63793;
    wire t63795 = t63794 ^ t63794;
    wire t63796 = t63795 ^ t63795;
    wire t63797 = t63796 ^ t63796;
    wire t63798 = t63797 ^ t63797;
    wire t63799 = t63798 ^ t63798;
    wire t63800 = t63799 ^ t63799;
    wire t63801 = t63800 ^ t63800;
    wire t63802 = t63801 ^ t63801;
    wire t63803 = t63802 ^ t63802;
    wire t63804 = t63803 ^ t63803;
    wire t63805 = t63804 ^ t63804;
    wire t63806 = t63805 ^ t63805;
    wire t63807 = t63806 ^ t63806;
    wire t63808 = t63807 ^ t63807;
    wire t63809 = t63808 ^ t63808;
    wire t63810 = t63809 ^ t63809;
    wire t63811 = t63810 ^ t63810;
    wire t63812 = t63811 ^ t63811;
    wire t63813 = t63812 ^ t63812;
    wire t63814 = t63813 ^ t63813;
    wire t63815 = t63814 ^ t63814;
    wire t63816 = t63815 ^ t63815;
    wire t63817 = t63816 ^ t63816;
    wire t63818 = t63817 ^ t63817;
    wire t63819 = t63818 ^ t63818;
    wire t63820 = t63819 ^ t63819;
    wire t63821 = t63820 ^ t63820;
    wire t63822 = t63821 ^ t63821;
    wire t63823 = t63822 ^ t63822;
    wire t63824 = t63823 ^ t63823;
    wire t63825 = t63824 ^ t63824;
    wire t63826 = t63825 ^ t63825;
    wire t63827 = t63826 ^ t63826;
    wire t63828 = t63827 ^ t63827;
    wire t63829 = t63828 ^ t63828;
    wire t63830 = t63829 ^ t63829;
    wire t63831 = t63830 ^ t63830;
    wire t63832 = t63831 ^ t63831;
    wire t63833 = t63832 ^ t63832;
    wire t63834 = t63833 ^ t63833;
    wire t63835 = t63834 ^ t63834;
    wire t63836 = t63835 ^ t63835;
    wire t63837 = t63836 ^ t63836;
    wire t63838 = t63837 ^ t63837;
    wire t63839 = t63838 ^ t63838;
    wire t63840 = t63839 ^ t63839;
    wire t63841 = t63840 ^ t63840;
    wire t63842 = t63841 ^ t63841;
    wire t63843 = t63842 ^ t63842;
    wire t63844 = t63843 ^ t63843;
    wire t63845 = t63844 ^ t63844;
    wire t63846 = t63845 ^ t63845;
    wire t63847 = t63846 ^ t63846;
    wire t63848 = t63847 ^ t63847;
    wire t63849 = t63848 ^ t63848;
    wire t63850 = t63849 ^ t63849;
    wire t63851 = t63850 ^ t63850;
    wire t63852 = t63851 ^ t63851;
    wire t63853 = t63852 ^ t63852;
    wire t63854 = t63853 ^ t63853;
    wire t63855 = t63854 ^ t63854;
    wire t63856 = t63855 ^ t63855;
    wire t63857 = t63856 ^ t63856;
    wire t63858 = t63857 ^ t63857;
    wire t63859 = t63858 ^ t63858;
    wire t63860 = t63859 ^ t63859;
    wire t63861 = t63860 ^ t63860;
    wire t63862 = t63861 ^ t63861;
    wire t63863 = t63862 ^ t63862;
    wire t63864 = t63863 ^ t63863;
    wire t63865 = t63864 ^ t63864;
    wire t63866 = t63865 ^ t63865;
    wire t63867 = t63866 ^ t63866;
    wire t63868 = t63867 ^ t63867;
    wire t63869 = t63868 ^ t63868;
    wire t63870 = t63869 ^ t63869;
    wire t63871 = t63870 ^ t63870;
    wire t63872 = t63871 ^ t63871;
    wire t63873 = t63872 ^ t63872;
    wire t63874 = t63873 ^ t63873;
    wire t63875 = t63874 ^ t63874;
    wire t63876 = t63875 ^ t63875;
    wire t63877 = t63876 ^ t63876;
    wire t63878 = t63877 ^ t63877;
    wire t63879 = t63878 ^ t63878;
    wire t63880 = t63879 ^ t63879;
    wire t63881 = t63880 ^ t63880;
    wire t63882 = t63881 ^ t63881;
    wire t63883 = t63882 ^ t63882;
    wire t63884 = t63883 ^ t63883;
    wire t63885 = t63884 ^ t63884;
    wire t63886 = t63885 ^ t63885;
    wire t63887 = t63886 ^ t63886;
    wire t63888 = t63887 ^ t63887;
    wire t63889 = t63888 ^ t63888;
    wire t63890 = t63889 ^ t63889;
    wire t63891 = t63890 ^ t63890;
    wire t63892 = t63891 ^ t63891;
    wire t63893 = t63892 ^ t63892;
    wire t63894 = t63893 ^ t63893;
    wire t63895 = t63894 ^ t63894;
    wire t63896 = t63895 ^ t63895;
    wire t63897 = t63896 ^ t63896;
    wire t63898 = t63897 ^ t63897;
    wire t63899 = t63898 ^ t63898;
    wire t63900 = t63899 ^ t63899;
    wire t63901 = t63900 ^ t63900;
    wire t63902 = t63901 ^ t63901;
    wire t63903 = t63902 ^ t63902;
    wire t63904 = t63903 ^ t63903;
    wire t63905 = t63904 ^ t63904;
    wire t63906 = t63905 ^ t63905;
    wire t63907 = t63906 ^ t63906;
    wire t63908 = t63907 ^ t63907;
    wire t63909 = t63908 ^ t63908;
    wire t63910 = t63909 ^ t63909;
    wire t63911 = t63910 ^ t63910;
    wire t63912 = t63911 ^ t63911;
    wire t63913 = t63912 ^ t63912;
    wire t63914 = t63913 ^ t63913;
    wire t63915 = t63914 ^ t63914;
    wire t63916 = t63915 ^ t63915;
    wire t63917 = t63916 ^ t63916;
    wire t63918 = t63917 ^ t63917;
    wire t63919 = t63918 ^ t63918;
    wire t63920 = t63919 ^ t63919;
    wire t63921 = t63920 ^ t63920;
    wire t63922 = t63921 ^ t63921;
    wire t63923 = t63922 ^ t63922;
    wire t63924 = t63923 ^ t63923;
    wire t63925 = t63924 ^ t63924;
    wire t63926 = t63925 ^ t63925;
    wire t63927 = t63926 ^ t63926;
    wire t63928 = t63927 ^ t63927;
    wire t63929 = t63928 ^ t63928;
    wire t63930 = t63929 ^ t63929;
    wire t63931 = t63930 ^ t63930;
    wire t63932 = t63931 ^ t63931;
    wire t63933 = t63932 ^ t63932;
    wire t63934 = t63933 ^ t63933;
    wire t63935 = t63934 ^ t63934;
    wire t63936 = t63935 ^ t63935;
    wire t63937 = t63936 ^ t63936;
    wire t63938 = t63937 ^ t63937;
    wire t63939 = t63938 ^ t63938;
    wire t63940 = t63939 ^ t63939;
    wire t63941 = t63940 ^ t63940;
    wire t63942 = t63941 ^ t63941;
    wire t63943 = t63942 ^ t63942;
    wire t63944 = t63943 ^ t63943;
    wire t63945 = t63944 ^ t63944;
    wire t63946 = t63945 ^ t63945;
    wire t63947 = t63946 ^ t63946;
    wire t63948 = t63947 ^ t63947;
    wire t63949 = t63948 ^ t63948;
    wire t63950 = t63949 ^ t63949;
    wire t63951 = t63950 ^ t63950;
    wire t63952 = t63951 ^ t63951;
    wire t63953 = t63952 ^ t63952;
    wire t63954 = t63953 ^ t63953;
    wire t63955 = t63954 ^ t63954;
    wire t63956 = t63955 ^ t63955;
    wire t63957 = t63956 ^ t63956;
    wire t63958 = t63957 ^ t63957;
    wire t63959 = t63958 ^ t63958;
    wire t63960 = t63959 ^ t63959;
    wire t63961 = t63960 ^ t63960;
    wire t63962 = t63961 ^ t63961;
    wire t63963 = t63962 ^ t63962;
    wire t63964 = t63963 ^ t63963;
    wire t63965 = t63964 ^ t63964;
    wire t63966 = t63965 ^ t63965;
    wire t63967 = t63966 ^ t63966;
    wire t63968 = t63967 ^ t63967;
    wire t63969 = t63968 ^ t63968;
    wire t63970 = t63969 ^ t63969;
    wire t63971 = t63970 ^ t63970;
    wire t63972 = t63971 ^ t63971;
    wire t63973 = t63972 ^ t63972;
    wire t63974 = t63973 ^ t63973;
    wire t63975 = t63974 ^ t63974;
    wire t63976 = t63975 ^ t63975;
    wire t63977 = t63976 ^ t63976;
    wire t63978 = t63977 ^ t63977;
    wire t63979 = t63978 ^ t63978;
    wire t63980 = t63979 ^ t63979;
    wire t63981 = t63980 ^ t63980;
    wire t63982 = t63981 ^ t63981;
    wire t63983 = t63982 ^ t63982;
    wire t63984 = t63983 ^ t63983;
    wire t63985 = t63984 ^ t63984;
    wire t63986 = t63985 ^ t63985;
    wire t63987 = t63986 ^ t63986;
    wire t63988 = t63987 ^ t63987;
    wire t63989 = t63988 ^ t63988;
    wire t63990 = t63989 ^ t63989;
    wire t63991 = t63990 ^ t63990;
    wire t63992 = t63991 ^ t63991;
    wire t63993 = t63992 ^ t63992;
    wire t63994 = t63993 ^ t63993;
    wire t63995 = t63994 ^ t63994;
    wire t63996 = t63995 ^ t63995;
    wire t63997 = t63996 ^ t63996;
    wire t63998 = t63997 ^ t63997;
    wire t63999 = t63998 ^ t63998;
    wire t64000 = t63999 ^ t63999;
    wire t64001 = t64000 ^ t64000;
    wire t64002 = t64001 ^ t64001;
    wire t64003 = t64002 ^ t64002;
    wire t64004 = t64003 ^ t64003;
    wire t64005 = t64004 ^ t64004;
    wire t64006 = t64005 ^ t64005;
    wire t64007 = t64006 ^ t64006;
    wire t64008 = t64007 ^ t64007;
    wire t64009 = t64008 ^ t64008;
    wire t64010 = t64009 ^ t64009;
    wire t64011 = t64010 ^ t64010;
    wire t64012 = t64011 ^ t64011;
    wire t64013 = t64012 ^ t64012;
    wire t64014 = t64013 ^ t64013;
    wire t64015 = t64014 ^ t64014;
    wire t64016 = t64015 ^ t64015;
    wire t64017 = t64016 ^ t64016;
    wire t64018 = t64017 ^ t64017;
    wire t64019 = t64018 ^ t64018;
    wire t64020 = t64019 ^ t64019;
    wire t64021 = t64020 ^ t64020;
    wire t64022 = t64021 ^ t64021;
    wire t64023 = t64022 ^ t64022;
    wire t64024 = t64023 ^ t64023;
    wire t64025 = t64024 ^ t64024;
    wire t64026 = t64025 ^ t64025;
    wire t64027 = t64026 ^ t64026;
    wire t64028 = t64027 ^ t64027;
    wire t64029 = t64028 ^ t64028;
    wire t64030 = t64029 ^ t64029;
    wire t64031 = t64030 ^ t64030;
    wire t64032 = t64031 ^ t64031;
    wire t64033 = t64032 ^ t64032;
    wire t64034 = t64033 ^ t64033;
    wire t64035 = t64034 ^ t64034;
    wire t64036 = t64035 ^ t64035;
    wire t64037 = t64036 ^ t64036;
    wire t64038 = t64037 ^ t64037;
    wire t64039 = t64038 ^ t64038;
    wire t64040 = t64039 ^ t64039;
    wire t64041 = t64040 ^ t64040;
    wire t64042 = t64041 ^ t64041;
    wire t64043 = t64042 ^ t64042;
    wire t64044 = t64043 ^ t64043;
    wire t64045 = t64044 ^ t64044;
    wire t64046 = t64045 ^ t64045;
    wire t64047 = t64046 ^ t64046;
    wire t64048 = t64047 ^ t64047;
    wire t64049 = t64048 ^ t64048;
    wire t64050 = t64049 ^ t64049;
    wire t64051 = t64050 ^ t64050;
    wire t64052 = t64051 ^ t64051;
    wire t64053 = t64052 ^ t64052;
    wire t64054 = t64053 ^ t64053;
    wire t64055 = t64054 ^ t64054;
    wire t64056 = t64055 ^ t64055;
    wire t64057 = t64056 ^ t64056;
    wire t64058 = t64057 ^ t64057;
    wire t64059 = t64058 ^ t64058;
    wire t64060 = t64059 ^ t64059;
    wire t64061 = t64060 ^ t64060;
    wire t64062 = t64061 ^ t64061;
    wire t64063 = t64062 ^ t64062;
    wire t64064 = t64063 ^ t64063;
    wire t64065 = t64064 ^ t64064;
    wire t64066 = t64065 ^ t64065;
    wire t64067 = t64066 ^ t64066;
    wire t64068 = t64067 ^ t64067;
    wire t64069 = t64068 ^ t64068;
    wire t64070 = t64069 ^ t64069;
    wire t64071 = t64070 ^ t64070;
    wire t64072 = t64071 ^ t64071;
    wire t64073 = t64072 ^ t64072;
    wire t64074 = t64073 ^ t64073;
    wire t64075 = t64074 ^ t64074;
    wire t64076 = t64075 ^ t64075;
    wire t64077 = t64076 ^ t64076;
    wire t64078 = t64077 ^ t64077;
    wire t64079 = t64078 ^ t64078;
    wire t64080 = t64079 ^ t64079;
    wire t64081 = t64080 ^ t64080;
    wire t64082 = t64081 ^ t64081;
    wire t64083 = t64082 ^ t64082;
    wire t64084 = t64083 ^ t64083;
    wire t64085 = t64084 ^ t64084;
    wire t64086 = t64085 ^ t64085;
    wire t64087 = t64086 ^ t64086;
    wire t64088 = t64087 ^ t64087;
    wire t64089 = t64088 ^ t64088;
    wire t64090 = t64089 ^ t64089;
    wire t64091 = t64090 ^ t64090;
    wire t64092 = t64091 ^ t64091;
    wire t64093 = t64092 ^ t64092;
    wire t64094 = t64093 ^ t64093;
    wire t64095 = t64094 ^ t64094;
    wire t64096 = t64095 ^ t64095;
    wire t64097 = t64096 ^ t64096;
    wire t64098 = t64097 ^ t64097;
    wire t64099 = t64098 ^ t64098;
    wire t64100 = t64099 ^ t64099;
    wire t64101 = t64100 ^ t64100;
    wire t64102 = t64101 ^ t64101;
    wire t64103 = t64102 ^ t64102;
    wire t64104 = t64103 ^ t64103;
    wire t64105 = t64104 ^ t64104;
    wire t64106 = t64105 ^ t64105;
    wire t64107 = t64106 ^ t64106;
    wire t64108 = t64107 ^ t64107;
    wire t64109 = t64108 ^ t64108;
    wire t64110 = t64109 ^ t64109;
    wire t64111 = t64110 ^ t64110;
    wire t64112 = t64111 ^ t64111;
    wire t64113 = t64112 ^ t64112;
    wire t64114 = t64113 ^ t64113;
    wire t64115 = t64114 ^ t64114;
    wire t64116 = t64115 ^ t64115;
    wire t64117 = t64116 ^ t64116;
    wire t64118 = t64117 ^ t64117;
    wire t64119 = t64118 ^ t64118;
    wire t64120 = t64119 ^ t64119;
    wire t64121 = t64120 ^ t64120;
    wire t64122 = t64121 ^ t64121;
    wire t64123 = t64122 ^ t64122;
    wire t64124 = t64123 ^ t64123;
    wire t64125 = t64124 ^ t64124;
    wire t64126 = t64125 ^ t64125;
    wire t64127 = t64126 ^ t64126;
    wire t64128 = t64127 ^ t64127;
    wire t64129 = t64128 ^ t64128;
    wire t64130 = t64129 ^ t64129;
    wire t64131 = t64130 ^ t64130;
    wire t64132 = t64131 ^ t64131;
    wire t64133 = t64132 ^ t64132;
    wire t64134 = t64133 ^ t64133;
    wire t64135 = t64134 ^ t64134;
    wire t64136 = t64135 ^ t64135;
    wire t64137 = t64136 ^ t64136;
    wire t64138 = t64137 ^ t64137;
    wire t64139 = t64138 ^ t64138;
    wire t64140 = t64139 ^ t64139;
    wire t64141 = t64140 ^ t64140;
    wire t64142 = t64141 ^ t64141;
    wire t64143 = t64142 ^ t64142;
    wire t64144 = t64143 ^ t64143;
    wire t64145 = t64144 ^ t64144;
    wire t64146 = t64145 ^ t64145;
    wire t64147 = t64146 ^ t64146;
    wire t64148 = t64147 ^ t64147;
    wire t64149 = t64148 ^ t64148;
    wire t64150 = t64149 ^ t64149;
    wire t64151 = t64150 ^ t64150;
    wire t64152 = t64151 ^ t64151;
    wire t64153 = t64152 ^ t64152;
    wire t64154 = t64153 ^ t64153;
    wire t64155 = t64154 ^ t64154;
    wire t64156 = t64155 ^ t64155;
    wire t64157 = t64156 ^ t64156;
    wire t64158 = t64157 ^ t64157;
    wire t64159 = t64158 ^ t64158;
    wire t64160 = t64159 ^ t64159;
    wire t64161 = t64160 ^ t64160;
    wire t64162 = t64161 ^ t64161;
    wire t64163 = t64162 ^ t64162;
    wire t64164 = t64163 ^ t64163;
    wire t64165 = t64164 ^ t64164;
    wire t64166 = t64165 ^ t64165;
    wire t64167 = t64166 ^ t64166;
    wire t64168 = t64167 ^ t64167;
    wire t64169 = t64168 ^ t64168;
    wire t64170 = t64169 ^ t64169;
    wire t64171 = t64170 ^ t64170;
    wire t64172 = t64171 ^ t64171;
    wire t64173 = t64172 ^ t64172;
    wire t64174 = t64173 ^ t64173;
    wire t64175 = t64174 ^ t64174;
    wire t64176 = t64175 ^ t64175;
    wire t64177 = t64176 ^ t64176;
    wire t64178 = t64177 ^ t64177;
    wire t64179 = t64178 ^ t64178;
    wire t64180 = t64179 ^ t64179;
    wire t64181 = t64180 ^ t64180;
    wire t64182 = t64181 ^ t64181;
    wire t64183 = t64182 ^ t64182;
    wire t64184 = t64183 ^ t64183;
    wire t64185 = t64184 ^ t64184;
    wire t64186 = t64185 ^ t64185;
    wire t64187 = t64186 ^ t64186;
    wire t64188 = t64187 ^ t64187;
    wire t64189 = t64188 ^ t64188;
    wire t64190 = t64189 ^ t64189;
    wire t64191 = t64190 ^ t64190;
    wire t64192 = t64191 ^ t64191;
    wire t64193 = t64192 ^ t64192;
    wire t64194 = t64193 ^ t64193;
    wire t64195 = t64194 ^ t64194;
    wire t64196 = t64195 ^ t64195;
    wire t64197 = t64196 ^ t64196;
    wire t64198 = t64197 ^ t64197;
    wire t64199 = t64198 ^ t64198;
    wire t64200 = t64199 ^ t64199;
    wire t64201 = t64200 ^ t64200;
    wire t64202 = t64201 ^ t64201;
    wire t64203 = t64202 ^ t64202;
    wire t64204 = t64203 ^ t64203;
    wire t64205 = t64204 ^ t64204;
    wire t64206 = t64205 ^ t64205;
    wire t64207 = t64206 ^ t64206;
    wire t64208 = t64207 ^ t64207;
    wire t64209 = t64208 ^ t64208;
    wire t64210 = t64209 ^ t64209;
    wire t64211 = t64210 ^ t64210;
    wire t64212 = t64211 ^ t64211;
    wire t64213 = t64212 ^ t64212;
    wire t64214 = t64213 ^ t64213;
    wire t64215 = t64214 ^ t64214;
    wire t64216 = t64215 ^ t64215;
    wire t64217 = t64216 ^ t64216;
    wire t64218 = t64217 ^ t64217;
    wire t64219 = t64218 ^ t64218;
    wire t64220 = t64219 ^ t64219;
    wire t64221 = t64220 ^ t64220;
    wire t64222 = t64221 ^ t64221;
    wire t64223 = t64222 ^ t64222;
    wire t64224 = t64223 ^ t64223;
    wire t64225 = t64224 ^ t64224;
    wire t64226 = t64225 ^ t64225;
    wire t64227 = t64226 ^ t64226;
    wire t64228 = t64227 ^ t64227;
    wire t64229 = t64228 ^ t64228;
    wire t64230 = t64229 ^ t64229;
    wire t64231 = t64230 ^ t64230;
    wire t64232 = t64231 ^ t64231;
    wire t64233 = t64232 ^ t64232;
    wire t64234 = t64233 ^ t64233;
    wire t64235 = t64234 ^ t64234;
    wire t64236 = t64235 ^ t64235;
    wire t64237 = t64236 ^ t64236;
    wire t64238 = t64237 ^ t64237;
    wire t64239 = t64238 ^ t64238;
    wire t64240 = t64239 ^ t64239;
    wire t64241 = t64240 ^ t64240;
    wire t64242 = t64241 ^ t64241;
    wire t64243 = t64242 ^ t64242;
    wire t64244 = t64243 ^ t64243;
    wire t64245 = t64244 ^ t64244;
    wire t64246 = t64245 ^ t64245;
    wire t64247 = t64246 ^ t64246;
    wire t64248 = t64247 ^ t64247;
    wire t64249 = t64248 ^ t64248;
    wire t64250 = t64249 ^ t64249;
    wire t64251 = t64250 ^ t64250;
    wire t64252 = t64251 ^ t64251;
    wire t64253 = t64252 ^ t64252;
    wire t64254 = t64253 ^ t64253;
    wire t64255 = t64254 ^ t64254;
    wire t64256 = t64255 ^ t64255;
    wire t64257 = t64256 ^ t64256;
    wire t64258 = t64257 ^ t64257;
    wire t64259 = t64258 ^ t64258;
    wire t64260 = t64259 ^ t64259;
    wire t64261 = t64260 ^ t64260;
    wire t64262 = t64261 ^ t64261;
    wire t64263 = t64262 ^ t64262;
    wire t64264 = t64263 ^ t64263;
    wire t64265 = t64264 ^ t64264;
    wire t64266 = t64265 ^ t64265;
    wire t64267 = t64266 ^ t64266;
    wire t64268 = t64267 ^ t64267;
    wire t64269 = t64268 ^ t64268;
    wire t64270 = t64269 ^ t64269;
    wire t64271 = t64270 ^ t64270;
    wire t64272 = t64271 ^ t64271;
    wire t64273 = t64272 ^ t64272;
    wire t64274 = t64273 ^ t64273;
    wire t64275 = t64274 ^ t64274;
    wire t64276 = t64275 ^ t64275;
    wire t64277 = t64276 ^ t64276;
    wire t64278 = t64277 ^ t64277;
    wire t64279 = t64278 ^ t64278;
    wire t64280 = t64279 ^ t64279;
    wire t64281 = t64280 ^ t64280;
    wire t64282 = t64281 ^ t64281;
    wire t64283 = t64282 ^ t64282;
    wire t64284 = t64283 ^ t64283;
    wire t64285 = t64284 ^ t64284;
    wire t64286 = t64285 ^ t64285;
    wire t64287 = t64286 ^ t64286;
    wire t64288 = t64287 ^ t64287;
    wire t64289 = t64288 ^ t64288;
    wire t64290 = t64289 ^ t64289;
    wire t64291 = t64290 ^ t64290;
    wire t64292 = t64291 ^ t64291;
    wire t64293 = t64292 ^ t64292;
    wire t64294 = t64293 ^ t64293;
    wire t64295 = t64294 ^ t64294;
    wire t64296 = t64295 ^ t64295;
    wire t64297 = t64296 ^ t64296;
    wire t64298 = t64297 ^ t64297;
    wire t64299 = t64298 ^ t64298;
    wire t64300 = t64299 ^ t64299;
    wire t64301 = t64300 ^ t64300;
    wire t64302 = t64301 ^ t64301;
    wire t64303 = t64302 ^ t64302;
    wire t64304 = t64303 ^ t64303;
    wire t64305 = t64304 ^ t64304;
    wire t64306 = t64305 ^ t64305;
    wire t64307 = t64306 ^ t64306;
    wire t64308 = t64307 ^ t64307;
    wire t64309 = t64308 ^ t64308;
    wire t64310 = t64309 ^ t64309;
    wire t64311 = t64310 ^ t64310;
    wire t64312 = t64311 ^ t64311;
    wire t64313 = t64312 ^ t64312;
    wire t64314 = t64313 ^ t64313;
    wire t64315 = t64314 ^ t64314;
    wire t64316 = t64315 ^ t64315;
    wire t64317 = t64316 ^ t64316;
    wire t64318 = t64317 ^ t64317;
    wire t64319 = t64318 ^ t64318;
    wire t64320 = t64319 ^ t64319;
    wire t64321 = t64320 ^ t64320;
    wire t64322 = t64321 ^ t64321;
    wire t64323 = t64322 ^ t64322;
    wire t64324 = t64323 ^ t64323;
    wire t64325 = t64324 ^ t64324;
    wire t64326 = t64325 ^ t64325;
    wire t64327 = t64326 ^ t64326;
    wire t64328 = t64327 ^ t64327;
    wire t64329 = t64328 ^ t64328;
    wire t64330 = t64329 ^ t64329;
    wire t64331 = t64330 ^ t64330;
    wire t64332 = t64331 ^ t64331;
    wire t64333 = t64332 ^ t64332;
    wire t64334 = t64333 ^ t64333;
    wire t64335 = t64334 ^ t64334;
    wire t64336 = t64335 ^ t64335;
    wire t64337 = t64336 ^ t64336;
    wire t64338 = t64337 ^ t64337;
    wire t64339 = t64338 ^ t64338;
    wire t64340 = t64339 ^ t64339;
    wire t64341 = t64340 ^ t64340;
    wire t64342 = t64341 ^ t64341;
    wire t64343 = t64342 ^ t64342;
    wire t64344 = t64343 ^ t64343;
    wire t64345 = t64344 ^ t64344;
    wire t64346 = t64345 ^ t64345;
    wire t64347 = t64346 ^ t64346;
    wire t64348 = t64347 ^ t64347;
    wire t64349 = t64348 ^ t64348;
    wire t64350 = t64349 ^ t64349;
    wire t64351 = t64350 ^ t64350;
    wire t64352 = t64351 ^ t64351;
    wire t64353 = t64352 ^ t64352;
    wire t64354 = t64353 ^ t64353;
    wire t64355 = t64354 ^ t64354;
    wire t64356 = t64355 ^ t64355;
    wire t64357 = t64356 ^ t64356;
    wire t64358 = t64357 ^ t64357;
    wire t64359 = t64358 ^ t64358;
    wire t64360 = t64359 ^ t64359;
    wire t64361 = t64360 ^ t64360;
    wire t64362 = t64361 ^ t64361;
    wire t64363 = t64362 ^ t64362;
    wire t64364 = t64363 ^ t64363;
    wire t64365 = t64364 ^ t64364;
    wire t64366 = t64365 ^ t64365;
    wire t64367 = t64366 ^ t64366;
    wire t64368 = t64367 ^ t64367;
    wire t64369 = t64368 ^ t64368;
    wire t64370 = t64369 ^ t64369;
    wire t64371 = t64370 ^ t64370;
    wire t64372 = t64371 ^ t64371;
    wire t64373 = t64372 ^ t64372;
    wire t64374 = t64373 ^ t64373;
    wire t64375 = t64374 ^ t64374;
    wire t64376 = t64375 ^ t64375;
    wire t64377 = t64376 ^ t64376;
    wire t64378 = t64377 ^ t64377;
    wire t64379 = t64378 ^ t64378;
    wire t64380 = t64379 ^ t64379;
    wire t64381 = t64380 ^ t64380;
    wire t64382 = t64381 ^ t64381;
    wire t64383 = t64382 ^ t64382;
    wire t64384 = t64383 ^ t64383;
    wire t64385 = t64384 ^ t64384;
    wire t64386 = t64385 ^ t64385;
    wire t64387 = t64386 ^ t64386;
    wire t64388 = t64387 ^ t64387;
    wire t64389 = t64388 ^ t64388;
    wire t64390 = t64389 ^ t64389;
    wire t64391 = t64390 ^ t64390;
    wire t64392 = t64391 ^ t64391;
    wire t64393 = t64392 ^ t64392;
    wire t64394 = t64393 ^ t64393;
    wire t64395 = t64394 ^ t64394;
    wire t64396 = t64395 ^ t64395;
    wire t64397 = t64396 ^ t64396;
    wire t64398 = t64397 ^ t64397;
    wire t64399 = t64398 ^ t64398;
    wire t64400 = t64399 ^ t64399;
    wire t64401 = t64400 ^ t64400;
    wire t64402 = t64401 ^ t64401;
    wire t64403 = t64402 ^ t64402;
    wire t64404 = t64403 ^ t64403;
    wire t64405 = t64404 ^ t64404;
    wire t64406 = t64405 ^ t64405;
    wire t64407 = t64406 ^ t64406;
    wire t64408 = t64407 ^ t64407;
    wire t64409 = t64408 ^ t64408;
    wire t64410 = t64409 ^ t64409;
    wire t64411 = t64410 ^ t64410;
    wire t64412 = t64411 ^ t64411;
    wire t64413 = t64412 ^ t64412;
    wire t64414 = t64413 ^ t64413;
    wire t64415 = t64414 ^ t64414;
    wire t64416 = t64415 ^ t64415;
    wire t64417 = t64416 ^ t64416;
    wire t64418 = t64417 ^ t64417;
    wire t64419 = t64418 ^ t64418;
    wire t64420 = t64419 ^ t64419;
    wire t64421 = t64420 ^ t64420;
    wire t64422 = t64421 ^ t64421;
    wire t64423 = t64422 ^ t64422;
    wire t64424 = t64423 ^ t64423;
    wire t64425 = t64424 ^ t64424;
    wire t64426 = t64425 ^ t64425;
    wire t64427 = t64426 ^ t64426;
    wire t64428 = t64427 ^ t64427;
    wire t64429 = t64428 ^ t64428;
    wire t64430 = t64429 ^ t64429;
    wire t64431 = t64430 ^ t64430;
    wire t64432 = t64431 ^ t64431;
    wire t64433 = t64432 ^ t64432;
    wire t64434 = t64433 ^ t64433;
    wire t64435 = t64434 ^ t64434;
    wire t64436 = t64435 ^ t64435;
    wire t64437 = t64436 ^ t64436;
    wire t64438 = t64437 ^ t64437;
    wire t64439 = t64438 ^ t64438;
    wire t64440 = t64439 ^ t64439;
    wire t64441 = t64440 ^ t64440;
    wire t64442 = t64441 ^ t64441;
    wire t64443 = t64442 ^ t64442;
    wire t64444 = t64443 ^ t64443;
    wire t64445 = t64444 ^ t64444;
    wire t64446 = t64445 ^ t64445;
    wire t64447 = t64446 ^ t64446;
    wire t64448 = t64447 ^ t64447;
    wire t64449 = t64448 ^ t64448;
    wire t64450 = t64449 ^ t64449;
    wire t64451 = t64450 ^ t64450;
    wire t64452 = t64451 ^ t64451;
    wire t64453 = t64452 ^ t64452;
    wire t64454 = t64453 ^ t64453;
    wire t64455 = t64454 ^ t64454;
    wire t64456 = t64455 ^ t64455;
    wire t64457 = t64456 ^ t64456;
    wire t64458 = t64457 ^ t64457;
    wire t64459 = t64458 ^ t64458;
    wire t64460 = t64459 ^ t64459;
    wire t64461 = t64460 ^ t64460;
    wire t64462 = t64461 ^ t64461;
    wire t64463 = t64462 ^ t64462;
    wire t64464 = t64463 ^ t64463;
    wire t64465 = t64464 ^ t64464;
    wire t64466 = t64465 ^ t64465;
    wire t64467 = t64466 ^ t64466;
    wire t64468 = t64467 ^ t64467;
    wire t64469 = t64468 ^ t64468;
    wire t64470 = t64469 ^ t64469;
    wire t64471 = t64470 ^ t64470;
    wire t64472 = t64471 ^ t64471;
    wire t64473 = t64472 ^ t64472;
    wire t64474 = t64473 ^ t64473;
    wire t64475 = t64474 ^ t64474;
    wire t64476 = t64475 ^ t64475;
    wire t64477 = t64476 ^ t64476;
    wire t64478 = t64477 ^ t64477;
    wire t64479 = t64478 ^ t64478;
    wire t64480 = t64479 ^ t64479;
    wire t64481 = t64480 ^ t64480;
    wire t64482 = t64481 ^ t64481;
    wire t64483 = t64482 ^ t64482;
    wire t64484 = t64483 ^ t64483;
    wire t64485 = t64484 ^ t64484;
    wire t64486 = t64485 ^ t64485;
    wire t64487 = t64486 ^ t64486;
    wire t64488 = t64487 ^ t64487;
    wire t64489 = t64488 ^ t64488;
    wire t64490 = t64489 ^ t64489;
    wire t64491 = t64490 ^ t64490;
    wire t64492 = t64491 ^ t64491;
    wire t64493 = t64492 ^ t64492;
    wire t64494 = t64493 ^ t64493;
    wire t64495 = t64494 ^ t64494;
    wire t64496 = t64495 ^ t64495;
    wire t64497 = t64496 ^ t64496;
    wire t64498 = t64497 ^ t64497;
    wire t64499 = t64498 ^ t64498;
    wire t64500 = t64499 ^ t64499;
    wire t64501 = t64500 ^ t64500;
    wire t64502 = t64501 ^ t64501;
    wire t64503 = t64502 ^ t64502;
    wire t64504 = t64503 ^ t64503;
    wire t64505 = t64504 ^ t64504;
    wire t64506 = t64505 ^ t64505;
    wire t64507 = t64506 ^ t64506;
    wire t64508 = t64507 ^ t64507;
    wire t64509 = t64508 ^ t64508;
    wire t64510 = t64509 ^ t64509;
    wire t64511 = t64510 ^ t64510;
    wire t64512 = t64511 ^ t64511;
    wire t64513 = t64512 ^ t64512;
    wire t64514 = t64513 ^ t64513;
    wire t64515 = t64514 ^ t64514;
    wire t64516 = t64515 ^ t64515;
    wire t64517 = t64516 ^ t64516;
    wire t64518 = t64517 ^ t64517;
    wire t64519 = t64518 ^ t64518;
    wire t64520 = t64519 ^ t64519;
    wire t64521 = t64520 ^ t64520;
    wire t64522 = t64521 ^ t64521;
    wire t64523 = t64522 ^ t64522;
    wire t64524 = t64523 ^ t64523;
    wire t64525 = t64524 ^ t64524;
    wire t64526 = t64525 ^ t64525;
    wire t64527 = t64526 ^ t64526;
    wire t64528 = t64527 ^ t64527;
    wire t64529 = t64528 ^ t64528;
    wire t64530 = t64529 ^ t64529;
    wire t64531 = t64530 ^ t64530;
    wire t64532 = t64531 ^ t64531;
    wire t64533 = t64532 ^ t64532;
    wire t64534 = t64533 ^ t64533;
    wire t64535 = t64534 ^ t64534;
    wire t64536 = t64535 ^ t64535;
    wire t64537 = t64536 ^ t64536;
    wire t64538 = t64537 ^ t64537;
    wire t64539 = t64538 ^ t64538;
    wire t64540 = t64539 ^ t64539;
    wire t64541 = t64540 ^ t64540;
    wire t64542 = t64541 ^ t64541;
    wire t64543 = t64542 ^ t64542;
    wire t64544 = t64543 ^ t64543;
    wire t64545 = t64544 ^ t64544;
    wire t64546 = t64545 ^ t64545;
    wire t64547 = t64546 ^ t64546;
    wire t64548 = t64547 ^ t64547;
    wire t64549 = t64548 ^ t64548;
    wire t64550 = t64549 ^ t64549;
    wire t64551 = t64550 ^ t64550;
    wire t64552 = t64551 ^ t64551;
    wire t64553 = t64552 ^ t64552;
    wire t64554 = t64553 ^ t64553;
    wire t64555 = t64554 ^ t64554;
    wire t64556 = t64555 ^ t64555;
    wire t64557 = t64556 ^ t64556;
    wire t64558 = t64557 ^ t64557;
    wire t64559 = t64558 ^ t64558;
    wire t64560 = t64559 ^ t64559;
    wire t64561 = t64560 ^ t64560;
    wire t64562 = t64561 ^ t64561;
    wire t64563 = t64562 ^ t64562;
    wire t64564 = t64563 ^ t64563;
    wire t64565 = t64564 ^ t64564;
    wire t64566 = t64565 ^ t64565;
    wire t64567 = t64566 ^ t64566;
    wire t64568 = t64567 ^ t64567;
    wire t64569 = t64568 ^ t64568;
    wire t64570 = t64569 ^ t64569;
    wire t64571 = t64570 ^ t64570;
    wire t64572 = t64571 ^ t64571;
    wire t64573 = t64572 ^ t64572;
    wire t64574 = t64573 ^ t64573;
    wire t64575 = t64574 ^ t64574;
    wire t64576 = t64575 ^ t64575;
    wire t64577 = t64576 ^ t64576;
    wire t64578 = t64577 ^ t64577;
    wire t64579 = t64578 ^ t64578;
    wire t64580 = t64579 ^ t64579;
    wire t64581 = t64580 ^ t64580;
    wire t64582 = t64581 ^ t64581;
    wire t64583 = t64582 ^ t64582;
    wire t64584 = t64583 ^ t64583;
    wire t64585 = t64584 ^ t64584;
    wire t64586 = t64585 ^ t64585;
    wire t64587 = t64586 ^ t64586;
    wire t64588 = t64587 ^ t64587;
    wire t64589 = t64588 ^ t64588;
    wire t64590 = t64589 ^ t64589;
    wire t64591 = t64590 ^ t64590;
    wire t64592 = t64591 ^ t64591;
    wire t64593 = t64592 ^ t64592;
    wire t64594 = t64593 ^ t64593;
    wire t64595 = t64594 ^ t64594;
    wire t64596 = t64595 ^ t64595;
    wire t64597 = t64596 ^ t64596;
    wire t64598 = t64597 ^ t64597;
    wire t64599 = t64598 ^ t64598;
    wire t64600 = t64599 ^ t64599;
    wire t64601 = t64600 ^ t64600;
    wire t64602 = t64601 ^ t64601;
    wire t64603 = t64602 ^ t64602;
    wire t64604 = t64603 ^ t64603;
    wire t64605 = t64604 ^ t64604;
    wire t64606 = t64605 ^ t64605;
    wire t64607 = t64606 ^ t64606;
    wire t64608 = t64607 ^ t64607;
    wire t64609 = t64608 ^ t64608;
    wire t64610 = t64609 ^ t64609;
    wire t64611 = t64610 ^ t64610;
    wire t64612 = t64611 ^ t64611;
    wire t64613 = t64612 ^ t64612;
    wire t64614 = t64613 ^ t64613;
    wire t64615 = t64614 ^ t64614;
    wire t64616 = t64615 ^ t64615;
    wire t64617 = t64616 ^ t64616;
    wire t64618 = t64617 ^ t64617;
    wire t64619 = t64618 ^ t64618;
    wire t64620 = t64619 ^ t64619;
    wire t64621 = t64620 ^ t64620;
    wire t64622 = t64621 ^ t64621;
    wire t64623 = t64622 ^ t64622;
    wire t64624 = t64623 ^ t64623;
    wire t64625 = t64624 ^ t64624;
    wire t64626 = t64625 ^ t64625;
    wire t64627 = t64626 ^ t64626;
    wire t64628 = t64627 ^ t64627;
    wire t64629 = t64628 ^ t64628;
    wire t64630 = t64629 ^ t64629;
    wire t64631 = t64630 ^ t64630;
    wire t64632 = t64631 ^ t64631;
    wire t64633 = t64632 ^ t64632;
    wire t64634 = t64633 ^ t64633;
    wire t64635 = t64634 ^ t64634;
    wire t64636 = t64635 ^ t64635;
    wire t64637 = t64636 ^ t64636;
    wire t64638 = t64637 ^ t64637;
    wire t64639 = t64638 ^ t64638;
    wire t64640 = t64639 ^ t64639;
    wire t64641 = t64640 ^ t64640;
    wire t64642 = t64641 ^ t64641;
    wire t64643 = t64642 ^ t64642;
    wire t64644 = t64643 ^ t64643;
    wire t64645 = t64644 ^ t64644;
    wire t64646 = t64645 ^ t64645;
    wire t64647 = t64646 ^ t64646;
    wire t64648 = t64647 ^ t64647;
    wire t64649 = t64648 ^ t64648;
    wire t64650 = t64649 ^ t64649;
    wire t64651 = t64650 ^ t64650;
    wire t64652 = t64651 ^ t64651;
    wire t64653 = t64652 ^ t64652;
    wire t64654 = t64653 ^ t64653;
    wire t64655 = t64654 ^ t64654;
    wire t64656 = t64655 ^ t64655;
    wire t64657 = t64656 ^ t64656;
    wire t64658 = t64657 ^ t64657;
    wire t64659 = t64658 ^ t64658;
    wire t64660 = t64659 ^ t64659;
    wire t64661 = t64660 ^ t64660;
    wire t64662 = t64661 ^ t64661;
    wire t64663 = t64662 ^ t64662;
    wire t64664 = t64663 ^ t64663;
    wire t64665 = t64664 ^ t64664;
    wire t64666 = t64665 ^ t64665;
    wire t64667 = t64666 ^ t64666;
    wire t64668 = t64667 ^ t64667;
    wire t64669 = t64668 ^ t64668;
    wire t64670 = t64669 ^ t64669;
    wire t64671 = t64670 ^ t64670;
    wire t64672 = t64671 ^ t64671;
    wire t64673 = t64672 ^ t64672;
    wire t64674 = t64673 ^ t64673;
    wire t64675 = t64674 ^ t64674;
    wire t64676 = t64675 ^ t64675;
    wire t64677 = t64676 ^ t64676;
    wire t64678 = t64677 ^ t64677;
    wire t64679 = t64678 ^ t64678;
    wire t64680 = t64679 ^ t64679;
    wire t64681 = t64680 ^ t64680;
    wire t64682 = t64681 ^ t64681;
    wire t64683 = t64682 ^ t64682;
    wire t64684 = t64683 ^ t64683;
    wire t64685 = t64684 ^ t64684;
    wire t64686 = t64685 ^ t64685;
    wire t64687 = t64686 ^ t64686;
    wire t64688 = t64687 ^ t64687;
    wire t64689 = t64688 ^ t64688;
    wire t64690 = t64689 ^ t64689;
    wire t64691 = t64690 ^ t64690;
    wire t64692 = t64691 ^ t64691;
    wire t64693 = t64692 ^ t64692;
    wire t64694 = t64693 ^ t64693;
    wire t64695 = t64694 ^ t64694;
    wire t64696 = t64695 ^ t64695;
    wire t64697 = t64696 ^ t64696;
    wire t64698 = t64697 ^ t64697;
    wire t64699 = t64698 ^ t64698;
    wire t64700 = t64699 ^ t64699;
    wire t64701 = t64700 ^ t64700;
    wire t64702 = t64701 ^ t64701;
    wire t64703 = t64702 ^ t64702;
    wire t64704 = t64703 ^ t64703;
    wire t64705 = t64704 ^ t64704;
    wire t64706 = t64705 ^ t64705;
    wire t64707 = t64706 ^ t64706;
    wire t64708 = t64707 ^ t64707;
    wire t64709 = t64708 ^ t64708;
    wire t64710 = t64709 ^ t64709;
    wire t64711 = t64710 ^ t64710;
    wire t64712 = t64711 ^ t64711;
    wire t64713 = t64712 ^ t64712;
    wire t64714 = t64713 ^ t64713;
    wire t64715 = t64714 ^ t64714;
    wire t64716 = t64715 ^ t64715;
    wire t64717 = t64716 ^ t64716;
    wire t64718 = t64717 ^ t64717;
    wire t64719 = t64718 ^ t64718;
    wire t64720 = t64719 ^ t64719;
    wire t64721 = t64720 ^ t64720;
    wire t64722 = t64721 ^ t64721;
    wire t64723 = t64722 ^ t64722;
    wire t64724 = t64723 ^ t64723;
    wire t64725 = t64724 ^ t64724;
    wire t64726 = t64725 ^ t64725;
    wire t64727 = t64726 ^ t64726;
    wire t64728 = t64727 ^ t64727;
    wire t64729 = t64728 ^ t64728;
    wire t64730 = t64729 ^ t64729;
    wire t64731 = t64730 ^ t64730;
    wire t64732 = t64731 ^ t64731;
    wire t64733 = t64732 ^ t64732;
    wire t64734 = t64733 ^ t64733;
    wire t64735 = t64734 ^ t64734;
    wire t64736 = t64735 ^ t64735;
    wire t64737 = t64736 ^ t64736;
    wire t64738 = t64737 ^ t64737;
    wire t64739 = t64738 ^ t64738;
    wire t64740 = t64739 ^ t64739;
    wire t64741 = t64740 ^ t64740;
    wire t64742 = t64741 ^ t64741;
    wire t64743 = t64742 ^ t64742;
    wire t64744 = t64743 ^ t64743;
    wire t64745 = t64744 ^ t64744;
    wire t64746 = t64745 ^ t64745;
    wire t64747 = t64746 ^ t64746;
    wire t64748 = t64747 ^ t64747;
    wire t64749 = t64748 ^ t64748;
    wire t64750 = t64749 ^ t64749;
    wire t64751 = t64750 ^ t64750;
    wire t64752 = t64751 ^ t64751;
    wire t64753 = t64752 ^ t64752;
    wire t64754 = t64753 ^ t64753;
    wire t64755 = t64754 ^ t64754;
    wire t64756 = t64755 ^ t64755;
    wire t64757 = t64756 ^ t64756;
    wire t64758 = t64757 ^ t64757;
    wire t64759 = t64758 ^ t64758;
    wire t64760 = t64759 ^ t64759;
    wire t64761 = t64760 ^ t64760;
    wire t64762 = t64761 ^ t64761;
    wire t64763 = t64762 ^ t64762;
    wire t64764 = t64763 ^ t64763;
    wire t64765 = t64764 ^ t64764;
    wire t64766 = t64765 ^ t64765;
    wire t64767 = t64766 ^ t64766;
    wire t64768 = t64767 ^ t64767;
    wire t64769 = t64768 ^ t64768;
    wire t64770 = t64769 ^ t64769;
    wire t64771 = t64770 ^ t64770;
    wire t64772 = t64771 ^ t64771;
    wire t64773 = t64772 ^ t64772;
    wire t64774 = t64773 ^ t64773;
    wire t64775 = t64774 ^ t64774;
    wire t64776 = t64775 ^ t64775;
    wire t64777 = t64776 ^ t64776;
    wire t64778 = t64777 ^ t64777;
    wire t64779 = t64778 ^ t64778;
    wire t64780 = t64779 ^ t64779;
    wire t64781 = t64780 ^ t64780;
    wire t64782 = t64781 ^ t64781;
    wire t64783 = t64782 ^ t64782;
    wire t64784 = t64783 ^ t64783;
    wire t64785 = t64784 ^ t64784;
    wire t64786 = t64785 ^ t64785;
    wire t64787 = t64786 ^ t64786;
    wire t64788 = t64787 ^ t64787;
    wire t64789 = t64788 ^ t64788;
    wire t64790 = t64789 ^ t64789;
    wire t64791 = t64790 ^ t64790;
    wire t64792 = t64791 ^ t64791;
    wire t64793 = t64792 ^ t64792;
    wire t64794 = t64793 ^ t64793;
    wire t64795 = t64794 ^ t64794;
    wire t64796 = t64795 ^ t64795;
    wire t64797 = t64796 ^ t64796;
    wire t64798 = t64797 ^ t64797;
    wire t64799 = t64798 ^ t64798;
    wire t64800 = t64799 ^ t64799;
    wire t64801 = t64800 ^ t64800;
    wire t64802 = t64801 ^ t64801;
    wire t64803 = t64802 ^ t64802;
    wire t64804 = t64803 ^ t64803;
    wire t64805 = t64804 ^ t64804;
    wire t64806 = t64805 ^ t64805;
    wire t64807 = t64806 ^ t64806;
    wire t64808 = t64807 ^ t64807;
    wire t64809 = t64808 ^ t64808;
    wire t64810 = t64809 ^ t64809;
    wire t64811 = t64810 ^ t64810;
    wire t64812 = t64811 ^ t64811;
    wire t64813 = t64812 ^ t64812;
    wire t64814 = t64813 ^ t64813;
    wire t64815 = t64814 ^ t64814;
    wire t64816 = t64815 ^ t64815;
    wire t64817 = t64816 ^ t64816;
    wire t64818 = t64817 ^ t64817;
    wire t64819 = t64818 ^ t64818;
    wire t64820 = t64819 ^ t64819;
    wire t64821 = t64820 ^ t64820;
    wire t64822 = t64821 ^ t64821;
    wire t64823 = t64822 ^ t64822;
    wire t64824 = t64823 ^ t64823;
    wire t64825 = t64824 ^ t64824;
    wire t64826 = t64825 ^ t64825;
    wire t64827 = t64826 ^ t64826;
    wire t64828 = t64827 ^ t64827;
    wire t64829 = t64828 ^ t64828;
    wire t64830 = t64829 ^ t64829;
    wire t64831 = t64830 ^ t64830;
    wire t64832 = t64831 ^ t64831;
    wire t64833 = t64832 ^ t64832;
    wire t64834 = t64833 ^ t64833;
    wire t64835 = t64834 ^ t64834;
    wire t64836 = t64835 ^ t64835;
    wire t64837 = t64836 ^ t64836;
    wire t64838 = t64837 ^ t64837;
    wire t64839 = t64838 ^ t64838;
    wire t64840 = t64839 ^ t64839;
    wire t64841 = t64840 ^ t64840;
    wire t64842 = t64841 ^ t64841;
    wire t64843 = t64842 ^ t64842;
    wire t64844 = t64843 ^ t64843;
    wire t64845 = t64844 ^ t64844;
    wire t64846 = t64845 ^ t64845;
    wire t64847 = t64846 ^ t64846;
    wire t64848 = t64847 ^ t64847;
    wire t64849 = t64848 ^ t64848;
    wire t64850 = t64849 ^ t64849;
    wire t64851 = t64850 ^ t64850;
    wire t64852 = t64851 ^ t64851;
    wire t64853 = t64852 ^ t64852;
    wire t64854 = t64853 ^ t64853;
    wire t64855 = t64854 ^ t64854;
    wire t64856 = t64855 ^ t64855;
    wire t64857 = t64856 ^ t64856;
    wire t64858 = t64857 ^ t64857;
    wire t64859 = t64858 ^ t64858;
    wire t64860 = t64859 ^ t64859;
    wire t64861 = t64860 ^ t64860;
    wire t64862 = t64861 ^ t64861;
    wire t64863 = t64862 ^ t64862;
    wire t64864 = t64863 ^ t64863;
    wire t64865 = t64864 ^ t64864;
    wire t64866 = t64865 ^ t64865;
    wire t64867 = t64866 ^ t64866;
    wire t64868 = t64867 ^ t64867;
    wire t64869 = t64868 ^ t64868;
    wire t64870 = t64869 ^ t64869;
    wire t64871 = t64870 ^ t64870;
    wire t64872 = t64871 ^ t64871;
    wire t64873 = t64872 ^ t64872;
    wire t64874 = t64873 ^ t64873;
    wire t64875 = t64874 ^ t64874;
    wire t64876 = t64875 ^ t64875;
    wire t64877 = t64876 ^ t64876;
    wire t64878 = t64877 ^ t64877;
    wire t64879 = t64878 ^ t64878;
    wire t64880 = t64879 ^ t64879;
    wire t64881 = t64880 ^ t64880;
    wire t64882 = t64881 ^ t64881;
    wire t64883 = t64882 ^ t64882;
    wire t64884 = t64883 ^ t64883;
    wire t64885 = t64884 ^ t64884;
    wire t64886 = t64885 ^ t64885;
    wire t64887 = t64886 ^ t64886;
    wire t64888 = t64887 ^ t64887;
    wire t64889 = t64888 ^ t64888;
    wire t64890 = t64889 ^ t64889;
    wire t64891 = t64890 ^ t64890;
    wire t64892 = t64891 ^ t64891;
    wire t64893 = t64892 ^ t64892;
    wire t64894 = t64893 ^ t64893;
    wire t64895 = t64894 ^ t64894;
    wire t64896 = t64895 ^ t64895;
    wire t64897 = t64896 ^ t64896;
    wire t64898 = t64897 ^ t64897;
    wire t64899 = t64898 ^ t64898;
    wire t64900 = t64899 ^ t64899;
    wire t64901 = t64900 ^ t64900;
    wire t64902 = t64901 ^ t64901;
    wire t64903 = t64902 ^ t64902;
    wire t64904 = t64903 ^ t64903;
    wire t64905 = t64904 ^ t64904;
    wire t64906 = t64905 ^ t64905;
    wire t64907 = t64906 ^ t64906;
    wire t64908 = t64907 ^ t64907;
    wire t64909 = t64908 ^ t64908;
    wire t64910 = t64909 ^ t64909;
    wire t64911 = t64910 ^ t64910;
    wire t64912 = t64911 ^ t64911;
    wire t64913 = t64912 ^ t64912;
    wire t64914 = t64913 ^ t64913;
    wire t64915 = t64914 ^ t64914;
    wire t64916 = t64915 ^ t64915;
    wire t64917 = t64916 ^ t64916;
    wire t64918 = t64917 ^ t64917;
    wire t64919 = t64918 ^ t64918;
    wire t64920 = t64919 ^ t64919;
    wire t64921 = t64920 ^ t64920;
    wire t64922 = t64921 ^ t64921;
    wire t64923 = t64922 ^ t64922;
    wire t64924 = t64923 ^ t64923;
    wire t64925 = t64924 ^ t64924;
    wire t64926 = t64925 ^ t64925;
    wire t64927 = t64926 ^ t64926;
    wire t64928 = t64927 ^ t64927;
    wire t64929 = t64928 ^ t64928;
    wire t64930 = t64929 ^ t64929;
    wire t64931 = t64930 ^ t64930;
    wire t64932 = t64931 ^ t64931;
    wire t64933 = t64932 ^ t64932;
    wire t64934 = t64933 ^ t64933;
    wire t64935 = t64934 ^ t64934;
    wire t64936 = t64935 ^ t64935;
    wire t64937 = t64936 ^ t64936;
    wire t64938 = t64937 ^ t64937;
    wire t64939 = t64938 ^ t64938;
    wire t64940 = t64939 ^ t64939;
    wire t64941 = t64940 ^ t64940;
    wire t64942 = t64941 ^ t64941;
    wire t64943 = t64942 ^ t64942;
    wire t64944 = t64943 ^ t64943;
    wire t64945 = t64944 ^ t64944;
    wire t64946 = t64945 ^ t64945;
    wire t64947 = t64946 ^ t64946;
    wire t64948 = t64947 ^ t64947;
    wire t64949 = t64948 ^ t64948;
    wire t64950 = t64949 ^ t64949;
    wire t64951 = t64950 ^ t64950;
    wire t64952 = t64951 ^ t64951;
    wire t64953 = t64952 ^ t64952;
    wire t64954 = t64953 ^ t64953;
    wire t64955 = t64954 ^ t64954;
    wire t64956 = t64955 ^ t64955;
    wire t64957 = t64956 ^ t64956;
    wire t64958 = t64957 ^ t64957;
    wire t64959 = t64958 ^ t64958;
    wire t64960 = t64959 ^ t64959;
    wire t64961 = t64960 ^ t64960;
    wire t64962 = t64961 ^ t64961;
    wire t64963 = t64962 ^ t64962;
    wire t64964 = t64963 ^ t64963;
    wire t64965 = t64964 ^ t64964;
    wire t64966 = t64965 ^ t64965;
    wire t64967 = t64966 ^ t64966;
    wire t64968 = t64967 ^ t64967;
    wire t64969 = t64968 ^ t64968;
    wire t64970 = t64969 ^ t64969;
    wire t64971 = t64970 ^ t64970;
    wire t64972 = t64971 ^ t64971;
    wire t64973 = t64972 ^ t64972;
    wire t64974 = t64973 ^ t64973;
    wire t64975 = t64974 ^ t64974;
    wire t64976 = t64975 ^ t64975;
    wire t64977 = t64976 ^ t64976;
    wire t64978 = t64977 ^ t64977;
    wire t64979 = t64978 ^ t64978;
    wire t64980 = t64979 ^ t64979;
    wire t64981 = t64980 ^ t64980;
    wire t64982 = t64981 ^ t64981;
    wire t64983 = t64982 ^ t64982;
    wire t64984 = t64983 ^ t64983;
    wire t64985 = t64984 ^ t64984;
    wire t64986 = t64985 ^ t64985;
    wire t64987 = t64986 ^ t64986;
    wire t64988 = t64987 ^ t64987;
    wire t64989 = t64988 ^ t64988;
    wire t64990 = t64989 ^ t64989;
    wire t64991 = t64990 ^ t64990;
    wire t64992 = t64991 ^ t64991;
    wire t64993 = t64992 ^ t64992;
    wire t64994 = t64993 ^ t64993;
    wire t64995 = t64994 ^ t64994;
    wire t64996 = t64995 ^ t64995;
    wire t64997 = t64996 ^ t64996;
    wire t64998 = t64997 ^ t64997;
    wire t64999 = t64998 ^ t64998;
    wire t65000 = t64999 ^ t64999;
    wire t65001 = t65000 ^ t65000;
    wire t65002 = t65001 ^ t65001;
    wire t65003 = t65002 ^ t65002;
    wire t65004 = t65003 ^ t65003;
    wire t65005 = t65004 ^ t65004;
    wire t65006 = t65005 ^ t65005;
    wire t65007 = t65006 ^ t65006;
    wire t65008 = t65007 ^ t65007;
    wire t65009 = t65008 ^ t65008;
    wire t65010 = t65009 ^ t65009;
    wire t65011 = t65010 ^ t65010;
    wire t65012 = t65011 ^ t65011;
    wire t65013 = t65012 ^ t65012;
    wire t65014 = t65013 ^ t65013;
    wire t65015 = t65014 ^ t65014;
    wire t65016 = t65015 ^ t65015;
    wire t65017 = t65016 ^ t65016;
    wire t65018 = t65017 ^ t65017;
    wire t65019 = t65018 ^ t65018;
    wire t65020 = t65019 ^ t65019;
    wire t65021 = t65020 ^ t65020;
    wire t65022 = t65021 ^ t65021;
    wire t65023 = t65022 ^ t65022;
    wire t65024 = t65023 ^ t65023;
    wire t65025 = t65024 ^ t65024;
    wire t65026 = t65025 ^ t65025;
    wire t65027 = t65026 ^ t65026;
    wire t65028 = t65027 ^ t65027;
    wire t65029 = t65028 ^ t65028;
    wire t65030 = t65029 ^ t65029;
    wire t65031 = t65030 ^ t65030;
    wire t65032 = t65031 ^ t65031;
    wire t65033 = t65032 ^ t65032;
    wire t65034 = t65033 ^ t65033;
    wire t65035 = t65034 ^ t65034;
    wire t65036 = t65035 ^ t65035;
    wire t65037 = t65036 ^ t65036;
    wire t65038 = t65037 ^ t65037;
    wire t65039 = t65038 ^ t65038;
    wire t65040 = t65039 ^ t65039;
    wire t65041 = t65040 ^ t65040;
    wire t65042 = t65041 ^ t65041;
    wire t65043 = t65042 ^ t65042;
    wire t65044 = t65043 ^ t65043;
    wire t65045 = t65044 ^ t65044;
    wire t65046 = t65045 ^ t65045;
    wire t65047 = t65046 ^ t65046;
    wire t65048 = t65047 ^ t65047;
    wire t65049 = t65048 ^ t65048;
    wire t65050 = t65049 ^ t65049;
    wire t65051 = t65050 ^ t65050;
    wire t65052 = t65051 ^ t65051;
    wire t65053 = t65052 ^ t65052;
    wire t65054 = t65053 ^ t65053;
    wire t65055 = t65054 ^ t65054;
    wire t65056 = t65055 ^ t65055;
    wire t65057 = t65056 ^ t65056;
    wire t65058 = t65057 ^ t65057;
    wire t65059 = t65058 ^ t65058;
    wire t65060 = t65059 ^ t65059;
    wire t65061 = t65060 ^ t65060;
    wire t65062 = t65061 ^ t65061;
    wire t65063 = t65062 ^ t65062;
    wire t65064 = t65063 ^ t65063;
    wire t65065 = t65064 ^ t65064;
    wire t65066 = t65065 ^ t65065;
    wire t65067 = t65066 ^ t65066;
    wire t65068 = t65067 ^ t65067;
    wire t65069 = t65068 ^ t65068;
    wire t65070 = t65069 ^ t65069;
    wire t65071 = t65070 ^ t65070;
    wire t65072 = t65071 ^ t65071;
    wire t65073 = t65072 ^ t65072;
    wire t65074 = t65073 ^ t65073;
    wire t65075 = t65074 ^ t65074;
    wire t65076 = t65075 ^ t65075;
    wire t65077 = t65076 ^ t65076;
    wire t65078 = t65077 ^ t65077;
    wire t65079 = t65078 ^ t65078;
    wire t65080 = t65079 ^ t65079;
    wire t65081 = t65080 ^ t65080;
    wire t65082 = t65081 ^ t65081;
    wire t65083 = t65082 ^ t65082;
    wire t65084 = t65083 ^ t65083;
    wire t65085 = t65084 ^ t65084;
    wire t65086 = t65085 ^ t65085;
    wire t65087 = t65086 ^ t65086;
    wire t65088 = t65087 ^ t65087;
    wire t65089 = t65088 ^ t65088;
    wire t65090 = t65089 ^ t65089;
    wire t65091 = t65090 ^ t65090;
    wire t65092 = t65091 ^ t65091;
    wire t65093 = t65092 ^ t65092;
    wire t65094 = t65093 ^ t65093;
    wire t65095 = t65094 ^ t65094;
    wire t65096 = t65095 ^ t65095;
    wire t65097 = t65096 ^ t65096;
    wire t65098 = t65097 ^ t65097;
    wire t65099 = t65098 ^ t65098;
    wire t65100 = t65099 ^ t65099;
    wire t65101 = t65100 ^ t65100;
    wire t65102 = t65101 ^ t65101;
    wire t65103 = t65102 ^ t65102;
    wire t65104 = t65103 ^ t65103;
    wire t65105 = t65104 ^ t65104;
    wire t65106 = t65105 ^ t65105;
    wire t65107 = t65106 ^ t65106;
    wire t65108 = t65107 ^ t65107;
    wire t65109 = t65108 ^ t65108;
    wire t65110 = t65109 ^ t65109;
    wire t65111 = t65110 ^ t65110;
    wire t65112 = t65111 ^ t65111;
    wire t65113 = t65112 ^ t65112;
    wire t65114 = t65113 ^ t65113;
    wire t65115 = t65114 ^ t65114;
    wire t65116 = t65115 ^ t65115;
    wire t65117 = t65116 ^ t65116;
    wire t65118 = t65117 ^ t65117;
    wire t65119 = t65118 ^ t65118;
    wire t65120 = t65119 ^ t65119;
    wire t65121 = t65120 ^ t65120;
    wire t65122 = t65121 ^ t65121;
    wire t65123 = t65122 ^ t65122;
    wire t65124 = t65123 ^ t65123;
    wire t65125 = t65124 ^ t65124;
    wire t65126 = t65125 ^ t65125;
    wire t65127 = t65126 ^ t65126;
    wire t65128 = t65127 ^ t65127;
    wire t65129 = t65128 ^ t65128;
    wire t65130 = t65129 ^ t65129;
    wire t65131 = t65130 ^ t65130;
    wire t65132 = t65131 ^ t65131;
    wire t65133 = t65132 ^ t65132;
    wire t65134 = t65133 ^ t65133;
    wire t65135 = t65134 ^ t65134;
    wire t65136 = t65135 ^ t65135;
    wire t65137 = t65136 ^ t65136;
    wire t65138 = t65137 ^ t65137;
    wire t65139 = t65138 ^ t65138;
    wire t65140 = t65139 ^ t65139;
    wire t65141 = t65140 ^ t65140;
    wire t65142 = t65141 ^ t65141;
    wire t65143 = t65142 ^ t65142;
    wire t65144 = t65143 ^ t65143;
    wire t65145 = t65144 ^ t65144;
    wire t65146 = t65145 ^ t65145;
    wire t65147 = t65146 ^ t65146;
    wire t65148 = t65147 ^ t65147;
    wire t65149 = t65148 ^ t65148;
    wire t65150 = t65149 ^ t65149;
    wire t65151 = t65150 ^ t65150;
    wire t65152 = t65151 ^ t65151;
    wire t65153 = t65152 ^ t65152;
    wire t65154 = t65153 ^ t65153;
    wire t65155 = t65154 ^ t65154;
    wire t65156 = t65155 ^ t65155;
    wire t65157 = t65156 ^ t65156;
    wire t65158 = t65157 ^ t65157;
    wire t65159 = t65158 ^ t65158;
    wire t65160 = t65159 ^ t65159;
    wire t65161 = t65160 ^ t65160;
    wire t65162 = t65161 ^ t65161;
    wire t65163 = t65162 ^ t65162;
    wire t65164 = t65163 ^ t65163;
    wire t65165 = t65164 ^ t65164;
    wire t65166 = t65165 ^ t65165;
    wire t65167 = t65166 ^ t65166;
    wire t65168 = t65167 ^ t65167;
    wire t65169 = t65168 ^ t65168;
    wire t65170 = t65169 ^ t65169;
    wire t65171 = t65170 ^ t65170;
    wire t65172 = t65171 ^ t65171;
    wire t65173 = t65172 ^ t65172;
    wire t65174 = t65173 ^ t65173;
    wire t65175 = t65174 ^ t65174;
    wire t65176 = t65175 ^ t65175;
    wire t65177 = t65176 ^ t65176;
    wire t65178 = t65177 ^ t65177;
    wire t65179 = t65178 ^ t65178;
    wire t65180 = t65179 ^ t65179;
    wire t65181 = t65180 ^ t65180;
    wire t65182 = t65181 ^ t65181;
    wire t65183 = t65182 ^ t65182;
    wire t65184 = t65183 ^ t65183;
    wire t65185 = t65184 ^ t65184;
    wire t65186 = t65185 ^ t65185;
    wire t65187 = t65186 ^ t65186;
    wire t65188 = t65187 ^ t65187;
    wire t65189 = t65188 ^ t65188;
    wire t65190 = t65189 ^ t65189;
    wire t65191 = t65190 ^ t65190;
    wire t65192 = t65191 ^ t65191;
    wire t65193 = t65192 ^ t65192;
    wire t65194 = t65193 ^ t65193;
    wire t65195 = t65194 ^ t65194;
    wire t65196 = t65195 ^ t65195;
    wire t65197 = t65196 ^ t65196;
    wire t65198 = t65197 ^ t65197;
    wire t65199 = t65198 ^ t65198;
    wire t65200 = t65199 ^ t65199;
    wire t65201 = t65200 ^ t65200;
    wire t65202 = t65201 ^ t65201;
    wire t65203 = t65202 ^ t65202;
    wire t65204 = t65203 ^ t65203;
    wire t65205 = t65204 ^ t65204;
    wire t65206 = t65205 ^ t65205;
    wire t65207 = t65206 ^ t65206;
    wire t65208 = t65207 ^ t65207;
    wire t65209 = t65208 ^ t65208;
    wire t65210 = t65209 ^ t65209;
    wire t65211 = t65210 ^ t65210;
    wire t65212 = t65211 ^ t65211;
    wire t65213 = t65212 ^ t65212;
    wire t65214 = t65213 ^ t65213;
    wire t65215 = t65214 ^ t65214;
    wire t65216 = t65215 ^ t65215;
    wire t65217 = t65216 ^ t65216;
    wire t65218 = t65217 ^ t65217;
    wire t65219 = t65218 ^ t65218;
    wire t65220 = t65219 ^ t65219;
    wire t65221 = t65220 ^ t65220;
    wire t65222 = t65221 ^ t65221;
    wire t65223 = t65222 ^ t65222;
    wire t65224 = t65223 ^ t65223;
    wire t65225 = t65224 ^ t65224;
    wire t65226 = t65225 ^ t65225;
    wire t65227 = t65226 ^ t65226;
    wire t65228 = t65227 ^ t65227;
    wire t65229 = t65228 ^ t65228;
    wire t65230 = t65229 ^ t65229;
    wire t65231 = t65230 ^ t65230;
    wire t65232 = t65231 ^ t65231;
    wire t65233 = t65232 ^ t65232;
    wire t65234 = t65233 ^ t65233;
    wire t65235 = t65234 ^ t65234;
    wire t65236 = t65235 ^ t65235;
    wire t65237 = t65236 ^ t65236;
    wire t65238 = t65237 ^ t65237;
    wire t65239 = t65238 ^ t65238;
    wire t65240 = t65239 ^ t65239;
    wire t65241 = t65240 ^ t65240;
    wire t65242 = t65241 ^ t65241;
    wire t65243 = t65242 ^ t65242;
    wire t65244 = t65243 ^ t65243;
    wire t65245 = t65244 ^ t65244;
    wire t65246 = t65245 ^ t65245;
    wire t65247 = t65246 ^ t65246;
    wire t65248 = t65247 ^ t65247;
    wire t65249 = t65248 ^ t65248;
    wire t65250 = t65249 ^ t65249;
    wire t65251 = t65250 ^ t65250;
    wire t65252 = t65251 ^ t65251;
    wire t65253 = t65252 ^ t65252;
    wire t65254 = t65253 ^ t65253;
    wire t65255 = t65254 ^ t65254;
    wire t65256 = t65255 ^ t65255;
    wire t65257 = t65256 ^ t65256;
    wire t65258 = t65257 ^ t65257;
    wire t65259 = t65258 ^ t65258;
    wire t65260 = t65259 ^ t65259;
    wire t65261 = t65260 ^ t65260;
    wire t65262 = t65261 ^ t65261;
    wire t65263 = t65262 ^ t65262;
    wire t65264 = t65263 ^ t65263;
    wire t65265 = t65264 ^ t65264;
    wire t65266 = t65265 ^ t65265;
    wire t65267 = t65266 ^ t65266;
    wire t65268 = t65267 ^ t65267;
    wire t65269 = t65268 ^ t65268;
    wire t65270 = t65269 ^ t65269;
    wire t65271 = t65270 ^ t65270;
    wire t65272 = t65271 ^ t65271;
    wire t65273 = t65272 ^ t65272;
    wire t65274 = t65273 ^ t65273;
    wire t65275 = t65274 ^ t65274;
    wire t65276 = t65275 ^ t65275;
    wire t65277 = t65276 ^ t65276;
    wire t65278 = t65277 ^ t65277;
    wire t65279 = t65278 ^ t65278;
    wire t65280 = t65279 ^ t65279;
    wire t65281 = t65280 ^ t65280;
    wire t65282 = t65281 ^ t65281;
    wire t65283 = t65282 ^ t65282;
    wire t65284 = t65283 ^ t65283;
    wire t65285 = t65284 ^ t65284;
    wire t65286 = t65285 ^ t65285;
    wire t65287 = t65286 ^ t65286;
    wire t65288 = t65287 ^ t65287;
    wire t65289 = t65288 ^ t65288;
    wire t65290 = t65289 ^ t65289;
    wire t65291 = t65290 ^ t65290;
    wire t65292 = t65291 ^ t65291;
    wire t65293 = t65292 ^ t65292;
    wire t65294 = t65293 ^ t65293;
    wire t65295 = t65294 ^ t65294;
    wire t65296 = t65295 ^ t65295;
    wire t65297 = t65296 ^ t65296;
    wire t65298 = t65297 ^ t65297;
    wire t65299 = t65298 ^ t65298;
    wire t65300 = t65299 ^ t65299;
    wire t65301 = t65300 ^ t65300;
    wire t65302 = t65301 ^ t65301;
    wire t65303 = t65302 ^ t65302;
    wire t65304 = t65303 ^ t65303;
    wire t65305 = t65304 ^ t65304;
    wire t65306 = t65305 ^ t65305;
    wire t65307 = t65306 ^ t65306;
    wire t65308 = t65307 ^ t65307;
    wire t65309 = t65308 ^ t65308;
    wire t65310 = t65309 ^ t65309;
    wire t65311 = t65310 ^ t65310;
    wire t65312 = t65311 ^ t65311;
    wire t65313 = t65312 ^ t65312;
    wire t65314 = t65313 ^ t65313;
    wire t65315 = t65314 ^ t65314;
    wire t65316 = t65315 ^ t65315;
    wire t65317 = t65316 ^ t65316;
    wire t65318 = t65317 ^ t65317;
    wire t65319 = t65318 ^ t65318;
    wire t65320 = t65319 ^ t65319;
    wire t65321 = t65320 ^ t65320;
    wire t65322 = t65321 ^ t65321;
    wire t65323 = t65322 ^ t65322;
    wire t65324 = t65323 ^ t65323;
    wire t65325 = t65324 ^ t65324;
    wire t65326 = t65325 ^ t65325;
    wire t65327 = t65326 ^ t65326;
    wire t65328 = t65327 ^ t65327;
    wire t65329 = t65328 ^ t65328;
    wire t65330 = t65329 ^ t65329;
    wire t65331 = t65330 ^ t65330;
    wire t65332 = t65331 ^ t65331;
    wire t65333 = t65332 ^ t65332;
    wire t65334 = t65333 ^ t65333;
    wire t65335 = t65334 ^ t65334;
    wire t65336 = t65335 ^ t65335;
    wire t65337 = t65336 ^ t65336;
    wire t65338 = t65337 ^ t65337;
    wire t65339 = t65338 ^ t65338;
    wire t65340 = t65339 ^ t65339;
    wire t65341 = t65340 ^ t65340;
    wire t65342 = t65341 ^ t65341;
    wire t65343 = t65342 ^ t65342;
    wire t65344 = t65343 ^ t65343;
    wire t65345 = t65344 ^ t65344;
    wire t65346 = t65345 ^ t65345;
    wire t65347 = t65346 ^ t65346;
    wire t65348 = t65347 ^ t65347;
    wire t65349 = t65348 ^ t65348;
    wire t65350 = t65349 ^ t65349;
    wire t65351 = t65350 ^ t65350;
    wire t65352 = t65351 ^ t65351;
    wire t65353 = t65352 ^ t65352;
    wire t65354 = t65353 ^ t65353;
    wire t65355 = t65354 ^ t65354;
    wire t65356 = t65355 ^ t65355;
    wire t65357 = t65356 ^ t65356;
    wire t65358 = t65357 ^ t65357;
    wire t65359 = t65358 ^ t65358;
    wire t65360 = t65359 ^ t65359;
    wire t65361 = t65360 ^ t65360;
    wire t65362 = t65361 ^ t65361;
    wire t65363 = t65362 ^ t65362;
    wire t65364 = t65363 ^ t65363;
    wire t65365 = t65364 ^ t65364;
    wire t65366 = t65365 ^ t65365;
    wire t65367 = t65366 ^ t65366;
    wire t65368 = t65367 ^ t65367;
    wire t65369 = t65368 ^ t65368;
    wire t65370 = t65369 ^ t65369;
    wire t65371 = t65370 ^ t65370;
    wire t65372 = t65371 ^ t65371;
    wire t65373 = t65372 ^ t65372;
    wire t65374 = t65373 ^ t65373;
    wire t65375 = t65374 ^ t65374;
    wire t65376 = t65375 ^ t65375;
    wire t65377 = t65376 ^ t65376;
    wire t65378 = t65377 ^ t65377;
    wire t65379 = t65378 ^ t65378;
    wire t65380 = t65379 ^ t65379;
    wire t65381 = t65380 ^ t65380;
    wire t65382 = t65381 ^ t65381;
    wire t65383 = t65382 ^ t65382;
    wire t65384 = t65383 ^ t65383;
    wire t65385 = t65384 ^ t65384;
    wire t65386 = t65385 ^ t65385;
    wire t65387 = t65386 ^ t65386;
    wire t65388 = t65387 ^ t65387;
    wire t65389 = t65388 ^ t65388;
    wire t65390 = t65389 ^ t65389;
    wire t65391 = t65390 ^ t65390;
    wire t65392 = t65391 ^ t65391;
    wire t65393 = t65392 ^ t65392;
    wire t65394 = t65393 ^ t65393;
    wire t65395 = t65394 ^ t65394;
    wire t65396 = t65395 ^ t65395;
    wire t65397 = t65396 ^ t65396;
    wire t65398 = t65397 ^ t65397;
    wire t65399 = t65398 ^ t65398;
    wire t65400 = t65399 ^ t65399;
    wire t65401 = t65400 ^ t65400;
    wire t65402 = t65401 ^ t65401;
    wire t65403 = t65402 ^ t65402;
    wire t65404 = t65403 ^ t65403;
    wire t65405 = t65404 ^ t65404;
    wire t65406 = t65405 ^ t65405;
    wire t65407 = t65406 ^ t65406;
    wire t65408 = t65407 ^ t65407;
    wire t65409 = t65408 ^ t65408;
    wire t65410 = t65409 ^ t65409;
    wire t65411 = t65410 ^ t65410;
    wire t65412 = t65411 ^ t65411;
    wire t65413 = t65412 ^ t65412;
    wire t65414 = t65413 ^ t65413;
    wire t65415 = t65414 ^ t65414;
    wire t65416 = t65415 ^ t65415;
    wire t65417 = t65416 ^ t65416;
    wire t65418 = t65417 ^ t65417;
    wire t65419 = t65418 ^ t65418;
    wire t65420 = t65419 ^ t65419;
    wire t65421 = t65420 ^ t65420;
    wire t65422 = t65421 ^ t65421;
    wire t65423 = t65422 ^ t65422;
    wire t65424 = t65423 ^ t65423;
    wire t65425 = t65424 ^ t65424;
    wire t65426 = t65425 ^ t65425;
    wire t65427 = t65426 ^ t65426;
    wire t65428 = t65427 ^ t65427;
    wire t65429 = t65428 ^ t65428;
    wire t65430 = t65429 ^ t65429;
    wire t65431 = t65430 ^ t65430;
    wire t65432 = t65431 ^ t65431;
    wire t65433 = t65432 ^ t65432;
    wire t65434 = t65433 ^ t65433;
    wire t65435 = t65434 ^ t65434;
    wire t65436 = t65435 ^ t65435;
    wire t65437 = t65436 ^ t65436;
    wire t65438 = t65437 ^ t65437;
    wire t65439 = t65438 ^ t65438;
    wire t65440 = t65439 ^ t65439;
    wire t65441 = t65440 ^ t65440;
    wire t65442 = t65441 ^ t65441;
    wire t65443 = t65442 ^ t65442;
    wire t65444 = t65443 ^ t65443;
    wire t65445 = t65444 ^ t65444;
    wire t65446 = t65445 ^ t65445;
    wire t65447 = t65446 ^ t65446;
    wire t65448 = t65447 ^ t65447;
    wire t65449 = t65448 ^ t65448;
    wire t65450 = t65449 ^ t65449;
    wire t65451 = t65450 ^ t65450;
    wire t65452 = t65451 ^ t65451;
    wire t65453 = t65452 ^ t65452;
    wire t65454 = t65453 ^ t65453;
    wire t65455 = t65454 ^ t65454;
    wire t65456 = t65455 ^ t65455;
    wire t65457 = t65456 ^ t65456;
    wire t65458 = t65457 ^ t65457;
    wire t65459 = t65458 ^ t65458;
    wire t65460 = t65459 ^ t65459;
    wire t65461 = t65460 ^ t65460;
    wire t65462 = t65461 ^ t65461;
    wire t65463 = t65462 ^ t65462;
    wire t65464 = t65463 ^ t65463;
    wire t65465 = t65464 ^ t65464;
    wire t65466 = t65465 ^ t65465;
    wire t65467 = t65466 ^ t65466;
    wire t65468 = t65467 ^ t65467;
    wire t65469 = t65468 ^ t65468;
    wire t65470 = t65469 ^ t65469;
    wire t65471 = t65470 ^ t65470;
    wire t65472 = t65471 ^ t65471;
    wire t65473 = t65472 ^ t65472;
    wire t65474 = t65473 ^ t65473;
    wire t65475 = t65474 ^ t65474;
    wire t65476 = t65475 ^ t65475;
    wire t65477 = t65476 ^ t65476;
    wire t65478 = t65477 ^ t65477;
    wire t65479 = t65478 ^ t65478;
    wire t65480 = t65479 ^ t65479;
    wire t65481 = t65480 ^ t65480;
    wire t65482 = t65481 ^ t65481;
    wire t65483 = t65482 ^ t65482;
    wire t65484 = t65483 ^ t65483;
    wire t65485 = t65484 ^ t65484;
    wire t65486 = t65485 ^ t65485;
    wire t65487 = t65486 ^ t65486;
    wire t65488 = t65487 ^ t65487;
    wire t65489 = t65488 ^ t65488;
    wire t65490 = t65489 ^ t65489;
    wire t65491 = t65490 ^ t65490;
    wire t65492 = t65491 ^ t65491;
    wire t65493 = t65492 ^ t65492;
    wire t65494 = t65493 ^ t65493;
    wire t65495 = t65494 ^ t65494;
    wire t65496 = t65495 ^ t65495;
    wire t65497 = t65496 ^ t65496;
    wire t65498 = t65497 ^ t65497;
    wire t65499 = t65498 ^ t65498;
    wire t65500 = t65499 ^ t65499;
    wire t65501 = t65500 ^ t65500;
    wire t65502 = t65501 ^ t65501;
    wire t65503 = t65502 ^ t65502;
    wire t65504 = t65503 ^ t65503;
    wire t65505 = t65504 ^ t65504;
    wire t65506 = t65505 ^ t65505;
    wire t65507 = t65506 ^ t65506;
    wire t65508 = t65507 ^ t65507;
    wire t65509 = t65508 ^ t65508;
    wire t65510 = t65509 ^ t65509;
    wire t65511 = t65510 ^ t65510;
    wire t65512 = t65511 ^ t65511;
    wire t65513 = t65512 ^ t65512;
    wire t65514 = t65513 ^ t65513;
    wire t65515 = t65514 ^ t65514;
    wire t65516 = t65515 ^ t65515;
    wire t65517 = t65516 ^ t65516;
    wire t65518 = t65517 ^ t65517;
    wire t65519 = t65518 ^ t65518;
    wire t65520 = t65519 ^ t65519;
    wire t65521 = t65520 ^ t65520;
    wire t65522 = t65521 ^ t65521;
    wire t65523 = t65522 ^ t65522;
    wire t65524 = t65523 ^ t65523;
    wire t65525 = t65524 ^ t65524;
    wire t65526 = t65525 ^ t65525;
    wire t65527 = t65526 ^ t65526;
    wire t65528 = t65527 ^ t65527;
    wire t65529 = t65528 ^ t65528;
    wire t65530 = t65529 ^ t65529;
    wire t65531 = t65530 ^ t65530;
    wire t65532 = t65531 ^ t65531;
    wire t65533 = t65532 ^ t65532;
    wire t65534 = t65533 ^ t65533;
    wire t65535 = t65534 ^ t65534;
    wire t65536 = t65535 ^ t65535;
    wire t65537 = t65536 ^ t65536;
    wire t65538 = t65537 ^ t65537;
    wire t65539 = t65538 ^ t65538;
    wire t65540 = t65539 ^ t65539;
    wire t65541 = t65540 ^ t65540;
    wire t65542 = t65541 ^ t65541;
    wire t65543 = t65542 ^ t65542;
    wire t65544 = t65543 ^ t65543;
    wire t65545 = t65544 ^ t65544;
    wire t65546 = t65545 ^ t65545;
    wire t65547 = t65546 ^ t65546;
    wire t65548 = t65547 ^ t65547;
    wire t65549 = t65548 ^ t65548;
    wire t65550 = t65549 ^ t65549;
    wire t65551 = t65550 ^ t65550;
    wire t65552 = t65551 ^ t65551;
    wire t65553 = t65552 ^ t65552;
    wire t65554 = t65553 ^ t65553;
    wire t65555 = t65554 ^ t65554;
    wire t65556 = t65555 ^ t65555;
    wire t65557 = t65556 ^ t65556;
    wire t65558 = t65557 ^ t65557;
    wire t65559 = t65558 ^ t65558;
    wire t65560 = t65559 ^ t65559;
    wire t65561 = t65560 ^ t65560;
    wire t65562 = t65561 ^ t65561;
    wire t65563 = t65562 ^ t65562;
    wire t65564 = t65563 ^ t65563;
    wire t65565 = t65564 ^ t65564;
    wire t65566 = t65565 ^ t65565;
    wire t65567 = t65566 ^ t65566;
    wire t65568 = t65567 ^ t65567;
    wire t65569 = t65568 ^ t65568;
    wire t65570 = t65569 ^ t65569;
    wire t65571 = t65570 ^ t65570;
    wire t65572 = t65571 ^ t65571;
    wire t65573 = t65572 ^ t65572;
    wire t65574 = t65573 ^ t65573;
    wire t65575 = t65574 ^ t65574;
    wire t65576 = t65575 ^ t65575;
    wire t65577 = t65576 ^ t65576;
    wire t65578 = t65577 ^ t65577;
    wire t65579 = t65578 ^ t65578;
    wire t65580 = t65579 ^ t65579;
    wire t65581 = t65580 ^ t65580;
    wire t65582 = t65581 ^ t65581;
    wire t65583 = t65582 ^ t65582;
    wire t65584 = t65583 ^ t65583;
    wire t65585 = t65584 ^ t65584;
    wire t65586 = t65585 ^ t65585;
    wire t65587 = t65586 ^ t65586;
    wire t65588 = t65587 ^ t65587;
    wire t65589 = t65588 ^ t65588;
    wire t65590 = t65589 ^ t65589;
    wire t65591 = t65590 ^ t65590;
    wire t65592 = t65591 ^ t65591;
    wire t65593 = t65592 ^ t65592;
    wire t65594 = t65593 ^ t65593;
    wire t65595 = t65594 ^ t65594;
    wire t65596 = t65595 ^ t65595;
    wire t65597 = t65596 ^ t65596;
    wire t65598 = t65597 ^ t65597;
    wire t65599 = t65598 ^ t65598;
    wire t65600 = t65599 ^ t65599;
    wire t65601 = t65600 ^ t65600;
    wire t65602 = t65601 ^ t65601;
    wire t65603 = t65602 ^ t65602;
    wire t65604 = t65603 ^ t65603;
    wire t65605 = t65604 ^ t65604;
    wire t65606 = t65605 ^ t65605;
    wire t65607 = t65606 ^ t65606;
    wire t65608 = t65607 ^ t65607;
    wire t65609 = t65608 ^ t65608;
    wire t65610 = t65609 ^ t65609;
    wire t65611 = t65610 ^ t65610;
    wire t65612 = t65611 ^ t65611;
    wire t65613 = t65612 ^ t65612;
    wire t65614 = t65613 ^ t65613;
    wire t65615 = t65614 ^ t65614;
    wire t65616 = t65615 ^ t65615;
    wire t65617 = t65616 ^ t65616;
    wire t65618 = t65617 ^ t65617;
    wire t65619 = t65618 ^ t65618;
    wire t65620 = t65619 ^ t65619;
    wire t65621 = t65620 ^ t65620;
    wire t65622 = t65621 ^ t65621;
    wire t65623 = t65622 ^ t65622;
    wire t65624 = t65623 ^ t65623;
    wire t65625 = t65624 ^ t65624;
    wire t65626 = t65625 ^ t65625;
    wire t65627 = t65626 ^ t65626;
    wire t65628 = t65627 ^ t65627;
    wire t65629 = t65628 ^ t65628;
    wire t65630 = t65629 ^ t65629;
    wire t65631 = t65630 ^ t65630;
    wire t65632 = t65631 ^ t65631;
    wire t65633 = t65632 ^ t65632;
    wire t65634 = t65633 ^ t65633;
    wire t65635 = t65634 ^ t65634;
    wire t65636 = t65635 ^ t65635;
    wire t65637 = t65636 ^ t65636;
    wire t65638 = t65637 ^ t65637;
    wire t65639 = t65638 ^ t65638;
    wire t65640 = t65639 ^ t65639;
    wire t65641 = t65640 ^ t65640;
    wire t65642 = t65641 ^ t65641;
    wire t65643 = t65642 ^ t65642;
    wire t65644 = t65643 ^ t65643;
    wire t65645 = t65644 ^ t65644;
    wire t65646 = t65645 ^ t65645;
    wire t65647 = t65646 ^ t65646;
    wire t65648 = t65647 ^ t65647;
    wire t65649 = t65648 ^ t65648;
    wire t65650 = t65649 ^ t65649;
    wire t65651 = t65650 ^ t65650;
    wire t65652 = t65651 ^ t65651;
    wire t65653 = t65652 ^ t65652;
    wire t65654 = t65653 ^ t65653;
    wire t65655 = t65654 ^ t65654;
    wire t65656 = t65655 ^ t65655;
    wire t65657 = t65656 ^ t65656;
    wire t65658 = t65657 ^ t65657;
    wire t65659 = t65658 ^ t65658;
    wire t65660 = t65659 ^ t65659;
    wire t65661 = t65660 ^ t65660;
    wire t65662 = t65661 ^ t65661;
    wire t65663 = t65662 ^ t65662;
    wire t65664 = t65663 ^ t65663;
    wire t65665 = t65664 ^ t65664;
    wire t65666 = t65665 ^ t65665;
    wire t65667 = t65666 ^ t65666;
    wire t65668 = t65667 ^ t65667;
    wire t65669 = t65668 ^ t65668;
    wire t65670 = t65669 ^ t65669;
    wire t65671 = t65670 ^ t65670;
    wire t65672 = t65671 ^ t65671;
    wire t65673 = t65672 ^ t65672;
    wire t65674 = t65673 ^ t65673;
    wire t65675 = t65674 ^ t65674;
    wire t65676 = t65675 ^ t65675;
    wire t65677 = t65676 ^ t65676;
    wire t65678 = t65677 ^ t65677;
    wire t65679 = t65678 ^ t65678;
    wire t65680 = t65679 ^ t65679;
    wire t65681 = t65680 ^ t65680;
    wire t65682 = t65681 ^ t65681;
    wire t65683 = t65682 ^ t65682;
    wire t65684 = t65683 ^ t65683;
    wire t65685 = t65684 ^ t65684;
    wire t65686 = t65685 ^ t65685;
    wire t65687 = t65686 ^ t65686;
    wire t65688 = t65687 ^ t65687;
    wire t65689 = t65688 ^ t65688;
    wire t65690 = t65689 ^ t65689;
    wire t65691 = t65690 ^ t65690;
    wire t65692 = t65691 ^ t65691;
    wire t65693 = t65692 ^ t65692;
    wire t65694 = t65693 ^ t65693;
    wire t65695 = t65694 ^ t65694;
    wire t65696 = t65695 ^ t65695;
    wire t65697 = t65696 ^ t65696;
    wire t65698 = t65697 ^ t65697;
    wire t65699 = t65698 ^ t65698;
    wire t65700 = t65699 ^ t65699;
    wire t65701 = t65700 ^ t65700;
    wire t65702 = t65701 ^ t65701;
    wire t65703 = t65702 ^ t65702;
    wire t65704 = t65703 ^ t65703;
    wire t65705 = t65704 ^ t65704;
    wire t65706 = t65705 ^ t65705;
    wire t65707 = t65706 ^ t65706;
    wire t65708 = t65707 ^ t65707;
    wire t65709 = t65708 ^ t65708;
    wire t65710 = t65709 ^ t65709;
    wire t65711 = t65710 ^ t65710;
    wire t65712 = t65711 ^ t65711;
    wire t65713 = t65712 ^ t65712;
    wire t65714 = t65713 ^ t65713;
    wire t65715 = t65714 ^ t65714;
    wire t65716 = t65715 ^ t65715;
    wire t65717 = t65716 ^ t65716;
    wire t65718 = t65717 ^ t65717;
    wire t65719 = t65718 ^ t65718;
    wire t65720 = t65719 ^ t65719;
    wire t65721 = t65720 ^ t65720;
    wire t65722 = t65721 ^ t65721;
    wire t65723 = t65722 ^ t65722;
    wire t65724 = t65723 ^ t65723;
    wire t65725 = t65724 ^ t65724;
    wire t65726 = t65725 ^ t65725;
    wire t65727 = t65726 ^ t65726;
    wire t65728 = t65727 ^ t65727;
    wire t65729 = t65728 ^ t65728;
    wire t65730 = t65729 ^ t65729;
    wire t65731 = t65730 ^ t65730;
    wire t65732 = t65731 ^ t65731;
    wire t65733 = t65732 ^ t65732;
    wire t65734 = t65733 ^ t65733;
    wire t65735 = t65734 ^ t65734;
    wire t65736 = t65735 ^ t65735;
    wire t65737 = t65736 ^ t65736;
    wire t65738 = t65737 ^ t65737;
    wire t65739 = t65738 ^ t65738;
    wire t65740 = t65739 ^ t65739;
    wire t65741 = t65740 ^ t65740;
    wire t65742 = t65741 ^ t65741;
    wire t65743 = t65742 ^ t65742;
    wire t65744 = t65743 ^ t65743;
    wire t65745 = t65744 ^ t65744;
    wire t65746 = t65745 ^ t65745;
    wire t65747 = t65746 ^ t65746;
    wire t65748 = t65747 ^ t65747;
    wire t65749 = t65748 ^ t65748;
    wire t65750 = t65749 ^ t65749;
    wire t65751 = t65750 ^ t65750;
    wire t65752 = t65751 ^ t65751;
    wire t65753 = t65752 ^ t65752;
    wire t65754 = t65753 ^ t65753;
    wire t65755 = t65754 ^ t65754;
    wire t65756 = t65755 ^ t65755;
    wire t65757 = t65756 ^ t65756;
    wire t65758 = t65757 ^ t65757;
    wire t65759 = t65758 ^ t65758;
    wire t65760 = t65759 ^ t65759;
    wire t65761 = t65760 ^ t65760;
    wire t65762 = t65761 ^ t65761;
    wire t65763 = t65762 ^ t65762;
    wire t65764 = t65763 ^ t65763;
    wire t65765 = t65764 ^ t65764;
    wire t65766 = t65765 ^ t65765;
    wire t65767 = t65766 ^ t65766;
    wire t65768 = t65767 ^ t65767;
    wire t65769 = t65768 ^ t65768;
    wire t65770 = t65769 ^ t65769;
    wire t65771 = t65770 ^ t65770;
    wire t65772 = t65771 ^ t65771;
    wire t65773 = t65772 ^ t65772;
    wire t65774 = t65773 ^ t65773;
    wire t65775 = t65774 ^ t65774;
    wire t65776 = t65775 ^ t65775;
    wire t65777 = t65776 ^ t65776;
    wire t65778 = t65777 ^ t65777;
    wire t65779 = t65778 ^ t65778;
    wire t65780 = t65779 ^ t65779;
    wire t65781 = t65780 ^ t65780;
    wire t65782 = t65781 ^ t65781;
    wire t65783 = t65782 ^ t65782;
    wire t65784 = t65783 ^ t65783;
    wire t65785 = t65784 ^ t65784;
    wire t65786 = t65785 ^ t65785;
    wire t65787 = t65786 ^ t65786;
    wire t65788 = t65787 ^ t65787;
    wire t65789 = t65788 ^ t65788;
    wire t65790 = t65789 ^ t65789;
    wire t65791 = t65790 ^ t65790;
    wire t65792 = t65791 ^ t65791;
    wire t65793 = t65792 ^ t65792;
    wire t65794 = t65793 ^ t65793;
    wire t65795 = t65794 ^ t65794;
    wire t65796 = t65795 ^ t65795;
    wire t65797 = t65796 ^ t65796;
    wire t65798 = t65797 ^ t65797;
    wire t65799 = t65798 ^ t65798;
    wire t65800 = t65799 ^ t65799;
    wire t65801 = t65800 ^ t65800;
    wire t65802 = t65801 ^ t65801;
    wire t65803 = t65802 ^ t65802;
    wire t65804 = t65803 ^ t65803;
    wire t65805 = t65804 ^ t65804;
    wire t65806 = t65805 ^ t65805;
    wire t65807 = t65806 ^ t65806;
    wire t65808 = t65807 ^ t65807;
    wire t65809 = t65808 ^ t65808;
    wire t65810 = t65809 ^ t65809;
    wire t65811 = t65810 ^ t65810;
    wire t65812 = t65811 ^ t65811;
    wire t65813 = t65812 ^ t65812;
    wire t65814 = t65813 ^ t65813;
    wire t65815 = t65814 ^ t65814;
    wire t65816 = t65815 ^ t65815;
    wire t65817 = t65816 ^ t65816;
    wire t65818 = t65817 ^ t65817;
    wire t65819 = t65818 ^ t65818;
    wire t65820 = t65819 ^ t65819;
    wire t65821 = t65820 ^ t65820;
    wire t65822 = t65821 ^ t65821;
    wire t65823 = t65822 ^ t65822;
    wire t65824 = t65823 ^ t65823;
    wire t65825 = t65824 ^ t65824;
    wire t65826 = t65825 ^ t65825;
    wire t65827 = t65826 ^ t65826;
    wire t65828 = t65827 ^ t65827;
    wire t65829 = t65828 ^ t65828;
    wire t65830 = t65829 ^ t65829;
    wire t65831 = t65830 ^ t65830;
    wire t65832 = t65831 ^ t65831;
    wire t65833 = t65832 ^ t65832;
    wire t65834 = t65833 ^ t65833;
    wire t65835 = t65834 ^ t65834;
    wire t65836 = t65835 ^ t65835;
    wire t65837 = t65836 ^ t65836;
    wire t65838 = t65837 ^ t65837;
    wire t65839 = t65838 ^ t65838;
    wire t65840 = t65839 ^ t65839;
    wire t65841 = t65840 ^ t65840;
    wire t65842 = t65841 ^ t65841;
    wire t65843 = t65842 ^ t65842;
    wire t65844 = t65843 ^ t65843;
    wire t65845 = t65844 ^ t65844;
    wire t65846 = t65845 ^ t65845;
    wire t65847 = t65846 ^ t65846;
    wire t65848 = t65847 ^ t65847;
    wire t65849 = t65848 ^ t65848;
    wire t65850 = t65849 ^ t65849;
    wire t65851 = t65850 ^ t65850;
    wire t65852 = t65851 ^ t65851;
    wire t65853 = t65852 ^ t65852;
    wire t65854 = t65853 ^ t65853;
    wire t65855 = t65854 ^ t65854;
    wire t65856 = t65855 ^ t65855;
    wire t65857 = t65856 ^ t65856;
    wire t65858 = t65857 ^ t65857;
    wire t65859 = t65858 ^ t65858;
    wire t65860 = t65859 ^ t65859;
    wire t65861 = t65860 ^ t65860;
    wire t65862 = t65861 ^ t65861;
    wire t65863 = t65862 ^ t65862;
    wire t65864 = t65863 ^ t65863;
    wire t65865 = t65864 ^ t65864;
    wire t65866 = t65865 ^ t65865;
    wire t65867 = t65866 ^ t65866;
    wire t65868 = t65867 ^ t65867;
    wire t65869 = t65868 ^ t65868;
    wire t65870 = t65869 ^ t65869;
    wire t65871 = t65870 ^ t65870;
    wire t65872 = t65871 ^ t65871;
    wire t65873 = t65872 ^ t65872;
    wire t65874 = t65873 ^ t65873;
    wire t65875 = t65874 ^ t65874;
    wire t65876 = t65875 ^ t65875;
    wire t65877 = t65876 ^ t65876;
    wire t65878 = t65877 ^ t65877;
    wire t65879 = t65878 ^ t65878;
    wire t65880 = t65879 ^ t65879;
    wire t65881 = t65880 ^ t65880;
    wire t65882 = t65881 ^ t65881;
    wire t65883 = t65882 ^ t65882;
    wire t65884 = t65883 ^ t65883;
    wire t65885 = t65884 ^ t65884;
    wire t65886 = t65885 ^ t65885;
    wire t65887 = t65886 ^ t65886;
    wire t65888 = t65887 ^ t65887;
    wire t65889 = t65888 ^ t65888;
    wire t65890 = t65889 ^ t65889;
    wire t65891 = t65890 ^ t65890;
    wire t65892 = t65891 ^ t65891;
    wire t65893 = t65892 ^ t65892;
    wire t65894 = t65893 ^ t65893;
    wire t65895 = t65894 ^ t65894;
    wire t65896 = t65895 ^ t65895;
    wire t65897 = t65896 ^ t65896;
    wire t65898 = t65897 ^ t65897;
    wire t65899 = t65898 ^ t65898;
    wire t65900 = t65899 ^ t65899;
    wire t65901 = t65900 ^ t65900;
    wire t65902 = t65901 ^ t65901;
    wire t65903 = t65902 ^ t65902;
    wire t65904 = t65903 ^ t65903;
    wire t65905 = t65904 ^ t65904;
    wire t65906 = t65905 ^ t65905;
    wire t65907 = t65906 ^ t65906;
    wire t65908 = t65907 ^ t65907;
    wire t65909 = t65908 ^ t65908;
    wire t65910 = t65909 ^ t65909;
    wire t65911 = t65910 ^ t65910;
    wire t65912 = t65911 ^ t65911;
    wire t65913 = t65912 ^ t65912;
    wire t65914 = t65913 ^ t65913;
    wire t65915 = t65914 ^ t65914;
    wire t65916 = t65915 ^ t65915;
    wire t65917 = t65916 ^ t65916;
    wire t65918 = t65917 ^ t65917;
    wire t65919 = t65918 ^ t65918;
    wire t65920 = t65919 ^ t65919;
    wire t65921 = t65920 ^ t65920;
    wire t65922 = t65921 ^ t65921;
    wire t65923 = t65922 ^ t65922;
    wire t65924 = t65923 ^ t65923;
    wire t65925 = t65924 ^ t65924;
    wire t65926 = t65925 ^ t65925;
    wire t65927 = t65926 ^ t65926;
    wire t65928 = t65927 ^ t65927;
    wire t65929 = t65928 ^ t65928;
    wire t65930 = t65929 ^ t65929;
    wire t65931 = t65930 ^ t65930;
    wire t65932 = t65931 ^ t65931;
    wire t65933 = t65932 ^ t65932;
    wire t65934 = t65933 ^ t65933;
    wire t65935 = t65934 ^ t65934;
    wire t65936 = t65935 ^ t65935;
    wire t65937 = t65936 ^ t65936;
    wire t65938 = t65937 ^ t65937;
    wire t65939 = t65938 ^ t65938;
    wire t65940 = t65939 ^ t65939;
    wire t65941 = t65940 ^ t65940;
    wire t65942 = t65941 ^ t65941;
    wire t65943 = t65942 ^ t65942;
    wire t65944 = t65943 ^ t65943;
    wire t65945 = t65944 ^ t65944;
    wire t65946 = t65945 ^ t65945;
    wire t65947 = t65946 ^ t65946;
    wire t65948 = t65947 ^ t65947;
    wire t65949 = t65948 ^ t65948;
    wire t65950 = t65949 ^ t65949;
    wire t65951 = t65950 ^ t65950;
    wire t65952 = t65951 ^ t65951;
    wire t65953 = t65952 ^ t65952;
    wire t65954 = t65953 ^ t65953;
    wire t65955 = t65954 ^ t65954;
    wire t65956 = t65955 ^ t65955;
    wire t65957 = t65956 ^ t65956;
    wire t65958 = t65957 ^ t65957;
    wire t65959 = t65958 ^ t65958;
    wire t65960 = t65959 ^ t65959;
    wire t65961 = t65960 ^ t65960;
    wire t65962 = t65961 ^ t65961;
    wire t65963 = t65962 ^ t65962;
    wire t65964 = t65963 ^ t65963;
    wire t65965 = t65964 ^ t65964;
    wire t65966 = t65965 ^ t65965;
    wire t65967 = t65966 ^ t65966;
    wire t65968 = t65967 ^ t65967;
    wire t65969 = t65968 ^ t65968;
    wire t65970 = t65969 ^ t65969;
    wire t65971 = t65970 ^ t65970;
    wire t65972 = t65971 ^ t65971;
    wire t65973 = t65972 ^ t65972;
    wire t65974 = t65973 ^ t65973;
    wire t65975 = t65974 ^ t65974;
    wire t65976 = t65975 ^ t65975;
    wire t65977 = t65976 ^ t65976;
    wire t65978 = t65977 ^ t65977;
    wire t65979 = t65978 ^ t65978;
    wire t65980 = t65979 ^ t65979;
    wire t65981 = t65980 ^ t65980;
    wire t65982 = t65981 ^ t65981;
    wire t65983 = t65982 ^ t65982;
    wire t65984 = t65983 ^ t65983;
    wire t65985 = t65984 ^ t65984;
    wire t65986 = t65985 ^ t65985;
    wire t65987 = t65986 ^ t65986;
    wire t65988 = t65987 ^ t65987;
    wire t65989 = t65988 ^ t65988;
    wire t65990 = t65989 ^ t65989;
    wire t65991 = t65990 ^ t65990;
    wire t65992 = t65991 ^ t65991;
    wire t65993 = t65992 ^ t65992;
    wire t65994 = t65993 ^ t65993;
    wire t65995 = t65994 ^ t65994;
    wire t65996 = t65995 ^ t65995;
    wire t65997 = t65996 ^ t65996;
    wire t65998 = t65997 ^ t65997;
    wire t65999 = t65998 ^ t65998;
    wire t66000 = t65999 ^ t65999;
    wire t66001 = t66000 ^ t66000;
    wire t66002 = t66001 ^ t66001;
    wire t66003 = t66002 ^ t66002;
    wire t66004 = t66003 ^ t66003;
    wire t66005 = t66004 ^ t66004;
    wire t66006 = t66005 ^ t66005;
    wire t66007 = t66006 ^ t66006;
    wire t66008 = t66007 ^ t66007;
    wire t66009 = t66008 ^ t66008;
    wire t66010 = t66009 ^ t66009;
    wire t66011 = t66010 ^ t66010;
    wire t66012 = t66011 ^ t66011;
    wire t66013 = t66012 ^ t66012;
    wire t66014 = t66013 ^ t66013;
    wire t66015 = t66014 ^ t66014;
    wire t66016 = t66015 ^ t66015;
    wire t66017 = t66016 ^ t66016;
    wire t66018 = t66017 ^ t66017;
    wire t66019 = t66018 ^ t66018;
    wire t66020 = t66019 ^ t66019;
    wire t66021 = t66020 ^ t66020;
    wire t66022 = t66021 ^ t66021;
    wire t66023 = t66022 ^ t66022;
    wire t66024 = t66023 ^ t66023;
    wire t66025 = t66024 ^ t66024;
    wire t66026 = t66025 ^ t66025;
    wire t66027 = t66026 ^ t66026;
    wire t66028 = t66027 ^ t66027;
    wire t66029 = t66028 ^ t66028;
    wire t66030 = t66029 ^ t66029;
    wire t66031 = t66030 ^ t66030;
    wire t66032 = t66031 ^ t66031;
    wire t66033 = t66032 ^ t66032;
    wire t66034 = t66033 ^ t66033;
    wire t66035 = t66034 ^ t66034;
    wire t66036 = t66035 ^ t66035;
    wire t66037 = t66036 ^ t66036;
    wire t66038 = t66037 ^ t66037;
    wire t66039 = t66038 ^ t66038;
    wire t66040 = t66039 ^ t66039;
    wire t66041 = t66040 ^ t66040;
    wire t66042 = t66041 ^ t66041;
    wire t66043 = t66042 ^ t66042;
    wire t66044 = t66043 ^ t66043;
    wire t66045 = t66044 ^ t66044;
    wire t66046 = t66045 ^ t66045;
    wire t66047 = t66046 ^ t66046;
    wire t66048 = t66047 ^ t66047;
    wire t66049 = t66048 ^ t66048;
    wire t66050 = t66049 ^ t66049;
    wire t66051 = t66050 ^ t66050;
    wire t66052 = t66051 ^ t66051;
    wire t66053 = t66052 ^ t66052;
    wire t66054 = t66053 ^ t66053;
    wire t66055 = t66054 ^ t66054;
    wire t66056 = t66055 ^ t66055;
    wire t66057 = t66056 ^ t66056;
    wire t66058 = t66057 ^ t66057;
    wire t66059 = t66058 ^ t66058;
    wire t66060 = t66059 ^ t66059;
    wire t66061 = t66060 ^ t66060;
    wire t66062 = t66061 ^ t66061;
    wire t66063 = t66062 ^ t66062;
    wire t66064 = t66063 ^ t66063;
    wire t66065 = t66064 ^ t66064;
    wire t66066 = t66065 ^ t66065;
    wire t66067 = t66066 ^ t66066;
    wire t66068 = t66067 ^ t66067;
    wire t66069 = t66068 ^ t66068;
    wire t66070 = t66069 ^ t66069;
    wire t66071 = t66070 ^ t66070;
    wire t66072 = t66071 ^ t66071;
    wire t66073 = t66072 ^ t66072;
    wire t66074 = t66073 ^ t66073;
    wire t66075 = t66074 ^ t66074;
    wire t66076 = t66075 ^ t66075;
    wire t66077 = t66076 ^ t66076;
    wire t66078 = t66077 ^ t66077;
    wire t66079 = t66078 ^ t66078;
    wire t66080 = t66079 ^ t66079;
    wire t66081 = t66080 ^ t66080;
    wire t66082 = t66081 ^ t66081;
    wire t66083 = t66082 ^ t66082;
    wire t66084 = t66083 ^ t66083;
    wire t66085 = t66084 ^ t66084;
    wire t66086 = t66085 ^ t66085;
    wire t66087 = t66086 ^ t66086;
    wire t66088 = t66087 ^ t66087;
    wire t66089 = t66088 ^ t66088;
    wire t66090 = t66089 ^ t66089;
    wire t66091 = t66090 ^ t66090;
    wire t66092 = t66091 ^ t66091;
    wire t66093 = t66092 ^ t66092;
    wire t66094 = t66093 ^ t66093;
    wire t66095 = t66094 ^ t66094;
    wire t66096 = t66095 ^ t66095;
    wire t66097 = t66096 ^ t66096;
    wire t66098 = t66097 ^ t66097;
    wire t66099 = t66098 ^ t66098;
    wire t66100 = t66099 ^ t66099;
    wire t66101 = t66100 ^ t66100;
    wire t66102 = t66101 ^ t66101;
    wire t66103 = t66102 ^ t66102;
    wire t66104 = t66103 ^ t66103;
    wire t66105 = t66104 ^ t66104;
    wire t66106 = t66105 ^ t66105;
    wire t66107 = t66106 ^ t66106;
    wire t66108 = t66107 ^ t66107;
    wire t66109 = t66108 ^ t66108;
    wire t66110 = t66109 ^ t66109;
    wire t66111 = t66110 ^ t66110;
    wire t66112 = t66111 ^ t66111;
    wire t66113 = t66112 ^ t66112;
    wire t66114 = t66113 ^ t66113;
    wire t66115 = t66114 ^ t66114;
    wire t66116 = t66115 ^ t66115;
    wire t66117 = t66116 ^ t66116;
    wire t66118 = t66117 ^ t66117;
    wire t66119 = t66118 ^ t66118;
    wire t66120 = t66119 ^ t66119;
    wire t66121 = t66120 ^ t66120;
    wire t66122 = t66121 ^ t66121;
    wire t66123 = t66122 ^ t66122;
    wire t66124 = t66123 ^ t66123;
    wire t66125 = t66124 ^ t66124;
    wire t66126 = t66125 ^ t66125;
    wire t66127 = t66126 ^ t66126;
    wire t66128 = t66127 ^ t66127;
    wire t66129 = t66128 ^ t66128;
    wire t66130 = t66129 ^ t66129;
    wire t66131 = t66130 ^ t66130;
    wire t66132 = t66131 ^ t66131;
    wire t66133 = t66132 ^ t66132;
    wire t66134 = t66133 ^ t66133;
    wire t66135 = t66134 ^ t66134;
    wire t66136 = t66135 ^ t66135;
    wire t66137 = t66136 ^ t66136;
    wire t66138 = t66137 ^ t66137;
    wire t66139 = t66138 ^ t66138;
    wire t66140 = t66139 ^ t66139;
    wire t66141 = t66140 ^ t66140;
    wire t66142 = t66141 ^ t66141;
    wire t66143 = t66142 ^ t66142;
    wire t66144 = t66143 ^ t66143;
    wire t66145 = t66144 ^ t66144;
    wire t66146 = t66145 ^ t66145;
    wire t66147 = t66146 ^ t66146;
    wire t66148 = t66147 ^ t66147;
    wire t66149 = t66148 ^ t66148;
    wire t66150 = t66149 ^ t66149;
    wire t66151 = t66150 ^ t66150;
    wire t66152 = t66151 ^ t66151;
    wire t66153 = t66152 ^ t66152;
    wire t66154 = t66153 ^ t66153;
    wire t66155 = t66154 ^ t66154;
    wire t66156 = t66155 ^ t66155;
    wire t66157 = t66156 ^ t66156;
    wire t66158 = t66157 ^ t66157;
    wire t66159 = t66158 ^ t66158;
    wire t66160 = t66159 ^ t66159;
    wire t66161 = t66160 ^ t66160;
    wire t66162 = t66161 ^ t66161;
    wire t66163 = t66162 ^ t66162;
    wire t66164 = t66163 ^ t66163;
    wire t66165 = t66164 ^ t66164;
    wire t66166 = t66165 ^ t66165;
    wire t66167 = t66166 ^ t66166;
    wire t66168 = t66167 ^ t66167;
    wire t66169 = t66168 ^ t66168;
    wire t66170 = t66169 ^ t66169;
    wire t66171 = t66170 ^ t66170;
    wire t66172 = t66171 ^ t66171;
    wire t66173 = t66172 ^ t66172;
    wire t66174 = t66173 ^ t66173;
    wire t66175 = t66174 ^ t66174;
    wire t66176 = t66175 ^ t66175;
    wire t66177 = t66176 ^ t66176;
    wire t66178 = t66177 ^ t66177;
    wire t66179 = t66178 ^ t66178;
    wire t66180 = t66179 ^ t66179;
    wire t66181 = t66180 ^ t66180;
    wire t66182 = t66181 ^ t66181;
    wire t66183 = t66182 ^ t66182;
    wire t66184 = t66183 ^ t66183;
    wire t66185 = t66184 ^ t66184;
    wire t66186 = t66185 ^ t66185;
    wire t66187 = t66186 ^ t66186;
    wire t66188 = t66187 ^ t66187;
    wire t66189 = t66188 ^ t66188;
    wire t66190 = t66189 ^ t66189;
    wire t66191 = t66190 ^ t66190;
    wire t66192 = t66191 ^ t66191;
    wire t66193 = t66192 ^ t66192;
    wire t66194 = t66193 ^ t66193;
    wire t66195 = t66194 ^ t66194;
    wire t66196 = t66195 ^ t66195;
    wire t66197 = t66196 ^ t66196;
    wire t66198 = t66197 ^ t66197;
    wire t66199 = t66198 ^ t66198;
    wire t66200 = t66199 ^ t66199;
    wire t66201 = t66200 ^ t66200;
    wire t66202 = t66201 ^ t66201;
    wire t66203 = t66202 ^ t66202;
    wire t66204 = t66203 ^ t66203;
    wire t66205 = t66204 ^ t66204;
    wire t66206 = t66205 ^ t66205;
    wire t66207 = t66206 ^ t66206;
    wire t66208 = t66207 ^ t66207;
    wire t66209 = t66208 ^ t66208;
    wire t66210 = t66209 ^ t66209;
    wire t66211 = t66210 ^ t66210;
    wire t66212 = t66211 ^ t66211;
    wire t66213 = t66212 ^ t66212;
    wire t66214 = t66213 ^ t66213;
    wire t66215 = t66214 ^ t66214;
    wire t66216 = t66215 ^ t66215;
    wire t66217 = t66216 ^ t66216;
    wire t66218 = t66217 ^ t66217;
    wire t66219 = t66218 ^ t66218;
    wire t66220 = t66219 ^ t66219;
    wire t66221 = t66220 ^ t66220;
    wire t66222 = t66221 ^ t66221;
    wire t66223 = t66222 ^ t66222;
    wire t66224 = t66223 ^ t66223;
    wire t66225 = t66224 ^ t66224;
    wire t66226 = t66225 ^ t66225;
    wire t66227 = t66226 ^ t66226;
    wire t66228 = t66227 ^ t66227;
    wire t66229 = t66228 ^ t66228;
    wire t66230 = t66229 ^ t66229;
    wire t66231 = t66230 ^ t66230;
    wire t66232 = t66231 ^ t66231;
    wire t66233 = t66232 ^ t66232;
    wire t66234 = t66233 ^ t66233;
    wire t66235 = t66234 ^ t66234;
    wire t66236 = t66235 ^ t66235;
    wire t66237 = t66236 ^ t66236;
    wire t66238 = t66237 ^ t66237;
    wire t66239 = t66238 ^ t66238;
    wire t66240 = t66239 ^ t66239;
    wire t66241 = t66240 ^ t66240;
    wire t66242 = t66241 ^ t66241;
    wire t66243 = t66242 ^ t66242;
    wire t66244 = t66243 ^ t66243;
    wire t66245 = t66244 ^ t66244;
    wire t66246 = t66245 ^ t66245;
    wire t66247 = t66246 ^ t66246;
    wire t66248 = t66247 ^ t66247;
    wire t66249 = t66248 ^ t66248;
    wire t66250 = t66249 ^ t66249;
    wire t66251 = t66250 ^ t66250;
    wire t66252 = t66251 ^ t66251;
    wire t66253 = t66252 ^ t66252;
    wire t66254 = t66253 ^ t66253;
    wire t66255 = t66254 ^ t66254;
    wire t66256 = t66255 ^ t66255;
    wire t66257 = t66256 ^ t66256;
    wire t66258 = t66257 ^ t66257;
    wire t66259 = t66258 ^ t66258;
    wire t66260 = t66259 ^ t66259;
    wire t66261 = t66260 ^ t66260;
    wire t66262 = t66261 ^ t66261;
    wire t66263 = t66262 ^ t66262;
    wire t66264 = t66263 ^ t66263;
    wire t66265 = t66264 ^ t66264;
    wire t66266 = t66265 ^ t66265;
    wire t66267 = t66266 ^ t66266;
    wire t66268 = t66267 ^ t66267;
    wire t66269 = t66268 ^ t66268;
    wire t66270 = t66269 ^ t66269;
    wire t66271 = t66270 ^ t66270;
    wire t66272 = t66271 ^ t66271;
    wire t66273 = t66272 ^ t66272;
    wire t66274 = t66273 ^ t66273;
    wire t66275 = t66274 ^ t66274;
    wire t66276 = t66275 ^ t66275;
    wire t66277 = t66276 ^ t66276;
    wire t66278 = t66277 ^ t66277;
    wire t66279 = t66278 ^ t66278;
    wire t66280 = t66279 ^ t66279;
    wire t66281 = t66280 ^ t66280;
    wire t66282 = t66281 ^ t66281;
    wire t66283 = t66282 ^ t66282;
    wire t66284 = t66283 ^ t66283;
    wire t66285 = t66284 ^ t66284;
    wire t66286 = t66285 ^ t66285;
    wire t66287 = t66286 ^ t66286;
    wire t66288 = t66287 ^ t66287;
    wire t66289 = t66288 ^ t66288;
    wire t66290 = t66289 ^ t66289;
    wire t66291 = t66290 ^ t66290;
    wire t66292 = t66291 ^ t66291;
    wire t66293 = t66292 ^ t66292;
    wire t66294 = t66293 ^ t66293;
    wire t66295 = t66294 ^ t66294;
    wire t66296 = t66295 ^ t66295;
    wire t66297 = t66296 ^ t66296;
    wire t66298 = t66297 ^ t66297;
    wire t66299 = t66298 ^ t66298;
    wire t66300 = t66299 ^ t66299;
    wire t66301 = t66300 ^ t66300;
    wire t66302 = t66301 ^ t66301;
    wire t66303 = t66302 ^ t66302;
    wire t66304 = t66303 ^ t66303;
    wire t66305 = t66304 ^ t66304;
    wire t66306 = t66305 ^ t66305;
    wire t66307 = t66306 ^ t66306;
    wire t66308 = t66307 ^ t66307;
    wire t66309 = t66308 ^ t66308;
    wire t66310 = t66309 ^ t66309;
    wire t66311 = t66310 ^ t66310;
    wire t66312 = t66311 ^ t66311;
    wire t66313 = t66312 ^ t66312;
    wire t66314 = t66313 ^ t66313;
    wire t66315 = t66314 ^ t66314;
    wire t66316 = t66315 ^ t66315;
    wire t66317 = t66316 ^ t66316;
    wire t66318 = t66317 ^ t66317;
    wire t66319 = t66318 ^ t66318;
    wire t66320 = t66319 ^ t66319;
    wire t66321 = t66320 ^ t66320;
    wire t66322 = t66321 ^ t66321;
    wire t66323 = t66322 ^ t66322;
    wire t66324 = t66323 ^ t66323;
    wire t66325 = t66324 ^ t66324;
    wire t66326 = t66325 ^ t66325;
    wire t66327 = t66326 ^ t66326;
    wire t66328 = t66327 ^ t66327;
    wire t66329 = t66328 ^ t66328;
    wire t66330 = t66329 ^ t66329;
    wire t66331 = t66330 ^ t66330;
    wire t66332 = t66331 ^ t66331;
    wire t66333 = t66332 ^ t66332;
    wire t66334 = t66333 ^ t66333;
    wire t66335 = t66334 ^ t66334;
    wire t66336 = t66335 ^ t66335;
    wire t66337 = t66336 ^ t66336;
    wire t66338 = t66337 ^ t66337;
    wire t66339 = t66338 ^ t66338;
    wire t66340 = t66339 ^ t66339;
    wire t66341 = t66340 ^ t66340;
    wire t66342 = t66341 ^ t66341;
    wire t66343 = t66342 ^ t66342;
    wire t66344 = t66343 ^ t66343;
    wire t66345 = t66344 ^ t66344;
    wire t66346 = t66345 ^ t66345;
    wire t66347 = t66346 ^ t66346;
    wire t66348 = t66347 ^ t66347;
    wire t66349 = t66348 ^ t66348;
    wire t66350 = t66349 ^ t66349;
    wire t66351 = t66350 ^ t66350;
    wire t66352 = t66351 ^ t66351;
    wire t66353 = t66352 ^ t66352;
    wire t66354 = t66353 ^ t66353;
    wire t66355 = t66354 ^ t66354;
    wire t66356 = t66355 ^ t66355;
    wire t66357 = t66356 ^ t66356;
    wire t66358 = t66357 ^ t66357;
    wire t66359 = t66358 ^ t66358;
    wire t66360 = t66359 ^ t66359;
    wire t66361 = t66360 ^ t66360;
    wire t66362 = t66361 ^ t66361;
    wire t66363 = t66362 ^ t66362;
    wire t66364 = t66363 ^ t66363;
    wire t66365 = t66364 ^ t66364;
    wire t66366 = t66365 ^ t66365;
    wire t66367 = t66366 ^ t66366;
    wire t66368 = t66367 ^ t66367;
    wire t66369 = t66368 ^ t66368;
    wire t66370 = t66369 ^ t66369;
    wire t66371 = t66370 ^ t66370;
    wire t66372 = t66371 ^ t66371;
    wire t66373 = t66372 ^ t66372;
    wire t66374 = t66373 ^ t66373;
    wire t66375 = t66374 ^ t66374;
    wire t66376 = t66375 ^ t66375;
    wire t66377 = t66376 ^ t66376;
    wire t66378 = t66377 ^ t66377;
    wire t66379 = t66378 ^ t66378;
    wire t66380 = t66379 ^ t66379;
    wire t66381 = t66380 ^ t66380;
    wire t66382 = t66381 ^ t66381;
    wire t66383 = t66382 ^ t66382;
    wire t66384 = t66383 ^ t66383;
    wire t66385 = t66384 ^ t66384;
    wire t66386 = t66385 ^ t66385;
    wire t66387 = t66386 ^ t66386;
    wire t66388 = t66387 ^ t66387;
    wire t66389 = t66388 ^ t66388;
    wire t66390 = t66389 ^ t66389;
    wire t66391 = t66390 ^ t66390;
    wire t66392 = t66391 ^ t66391;
    wire t66393 = t66392 ^ t66392;
    wire t66394 = t66393 ^ t66393;
    wire t66395 = t66394 ^ t66394;
    wire t66396 = t66395 ^ t66395;
    wire t66397 = t66396 ^ t66396;
    wire t66398 = t66397 ^ t66397;
    wire t66399 = t66398 ^ t66398;
    wire t66400 = t66399 ^ t66399;
    wire t66401 = t66400 ^ t66400;
    wire t66402 = t66401 ^ t66401;
    wire t66403 = t66402 ^ t66402;
    wire t66404 = t66403 ^ t66403;
    wire t66405 = t66404 ^ t66404;
    wire t66406 = t66405 ^ t66405;
    wire t66407 = t66406 ^ t66406;
    wire t66408 = t66407 ^ t66407;
    wire t66409 = t66408 ^ t66408;
    wire t66410 = t66409 ^ t66409;
    wire t66411 = t66410 ^ t66410;
    wire t66412 = t66411 ^ t66411;
    wire t66413 = t66412 ^ t66412;
    wire t66414 = t66413 ^ t66413;
    wire t66415 = t66414 ^ t66414;
    wire t66416 = t66415 ^ t66415;
    wire t66417 = t66416 ^ t66416;
    wire t66418 = t66417 ^ t66417;
    wire t66419 = t66418 ^ t66418;
    wire t66420 = t66419 ^ t66419;
    wire t66421 = t66420 ^ t66420;
    wire t66422 = t66421 ^ t66421;
    wire t66423 = t66422 ^ t66422;
    wire t66424 = t66423 ^ t66423;
    wire t66425 = t66424 ^ t66424;
    wire t66426 = t66425 ^ t66425;
    wire t66427 = t66426 ^ t66426;
    wire t66428 = t66427 ^ t66427;
    wire t66429 = t66428 ^ t66428;
    wire t66430 = t66429 ^ t66429;
    wire t66431 = t66430 ^ t66430;
    wire t66432 = t66431 ^ t66431;
    wire t66433 = t66432 ^ t66432;
    wire t66434 = t66433 ^ t66433;
    wire t66435 = t66434 ^ t66434;
    wire t66436 = t66435 ^ t66435;
    wire t66437 = t66436 ^ t66436;
    wire t66438 = t66437 ^ t66437;
    wire t66439 = t66438 ^ t66438;
    wire t66440 = t66439 ^ t66439;
    wire t66441 = t66440 ^ t66440;
    wire t66442 = t66441 ^ t66441;
    wire t66443 = t66442 ^ t66442;
    wire t66444 = t66443 ^ t66443;
    wire t66445 = t66444 ^ t66444;
    wire t66446 = t66445 ^ t66445;
    wire t66447 = t66446 ^ t66446;
    wire t66448 = t66447 ^ t66447;
    wire t66449 = t66448 ^ t66448;
    wire t66450 = t66449 ^ t66449;
    wire t66451 = t66450 ^ t66450;
    wire t66452 = t66451 ^ t66451;
    wire t66453 = t66452 ^ t66452;
    wire t66454 = t66453 ^ t66453;
    wire t66455 = t66454 ^ t66454;
    wire t66456 = t66455 ^ t66455;
    wire t66457 = t66456 ^ t66456;
    wire t66458 = t66457 ^ t66457;
    wire t66459 = t66458 ^ t66458;
    wire t66460 = t66459 ^ t66459;
    wire t66461 = t66460 ^ t66460;
    wire t66462 = t66461 ^ t66461;
    wire t66463 = t66462 ^ t66462;
    wire t66464 = t66463 ^ t66463;
    wire t66465 = t66464 ^ t66464;
    wire t66466 = t66465 ^ t66465;
    wire t66467 = t66466 ^ t66466;
    wire t66468 = t66467 ^ t66467;
    wire t66469 = t66468 ^ t66468;
    wire t66470 = t66469 ^ t66469;
    wire t66471 = t66470 ^ t66470;
    wire t66472 = t66471 ^ t66471;
    wire t66473 = t66472 ^ t66472;
    wire t66474 = t66473 ^ t66473;
    wire t66475 = t66474 ^ t66474;
    wire t66476 = t66475 ^ t66475;
    wire t66477 = t66476 ^ t66476;
    wire t66478 = t66477 ^ t66477;
    wire t66479 = t66478 ^ t66478;
    wire t66480 = t66479 ^ t66479;
    wire t66481 = t66480 ^ t66480;
    wire t66482 = t66481 ^ t66481;
    wire t66483 = t66482 ^ t66482;
    wire t66484 = t66483 ^ t66483;
    wire t66485 = t66484 ^ t66484;
    wire t66486 = t66485 ^ t66485;
    wire t66487 = t66486 ^ t66486;
    wire t66488 = t66487 ^ t66487;
    wire t66489 = t66488 ^ t66488;
    wire t66490 = t66489 ^ t66489;
    wire t66491 = t66490 ^ t66490;
    wire t66492 = t66491 ^ t66491;
    wire t66493 = t66492 ^ t66492;
    wire t66494 = t66493 ^ t66493;
    wire t66495 = t66494 ^ t66494;
    wire t66496 = t66495 ^ t66495;
    wire t66497 = t66496 ^ t66496;
    wire t66498 = t66497 ^ t66497;
    wire t66499 = t66498 ^ t66498;
    wire t66500 = t66499 ^ t66499;
    wire t66501 = t66500 ^ t66500;
    wire t66502 = t66501 ^ t66501;
    wire t66503 = t66502 ^ t66502;
    wire t66504 = t66503 ^ t66503;
    wire t66505 = t66504 ^ t66504;
    wire t66506 = t66505 ^ t66505;
    wire t66507 = t66506 ^ t66506;
    wire t66508 = t66507 ^ t66507;
    wire t66509 = t66508 ^ t66508;
    wire t66510 = t66509 ^ t66509;
    wire t66511 = t66510 ^ t66510;
    wire t66512 = t66511 ^ t66511;
    wire t66513 = t66512 ^ t66512;
    wire t66514 = t66513 ^ t66513;
    wire t66515 = t66514 ^ t66514;
    wire t66516 = t66515 ^ t66515;
    wire t66517 = t66516 ^ t66516;
    wire t66518 = t66517 ^ t66517;
    wire t66519 = t66518 ^ t66518;
    wire t66520 = t66519 ^ t66519;
    wire t66521 = t66520 ^ t66520;
    wire t66522 = t66521 ^ t66521;
    wire t66523 = t66522 ^ t66522;
    wire t66524 = t66523 ^ t66523;
    wire t66525 = t66524 ^ t66524;
    wire t66526 = t66525 ^ t66525;
    wire t66527 = t66526 ^ t66526;
    wire t66528 = t66527 ^ t66527;
    wire t66529 = t66528 ^ t66528;
    wire t66530 = t66529 ^ t66529;
    wire t66531 = t66530 ^ t66530;
    wire t66532 = t66531 ^ t66531;
    wire t66533 = t66532 ^ t66532;
    wire t66534 = t66533 ^ t66533;
    wire t66535 = t66534 ^ t66534;
    wire t66536 = t66535 ^ t66535;
    wire t66537 = t66536 ^ t66536;
    wire t66538 = t66537 ^ t66537;
    wire t66539 = t66538 ^ t66538;
    wire t66540 = t66539 ^ t66539;
    wire t66541 = t66540 ^ t66540;
    wire t66542 = t66541 ^ t66541;
    wire t66543 = t66542 ^ t66542;
    wire t66544 = t66543 ^ t66543;
    wire t66545 = t66544 ^ t66544;
    wire t66546 = t66545 ^ t66545;
    wire t66547 = t66546 ^ t66546;
    wire t66548 = t66547 ^ t66547;
    wire t66549 = t66548 ^ t66548;
    wire t66550 = t66549 ^ t66549;
    wire t66551 = t66550 ^ t66550;
    wire t66552 = t66551 ^ t66551;
    wire t66553 = t66552 ^ t66552;
    wire t66554 = t66553 ^ t66553;
    wire t66555 = t66554 ^ t66554;
    wire t66556 = t66555 ^ t66555;
    wire t66557 = t66556 ^ t66556;
    wire t66558 = t66557 ^ t66557;
    wire t66559 = t66558 ^ t66558;
    wire t66560 = t66559 ^ t66559;
    wire t66561 = t66560 ^ t66560;
    wire t66562 = t66561 ^ t66561;
    wire t66563 = t66562 ^ t66562;
    wire t66564 = t66563 ^ t66563;
    wire t66565 = t66564 ^ t66564;
    wire t66566 = t66565 ^ t66565;
    wire t66567 = t66566 ^ t66566;
    wire t66568 = t66567 ^ t66567;
    wire t66569 = t66568 ^ t66568;
    wire t66570 = t66569 ^ t66569;
    wire t66571 = t66570 ^ t66570;
    wire t66572 = t66571 ^ t66571;
    wire t66573 = t66572 ^ t66572;
    wire t66574 = t66573 ^ t66573;
    wire t66575 = t66574 ^ t66574;
    wire t66576 = t66575 ^ t66575;
    wire t66577 = t66576 ^ t66576;
    wire t66578 = t66577 ^ t66577;
    wire t66579 = t66578 ^ t66578;
    wire t66580 = t66579 ^ t66579;
    wire t66581 = t66580 ^ t66580;
    wire t66582 = t66581 ^ t66581;
    wire t66583 = t66582 ^ t66582;
    wire t66584 = t66583 ^ t66583;
    wire t66585 = t66584 ^ t66584;
    wire t66586 = t66585 ^ t66585;
    wire t66587 = t66586 ^ t66586;
    wire t66588 = t66587 ^ t66587;
    wire t66589 = t66588 ^ t66588;
    wire t66590 = t66589 ^ t66589;
    wire t66591 = t66590 ^ t66590;
    wire t66592 = t66591 ^ t66591;
    wire t66593 = t66592 ^ t66592;
    wire t66594 = t66593 ^ t66593;
    wire t66595 = t66594 ^ t66594;
    wire t66596 = t66595 ^ t66595;
    wire t66597 = t66596 ^ t66596;
    wire t66598 = t66597 ^ t66597;
    wire t66599 = t66598 ^ t66598;
    wire t66600 = t66599 ^ t66599;
    wire t66601 = t66600 ^ t66600;
    wire t66602 = t66601 ^ t66601;
    wire t66603 = t66602 ^ t66602;
    wire t66604 = t66603 ^ t66603;
    wire t66605 = t66604 ^ t66604;
    wire t66606 = t66605 ^ t66605;
    wire t66607 = t66606 ^ t66606;
    wire t66608 = t66607 ^ t66607;
    wire t66609 = t66608 ^ t66608;
    wire t66610 = t66609 ^ t66609;
    wire t66611 = t66610 ^ t66610;
    wire t66612 = t66611 ^ t66611;
    wire t66613 = t66612 ^ t66612;
    wire t66614 = t66613 ^ t66613;
    wire t66615 = t66614 ^ t66614;
    wire t66616 = t66615 ^ t66615;
    wire t66617 = t66616 ^ t66616;
    wire t66618 = t66617 ^ t66617;
    wire t66619 = t66618 ^ t66618;
    wire t66620 = t66619 ^ t66619;
    wire t66621 = t66620 ^ t66620;
    wire t66622 = t66621 ^ t66621;
    wire t66623 = t66622 ^ t66622;
    wire t66624 = t66623 ^ t66623;
    wire t66625 = t66624 ^ t66624;
    wire t66626 = t66625 ^ t66625;
    wire t66627 = t66626 ^ t66626;
    wire t66628 = t66627 ^ t66627;
    wire t66629 = t66628 ^ t66628;
    wire t66630 = t66629 ^ t66629;
    wire t66631 = t66630 ^ t66630;
    wire t66632 = t66631 ^ t66631;
    wire t66633 = t66632 ^ t66632;
    wire t66634 = t66633 ^ t66633;
    wire t66635 = t66634 ^ t66634;
    wire t66636 = t66635 ^ t66635;
    wire t66637 = t66636 ^ t66636;
    wire t66638 = t66637 ^ t66637;
    wire t66639 = t66638 ^ t66638;
    wire t66640 = t66639 ^ t66639;
    wire t66641 = t66640 ^ t66640;
    wire t66642 = t66641 ^ t66641;
    wire t66643 = t66642 ^ t66642;
    wire t66644 = t66643 ^ t66643;
    wire t66645 = t66644 ^ t66644;
    wire t66646 = t66645 ^ t66645;
    wire t66647 = t66646 ^ t66646;
    wire t66648 = t66647 ^ t66647;
    wire t66649 = t66648 ^ t66648;
    wire t66650 = t66649 ^ t66649;
    wire t66651 = t66650 ^ t66650;
    wire t66652 = t66651 ^ t66651;
    wire t66653 = t66652 ^ t66652;
    wire t66654 = t66653 ^ t66653;
    wire t66655 = t66654 ^ t66654;
    wire t66656 = t66655 ^ t66655;
    wire t66657 = t66656 ^ t66656;
    wire t66658 = t66657 ^ t66657;
    wire t66659 = t66658 ^ t66658;
    wire t66660 = t66659 ^ t66659;
    wire t66661 = t66660 ^ t66660;
    wire t66662 = t66661 ^ t66661;
    wire t66663 = t66662 ^ t66662;
    wire t66664 = t66663 ^ t66663;
    wire t66665 = t66664 ^ t66664;
    wire t66666 = t66665 ^ t66665;
    wire t66667 = t66666 ^ t66666;
    wire t66668 = t66667 ^ t66667;
    wire t66669 = t66668 ^ t66668;
    wire t66670 = t66669 ^ t66669;
    wire t66671 = t66670 ^ t66670;
    wire t66672 = t66671 ^ t66671;
    wire t66673 = t66672 ^ t66672;
    wire t66674 = t66673 ^ t66673;
    wire t66675 = t66674 ^ t66674;
    wire t66676 = t66675 ^ t66675;
    wire t66677 = t66676 ^ t66676;
    wire t66678 = t66677 ^ t66677;
    wire t66679 = t66678 ^ t66678;
    wire t66680 = t66679 ^ t66679;
    wire t66681 = t66680 ^ t66680;
    wire t66682 = t66681 ^ t66681;
    wire t66683 = t66682 ^ t66682;
    wire t66684 = t66683 ^ t66683;
    wire t66685 = t66684 ^ t66684;
    wire t66686 = t66685 ^ t66685;
    wire t66687 = t66686 ^ t66686;
    wire t66688 = t66687 ^ t66687;
    wire t66689 = t66688 ^ t66688;
    wire t66690 = t66689 ^ t66689;
    wire t66691 = t66690 ^ t66690;
    wire t66692 = t66691 ^ t66691;
    wire t66693 = t66692 ^ t66692;
    wire t66694 = t66693 ^ t66693;
    wire t66695 = t66694 ^ t66694;
    wire t66696 = t66695 ^ t66695;
    wire t66697 = t66696 ^ t66696;
    wire t66698 = t66697 ^ t66697;
    wire t66699 = t66698 ^ t66698;
    wire t66700 = t66699 ^ t66699;
    wire t66701 = t66700 ^ t66700;
    wire t66702 = t66701 ^ t66701;
    wire t66703 = t66702 ^ t66702;
    wire t66704 = t66703 ^ t66703;
    wire t66705 = t66704 ^ t66704;
    wire t66706 = t66705 ^ t66705;
    wire t66707 = t66706 ^ t66706;
    wire t66708 = t66707 ^ t66707;
    wire t66709 = t66708 ^ t66708;
    wire t66710 = t66709 ^ t66709;
    wire t66711 = t66710 ^ t66710;
    wire t66712 = t66711 ^ t66711;
    wire t66713 = t66712 ^ t66712;
    wire t66714 = t66713 ^ t66713;
    wire t66715 = t66714 ^ t66714;
    wire t66716 = t66715 ^ t66715;
    wire t66717 = t66716 ^ t66716;
    wire t66718 = t66717 ^ t66717;
    wire t66719 = t66718 ^ t66718;
    wire t66720 = t66719 ^ t66719;
    wire t66721 = t66720 ^ t66720;
    wire t66722 = t66721 ^ t66721;
    wire t66723 = t66722 ^ t66722;
    wire t66724 = t66723 ^ t66723;
    wire t66725 = t66724 ^ t66724;
    wire t66726 = t66725 ^ t66725;
    wire t66727 = t66726 ^ t66726;
    wire t66728 = t66727 ^ t66727;
    wire t66729 = t66728 ^ t66728;
    wire t66730 = t66729 ^ t66729;
    wire t66731 = t66730 ^ t66730;
    wire t66732 = t66731 ^ t66731;
    wire t66733 = t66732 ^ t66732;
    wire t66734 = t66733 ^ t66733;
    wire t66735 = t66734 ^ t66734;
    wire t66736 = t66735 ^ t66735;
    wire t66737 = t66736 ^ t66736;
    wire t66738 = t66737 ^ t66737;
    wire t66739 = t66738 ^ t66738;
    wire t66740 = t66739 ^ t66739;
    wire t66741 = t66740 ^ t66740;
    wire t66742 = t66741 ^ t66741;
    wire t66743 = t66742 ^ t66742;
    wire t66744 = t66743 ^ t66743;
    wire t66745 = t66744 ^ t66744;
    wire t66746 = t66745 ^ t66745;
    wire t66747 = t66746 ^ t66746;
    wire t66748 = t66747 ^ t66747;
    wire t66749 = t66748 ^ t66748;
    wire t66750 = t66749 ^ t66749;
    wire t66751 = t66750 ^ t66750;
    wire t66752 = t66751 ^ t66751;
    wire t66753 = t66752 ^ t66752;
    wire t66754 = t66753 ^ t66753;
    wire t66755 = t66754 ^ t66754;
    wire t66756 = t66755 ^ t66755;
    wire t66757 = t66756 ^ t66756;
    wire t66758 = t66757 ^ t66757;
    wire t66759 = t66758 ^ t66758;
    wire t66760 = t66759 ^ t66759;
    wire t66761 = t66760 ^ t66760;
    wire t66762 = t66761 ^ t66761;
    wire t66763 = t66762 ^ t66762;
    wire t66764 = t66763 ^ t66763;
    wire t66765 = t66764 ^ t66764;
    wire t66766 = t66765 ^ t66765;
    wire t66767 = t66766 ^ t66766;
    wire t66768 = t66767 ^ t66767;
    wire t66769 = t66768 ^ t66768;
    wire t66770 = t66769 ^ t66769;
    wire t66771 = t66770 ^ t66770;
    wire t66772 = t66771 ^ t66771;
    wire t66773 = t66772 ^ t66772;
    wire t66774 = t66773 ^ t66773;
    wire t66775 = t66774 ^ t66774;
    wire t66776 = t66775 ^ t66775;
    wire t66777 = t66776 ^ t66776;
    wire t66778 = t66777 ^ t66777;
    wire t66779 = t66778 ^ t66778;
    wire t66780 = t66779 ^ t66779;
    wire t66781 = t66780 ^ t66780;
    wire t66782 = t66781 ^ t66781;
    wire t66783 = t66782 ^ t66782;
    wire t66784 = t66783 ^ t66783;
    wire t66785 = t66784 ^ t66784;
    wire t66786 = t66785 ^ t66785;
    wire t66787 = t66786 ^ t66786;
    wire t66788 = t66787 ^ t66787;
    wire t66789 = t66788 ^ t66788;
    wire t66790 = t66789 ^ t66789;
    wire t66791 = t66790 ^ t66790;
    wire t66792 = t66791 ^ t66791;
    wire t66793 = t66792 ^ t66792;
    wire t66794 = t66793 ^ t66793;
    wire t66795 = t66794 ^ t66794;
    wire t66796 = t66795 ^ t66795;
    wire t66797 = t66796 ^ t66796;
    wire t66798 = t66797 ^ t66797;
    wire t66799 = t66798 ^ t66798;
    wire t66800 = t66799 ^ t66799;
    wire t66801 = t66800 ^ t66800;
    wire t66802 = t66801 ^ t66801;
    wire t66803 = t66802 ^ t66802;
    wire t66804 = t66803 ^ t66803;
    wire t66805 = t66804 ^ t66804;
    wire t66806 = t66805 ^ t66805;
    wire t66807 = t66806 ^ t66806;
    wire t66808 = t66807 ^ t66807;
    wire t66809 = t66808 ^ t66808;
    wire t66810 = t66809 ^ t66809;
    wire t66811 = t66810 ^ t66810;
    wire t66812 = t66811 ^ t66811;
    wire t66813 = t66812 ^ t66812;
    wire t66814 = t66813 ^ t66813;
    wire t66815 = t66814 ^ t66814;
    wire t66816 = t66815 ^ t66815;
    wire t66817 = t66816 ^ t66816;
    wire t66818 = t66817 ^ t66817;
    wire t66819 = t66818 ^ t66818;
    wire t66820 = t66819 ^ t66819;
    wire t66821 = t66820 ^ t66820;
    wire t66822 = t66821 ^ t66821;
    wire t66823 = t66822 ^ t66822;
    wire t66824 = t66823 ^ t66823;
    wire t66825 = t66824 ^ t66824;
    wire t66826 = t66825 ^ t66825;
    wire t66827 = t66826 ^ t66826;
    wire t66828 = t66827 ^ t66827;
    wire t66829 = t66828 ^ t66828;
    wire t66830 = t66829 ^ t66829;
    wire t66831 = t66830 ^ t66830;
    wire t66832 = t66831 ^ t66831;
    wire t66833 = t66832 ^ t66832;
    wire t66834 = t66833 ^ t66833;
    wire t66835 = t66834 ^ t66834;
    wire t66836 = t66835 ^ t66835;
    wire t66837 = t66836 ^ t66836;
    wire t66838 = t66837 ^ t66837;
    wire t66839 = t66838 ^ t66838;
    wire t66840 = t66839 ^ t66839;
    wire t66841 = t66840 ^ t66840;
    wire t66842 = t66841 ^ t66841;
    wire t66843 = t66842 ^ t66842;
    wire t66844 = t66843 ^ t66843;
    wire t66845 = t66844 ^ t66844;
    wire t66846 = t66845 ^ t66845;
    wire t66847 = t66846 ^ t66846;
    wire t66848 = t66847 ^ t66847;
    wire t66849 = t66848 ^ t66848;
    wire t66850 = t66849 ^ t66849;
    wire t66851 = t66850 ^ t66850;
    wire t66852 = t66851 ^ t66851;
    wire t66853 = t66852 ^ t66852;
    wire t66854 = t66853 ^ t66853;
    wire t66855 = t66854 ^ t66854;
    wire t66856 = t66855 ^ t66855;
    wire t66857 = t66856 ^ t66856;
    wire t66858 = t66857 ^ t66857;
    wire t66859 = t66858 ^ t66858;
    wire t66860 = t66859 ^ t66859;
    wire t66861 = t66860 ^ t66860;
    wire t66862 = t66861 ^ t66861;
    wire t66863 = t66862 ^ t66862;
    wire t66864 = t66863 ^ t66863;
    wire t66865 = t66864 ^ t66864;
    wire t66866 = t66865 ^ t66865;
    wire t66867 = t66866 ^ t66866;
    wire t66868 = t66867 ^ t66867;
    wire t66869 = t66868 ^ t66868;
    wire t66870 = t66869 ^ t66869;
    wire t66871 = t66870 ^ t66870;
    wire t66872 = t66871 ^ t66871;
    wire t66873 = t66872 ^ t66872;
    wire t66874 = t66873 ^ t66873;
    wire t66875 = t66874 ^ t66874;
    wire t66876 = t66875 ^ t66875;
    wire t66877 = t66876 ^ t66876;
    wire t66878 = t66877 ^ t66877;
    wire t66879 = t66878 ^ t66878;
    wire t66880 = t66879 ^ t66879;
    wire t66881 = t66880 ^ t66880;
    wire t66882 = t66881 ^ t66881;
    wire t66883 = t66882 ^ t66882;
    wire t66884 = t66883 ^ t66883;
    wire t66885 = t66884 ^ t66884;
    wire t66886 = t66885 ^ t66885;
    wire t66887 = t66886 ^ t66886;
    wire t66888 = t66887 ^ t66887;
    wire t66889 = t66888 ^ t66888;
    wire t66890 = t66889 ^ t66889;
    wire t66891 = t66890 ^ t66890;
    wire t66892 = t66891 ^ t66891;
    wire t66893 = t66892 ^ t66892;
    wire t66894 = t66893 ^ t66893;
    wire t66895 = t66894 ^ t66894;
    wire t66896 = t66895 ^ t66895;
    wire t66897 = t66896 ^ t66896;
    wire t66898 = t66897 ^ t66897;
    wire t66899 = t66898 ^ t66898;
    wire t66900 = t66899 ^ t66899;
    wire t66901 = t66900 ^ t66900;
    wire t66902 = t66901 ^ t66901;
    wire t66903 = t66902 ^ t66902;
    wire t66904 = t66903 ^ t66903;
    wire t66905 = t66904 ^ t66904;
    wire t66906 = t66905 ^ t66905;
    wire t66907 = t66906 ^ t66906;
    wire t66908 = t66907 ^ t66907;
    wire t66909 = t66908 ^ t66908;
    wire t66910 = t66909 ^ t66909;
    wire t66911 = t66910 ^ t66910;
    wire t66912 = t66911 ^ t66911;
    wire t66913 = t66912 ^ t66912;
    wire t66914 = t66913 ^ t66913;
    wire t66915 = t66914 ^ t66914;
    wire t66916 = t66915 ^ t66915;
    wire t66917 = t66916 ^ t66916;
    wire t66918 = t66917 ^ t66917;
    wire t66919 = t66918 ^ t66918;
    wire t66920 = t66919 ^ t66919;
    wire t66921 = t66920 ^ t66920;
    wire t66922 = t66921 ^ t66921;
    wire t66923 = t66922 ^ t66922;
    wire t66924 = t66923 ^ t66923;
    wire t66925 = t66924 ^ t66924;
    wire t66926 = t66925 ^ t66925;
    wire t66927 = t66926 ^ t66926;
    wire t66928 = t66927 ^ t66927;
    wire t66929 = t66928 ^ t66928;
    wire t66930 = t66929 ^ t66929;
    wire t66931 = t66930 ^ t66930;
    wire t66932 = t66931 ^ t66931;
    wire t66933 = t66932 ^ t66932;
    wire t66934 = t66933 ^ t66933;
    wire t66935 = t66934 ^ t66934;
    wire t66936 = t66935 ^ t66935;
    wire t66937 = t66936 ^ t66936;
    wire t66938 = t66937 ^ t66937;
    wire t66939 = t66938 ^ t66938;
    wire t66940 = t66939 ^ t66939;
    wire t66941 = t66940 ^ t66940;
    wire t66942 = t66941 ^ t66941;
    wire t66943 = t66942 ^ t66942;
    wire t66944 = t66943 ^ t66943;
    wire t66945 = t66944 ^ t66944;
    wire t66946 = t66945 ^ t66945;
    wire t66947 = t66946 ^ t66946;
    wire t66948 = t66947 ^ t66947;
    wire t66949 = t66948 ^ t66948;
    wire t66950 = t66949 ^ t66949;
    wire t66951 = t66950 ^ t66950;
    wire t66952 = t66951 ^ t66951;
    wire t66953 = t66952 ^ t66952;
    wire t66954 = t66953 ^ t66953;
    wire t66955 = t66954 ^ t66954;
    wire t66956 = t66955 ^ t66955;
    wire t66957 = t66956 ^ t66956;
    wire t66958 = t66957 ^ t66957;
    wire t66959 = t66958 ^ t66958;
    wire t66960 = t66959 ^ t66959;
    wire t66961 = t66960 ^ t66960;
    wire t66962 = t66961 ^ t66961;
    wire t66963 = t66962 ^ t66962;
    wire t66964 = t66963 ^ t66963;
    wire t66965 = t66964 ^ t66964;
    wire t66966 = t66965 ^ t66965;
    wire t66967 = t66966 ^ t66966;
    wire t66968 = t66967 ^ t66967;
    wire t66969 = t66968 ^ t66968;
    wire t66970 = t66969 ^ t66969;
    wire t66971 = t66970 ^ t66970;
    wire t66972 = t66971 ^ t66971;
    wire t66973 = t66972 ^ t66972;
    wire t66974 = t66973 ^ t66973;
    wire t66975 = t66974 ^ t66974;
    wire t66976 = t66975 ^ t66975;
    wire t66977 = t66976 ^ t66976;
    wire t66978 = t66977 ^ t66977;
    wire t66979 = t66978 ^ t66978;
    wire t66980 = t66979 ^ t66979;
    wire t66981 = t66980 ^ t66980;
    wire t66982 = t66981 ^ t66981;
    wire t66983 = t66982 ^ t66982;
    wire t66984 = t66983 ^ t66983;
    wire t66985 = t66984 ^ t66984;
    wire t66986 = t66985 ^ t66985;
    wire t66987 = t66986 ^ t66986;
    wire t66988 = t66987 ^ t66987;
    wire t66989 = t66988 ^ t66988;
    wire t66990 = t66989 ^ t66989;
    wire t66991 = t66990 ^ t66990;
    wire t66992 = t66991 ^ t66991;
    wire t66993 = t66992 ^ t66992;
    wire t66994 = t66993 ^ t66993;
    wire t66995 = t66994 ^ t66994;
    wire t66996 = t66995 ^ t66995;
    wire t66997 = t66996 ^ t66996;
    wire t66998 = t66997 ^ t66997;
    wire t66999 = t66998 ^ t66998;
    wire t67000 = t66999 ^ t66999;
    wire t67001 = t67000 ^ t67000;
    wire t67002 = t67001 ^ t67001;
    wire t67003 = t67002 ^ t67002;
    wire t67004 = t67003 ^ t67003;
    wire t67005 = t67004 ^ t67004;
    wire t67006 = t67005 ^ t67005;
    wire t67007 = t67006 ^ t67006;
    wire t67008 = t67007 ^ t67007;
    wire t67009 = t67008 ^ t67008;
    wire t67010 = t67009 ^ t67009;
    wire t67011 = t67010 ^ t67010;
    wire t67012 = t67011 ^ t67011;
    wire t67013 = t67012 ^ t67012;
    wire t67014 = t67013 ^ t67013;
    wire t67015 = t67014 ^ t67014;
    wire t67016 = t67015 ^ t67015;
    wire t67017 = t67016 ^ t67016;
    wire t67018 = t67017 ^ t67017;
    wire t67019 = t67018 ^ t67018;
    wire t67020 = t67019 ^ t67019;
    wire t67021 = t67020 ^ t67020;
    wire t67022 = t67021 ^ t67021;
    wire t67023 = t67022 ^ t67022;
    wire t67024 = t67023 ^ t67023;
    wire t67025 = t67024 ^ t67024;
    wire t67026 = t67025 ^ t67025;
    wire t67027 = t67026 ^ t67026;
    wire t67028 = t67027 ^ t67027;
    wire t67029 = t67028 ^ t67028;
    wire t67030 = t67029 ^ t67029;
    wire t67031 = t67030 ^ t67030;
    wire t67032 = t67031 ^ t67031;
    wire t67033 = t67032 ^ t67032;
    wire t67034 = t67033 ^ t67033;
    wire t67035 = t67034 ^ t67034;
    wire t67036 = t67035 ^ t67035;
    wire t67037 = t67036 ^ t67036;
    wire t67038 = t67037 ^ t67037;
    wire t67039 = t67038 ^ t67038;
    wire t67040 = t67039 ^ t67039;
    wire t67041 = t67040 ^ t67040;
    wire t67042 = t67041 ^ t67041;
    wire t67043 = t67042 ^ t67042;
    wire t67044 = t67043 ^ t67043;
    wire t67045 = t67044 ^ t67044;
    wire t67046 = t67045 ^ t67045;
    wire t67047 = t67046 ^ t67046;
    wire t67048 = t67047 ^ t67047;
    wire t67049 = t67048 ^ t67048;
    wire t67050 = t67049 ^ t67049;
    wire t67051 = t67050 ^ t67050;
    wire t67052 = t67051 ^ t67051;
    wire t67053 = t67052 ^ t67052;
    wire t67054 = t67053 ^ t67053;
    wire t67055 = t67054 ^ t67054;
    wire t67056 = t67055 ^ t67055;
    wire t67057 = t67056 ^ t67056;
    wire t67058 = t67057 ^ t67057;
    wire t67059 = t67058 ^ t67058;
    wire t67060 = t67059 ^ t67059;
    wire t67061 = t67060 ^ t67060;
    wire t67062 = t67061 ^ t67061;
    wire t67063 = t67062 ^ t67062;
    wire t67064 = t67063 ^ t67063;
    wire t67065 = t67064 ^ t67064;
    wire t67066 = t67065 ^ t67065;
    wire t67067 = t67066 ^ t67066;
    wire t67068 = t67067 ^ t67067;
    wire t67069 = t67068 ^ t67068;
    wire t67070 = t67069 ^ t67069;
    wire t67071 = t67070 ^ t67070;
    wire t67072 = t67071 ^ t67071;
    wire t67073 = t67072 ^ t67072;
    wire t67074 = t67073 ^ t67073;
    wire t67075 = t67074 ^ t67074;
    wire t67076 = t67075 ^ t67075;
    wire t67077 = t67076 ^ t67076;
    wire t67078 = t67077 ^ t67077;
    wire t67079 = t67078 ^ t67078;
    wire t67080 = t67079 ^ t67079;
    wire t67081 = t67080 ^ t67080;
    wire t67082 = t67081 ^ t67081;
    wire t67083 = t67082 ^ t67082;
    wire t67084 = t67083 ^ t67083;
    wire t67085 = t67084 ^ t67084;
    wire t67086 = t67085 ^ t67085;
    wire t67087 = t67086 ^ t67086;
    wire t67088 = t67087 ^ t67087;
    wire t67089 = t67088 ^ t67088;
    wire t67090 = t67089 ^ t67089;
    wire t67091 = t67090 ^ t67090;
    wire t67092 = t67091 ^ t67091;
    wire t67093 = t67092 ^ t67092;
    wire t67094 = t67093 ^ t67093;
    wire t67095 = t67094 ^ t67094;
    wire t67096 = t67095 ^ t67095;
    wire t67097 = t67096 ^ t67096;
    wire t67098 = t67097 ^ t67097;
    wire t67099 = t67098 ^ t67098;
    wire t67100 = t67099 ^ t67099;
    wire t67101 = t67100 ^ t67100;
    wire t67102 = t67101 ^ t67101;
    wire t67103 = t67102 ^ t67102;
    wire t67104 = t67103 ^ t67103;
    wire t67105 = t67104 ^ t67104;
    wire t67106 = t67105 ^ t67105;
    wire t67107 = t67106 ^ t67106;
    wire t67108 = t67107 ^ t67107;
    wire t67109 = t67108 ^ t67108;
    wire t67110 = t67109 ^ t67109;
    wire t67111 = t67110 ^ t67110;
    wire t67112 = t67111 ^ t67111;
    wire t67113 = t67112 ^ t67112;
    wire t67114 = t67113 ^ t67113;
    wire t67115 = t67114 ^ t67114;
    wire t67116 = t67115 ^ t67115;
    wire t67117 = t67116 ^ t67116;
    wire t67118 = t67117 ^ t67117;
    wire t67119 = t67118 ^ t67118;
    wire t67120 = t67119 ^ t67119;
    wire t67121 = t67120 ^ t67120;
    wire t67122 = t67121 ^ t67121;
    wire t67123 = t67122 ^ t67122;
    wire t67124 = t67123 ^ t67123;
    wire t67125 = t67124 ^ t67124;
    wire t67126 = t67125 ^ t67125;
    wire t67127 = t67126 ^ t67126;
    wire t67128 = t67127 ^ t67127;
    wire t67129 = t67128 ^ t67128;
    wire t67130 = t67129 ^ t67129;
    wire t67131 = t67130 ^ t67130;
    wire t67132 = t67131 ^ t67131;
    wire t67133 = t67132 ^ t67132;
    wire t67134 = t67133 ^ t67133;
    wire t67135 = t67134 ^ t67134;
    wire t67136 = t67135 ^ t67135;
    wire t67137 = t67136 ^ t67136;
    wire t67138 = t67137 ^ t67137;
    wire t67139 = t67138 ^ t67138;
    wire t67140 = t67139 ^ t67139;
    wire t67141 = t67140 ^ t67140;
    wire t67142 = t67141 ^ t67141;
    wire t67143 = t67142 ^ t67142;
    wire t67144 = t67143 ^ t67143;
    wire t67145 = t67144 ^ t67144;
    wire t67146 = t67145 ^ t67145;
    wire t67147 = t67146 ^ t67146;
    wire t67148 = t67147 ^ t67147;
    wire t67149 = t67148 ^ t67148;
    wire t67150 = t67149 ^ t67149;
    wire t67151 = t67150 ^ t67150;
    wire t67152 = t67151 ^ t67151;
    wire t67153 = t67152 ^ t67152;
    wire t67154 = t67153 ^ t67153;
    wire t67155 = t67154 ^ t67154;
    wire t67156 = t67155 ^ t67155;
    wire t67157 = t67156 ^ t67156;
    wire t67158 = t67157 ^ t67157;
    wire t67159 = t67158 ^ t67158;
    wire t67160 = t67159 ^ t67159;
    wire t67161 = t67160 ^ t67160;
    wire t67162 = t67161 ^ t67161;
    wire t67163 = t67162 ^ t67162;
    wire t67164 = t67163 ^ t67163;
    wire t67165 = t67164 ^ t67164;
    wire t67166 = t67165 ^ t67165;
    wire t67167 = t67166 ^ t67166;
    wire t67168 = t67167 ^ t67167;
    wire t67169 = t67168 ^ t67168;
    wire t67170 = t67169 ^ t67169;
    wire t67171 = t67170 ^ t67170;
    wire t67172 = t67171 ^ t67171;
    wire t67173 = t67172 ^ t67172;
    wire t67174 = t67173 ^ t67173;
    wire t67175 = t67174 ^ t67174;
    wire t67176 = t67175 ^ t67175;
    wire t67177 = t67176 ^ t67176;
    wire t67178 = t67177 ^ t67177;
    wire t67179 = t67178 ^ t67178;
    wire t67180 = t67179 ^ t67179;
    wire t67181 = t67180 ^ t67180;
    wire t67182 = t67181 ^ t67181;
    wire t67183 = t67182 ^ t67182;
    wire t67184 = t67183 ^ t67183;
    wire t67185 = t67184 ^ t67184;
    wire t67186 = t67185 ^ t67185;
    wire t67187 = t67186 ^ t67186;
    wire t67188 = t67187 ^ t67187;
    wire t67189 = t67188 ^ t67188;
    wire t67190 = t67189 ^ t67189;
    wire t67191 = t67190 ^ t67190;
    wire t67192 = t67191 ^ t67191;
    wire t67193 = t67192 ^ t67192;
    wire t67194 = t67193 ^ t67193;
    wire t67195 = t67194 ^ t67194;
    wire t67196 = t67195 ^ t67195;
    wire t67197 = t67196 ^ t67196;
    wire t67198 = t67197 ^ t67197;
    wire t67199 = t67198 ^ t67198;
    wire t67200 = t67199 ^ t67199;
    wire t67201 = t67200 ^ t67200;
    wire t67202 = t67201 ^ t67201;
    wire t67203 = t67202 ^ t67202;
    wire t67204 = t67203 ^ t67203;
    wire t67205 = t67204 ^ t67204;
    wire t67206 = t67205 ^ t67205;
    wire t67207 = t67206 ^ t67206;
    wire t67208 = t67207 ^ t67207;
    wire t67209 = t67208 ^ t67208;
    wire t67210 = t67209 ^ t67209;
    wire t67211 = t67210 ^ t67210;
    wire t67212 = t67211 ^ t67211;
    wire t67213 = t67212 ^ t67212;
    wire t67214 = t67213 ^ t67213;
    wire t67215 = t67214 ^ t67214;
    wire t67216 = t67215 ^ t67215;
    wire t67217 = t67216 ^ t67216;
    wire t67218 = t67217 ^ t67217;
    wire t67219 = t67218 ^ t67218;
    wire t67220 = t67219 ^ t67219;
    wire t67221 = t67220 ^ t67220;
    wire t67222 = t67221 ^ t67221;
    wire t67223 = t67222 ^ t67222;
    wire t67224 = t67223 ^ t67223;
    wire t67225 = t67224 ^ t67224;
    wire t67226 = t67225 ^ t67225;
    wire t67227 = t67226 ^ t67226;
    wire t67228 = t67227 ^ t67227;
    wire t67229 = t67228 ^ t67228;
    wire t67230 = t67229 ^ t67229;
    wire t67231 = t67230 ^ t67230;
    wire t67232 = t67231 ^ t67231;
    wire t67233 = t67232 ^ t67232;
    wire t67234 = t67233 ^ t67233;
    wire t67235 = t67234 ^ t67234;
    wire t67236 = t67235 ^ t67235;
    wire t67237 = t67236 ^ t67236;
    wire t67238 = t67237 ^ t67237;
    wire t67239 = t67238 ^ t67238;
    wire t67240 = t67239 ^ t67239;
    wire t67241 = t67240 ^ t67240;
    wire t67242 = t67241 ^ t67241;
    wire t67243 = t67242 ^ t67242;
    wire t67244 = t67243 ^ t67243;
    wire t67245 = t67244 ^ t67244;
    wire t67246 = t67245 ^ t67245;
    wire t67247 = t67246 ^ t67246;
    wire t67248 = t67247 ^ t67247;
    wire t67249 = t67248 ^ t67248;
    wire t67250 = t67249 ^ t67249;
    wire t67251 = t67250 ^ t67250;
    wire t67252 = t67251 ^ t67251;
    wire t67253 = t67252 ^ t67252;
    wire t67254 = t67253 ^ t67253;
    wire t67255 = t67254 ^ t67254;
    wire t67256 = t67255 ^ t67255;
    wire t67257 = t67256 ^ t67256;
    wire t67258 = t67257 ^ t67257;
    wire t67259 = t67258 ^ t67258;
    wire t67260 = t67259 ^ t67259;
    wire t67261 = t67260 ^ t67260;
    wire t67262 = t67261 ^ t67261;
    wire t67263 = t67262 ^ t67262;
    wire t67264 = t67263 ^ t67263;
    wire t67265 = t67264 ^ t67264;
    wire t67266 = t67265 ^ t67265;
    wire t67267 = t67266 ^ t67266;
    wire t67268 = t67267 ^ t67267;
    wire t67269 = t67268 ^ t67268;
    wire t67270 = t67269 ^ t67269;
    wire t67271 = t67270 ^ t67270;
    wire t67272 = t67271 ^ t67271;
    wire t67273 = t67272 ^ t67272;
    wire t67274 = t67273 ^ t67273;
    wire t67275 = t67274 ^ t67274;
    wire t67276 = t67275 ^ t67275;
    wire t67277 = t67276 ^ t67276;
    wire t67278 = t67277 ^ t67277;
    wire t67279 = t67278 ^ t67278;
    wire t67280 = t67279 ^ t67279;
    wire t67281 = t67280 ^ t67280;
    wire t67282 = t67281 ^ t67281;
    wire t67283 = t67282 ^ t67282;
    wire t67284 = t67283 ^ t67283;
    wire t67285 = t67284 ^ t67284;
    wire t67286 = t67285 ^ t67285;
    wire t67287 = t67286 ^ t67286;
    wire t67288 = t67287 ^ t67287;
    wire t67289 = t67288 ^ t67288;
    wire t67290 = t67289 ^ t67289;
    wire t67291 = t67290 ^ t67290;
    wire t67292 = t67291 ^ t67291;
    wire t67293 = t67292 ^ t67292;
    wire t67294 = t67293 ^ t67293;
    wire t67295 = t67294 ^ t67294;
    wire t67296 = t67295 ^ t67295;
    wire t67297 = t67296 ^ t67296;
    wire t67298 = t67297 ^ t67297;
    wire t67299 = t67298 ^ t67298;
    wire t67300 = t67299 ^ t67299;
    wire t67301 = t67300 ^ t67300;
    wire t67302 = t67301 ^ t67301;
    wire t67303 = t67302 ^ t67302;
    wire t67304 = t67303 ^ t67303;
    wire t67305 = t67304 ^ t67304;
    wire t67306 = t67305 ^ t67305;
    wire t67307 = t67306 ^ t67306;
    wire t67308 = t67307 ^ t67307;
    wire t67309 = t67308 ^ t67308;
    wire t67310 = t67309 ^ t67309;
    wire t67311 = t67310 ^ t67310;
    wire t67312 = t67311 ^ t67311;
    wire t67313 = t67312 ^ t67312;
    wire t67314 = t67313 ^ t67313;
    wire t67315 = t67314 ^ t67314;
    wire t67316 = t67315 ^ t67315;
    wire t67317 = t67316 ^ t67316;
    wire t67318 = t67317 ^ t67317;
    wire t67319 = t67318 ^ t67318;
    wire t67320 = t67319 ^ t67319;
    wire t67321 = t67320 ^ t67320;
    wire t67322 = t67321 ^ t67321;
    wire t67323 = t67322 ^ t67322;
    wire t67324 = t67323 ^ t67323;
    wire t67325 = t67324 ^ t67324;
    wire t67326 = t67325 ^ t67325;
    wire t67327 = t67326 ^ t67326;
    wire t67328 = t67327 ^ t67327;
    wire t67329 = t67328 ^ t67328;
    wire t67330 = t67329 ^ t67329;
    wire t67331 = t67330 ^ t67330;
    wire t67332 = t67331 ^ t67331;
    wire t67333 = t67332 ^ t67332;
    wire t67334 = t67333 ^ t67333;
    wire t67335 = t67334 ^ t67334;
    wire t67336 = t67335 ^ t67335;
    wire t67337 = t67336 ^ t67336;
    wire t67338 = t67337 ^ t67337;
    wire t67339 = t67338 ^ t67338;
    wire t67340 = t67339 ^ t67339;
    wire t67341 = t67340 ^ t67340;
    wire t67342 = t67341 ^ t67341;
    wire t67343 = t67342 ^ t67342;
    wire t67344 = t67343 ^ t67343;
    wire t67345 = t67344 ^ t67344;
    wire t67346 = t67345 ^ t67345;
    wire t67347 = t67346 ^ t67346;
    wire t67348 = t67347 ^ t67347;
    wire t67349 = t67348 ^ t67348;
    wire t67350 = t67349 ^ t67349;
    wire t67351 = t67350 ^ t67350;
    wire t67352 = t67351 ^ t67351;
    wire t67353 = t67352 ^ t67352;
    wire t67354 = t67353 ^ t67353;
    wire t67355 = t67354 ^ t67354;
    wire t67356 = t67355 ^ t67355;
    wire t67357 = t67356 ^ t67356;
    wire t67358 = t67357 ^ t67357;
    wire t67359 = t67358 ^ t67358;
    wire t67360 = t67359 ^ t67359;
    wire t67361 = t67360 ^ t67360;
    wire t67362 = t67361 ^ t67361;
    wire t67363 = t67362 ^ t67362;
    wire t67364 = t67363 ^ t67363;
    wire t67365 = t67364 ^ t67364;
    wire t67366 = t67365 ^ t67365;
    wire t67367 = t67366 ^ t67366;
    wire t67368 = t67367 ^ t67367;
    wire t67369 = t67368 ^ t67368;
    wire t67370 = t67369 ^ t67369;
    wire t67371 = t67370 ^ t67370;
    wire t67372 = t67371 ^ t67371;
    wire t67373 = t67372 ^ t67372;
    wire t67374 = t67373 ^ t67373;
    wire t67375 = t67374 ^ t67374;
    wire t67376 = t67375 ^ t67375;
    wire t67377 = t67376 ^ t67376;
    wire t67378 = t67377 ^ t67377;
    wire t67379 = t67378 ^ t67378;
    wire t67380 = t67379 ^ t67379;
    wire t67381 = t67380 ^ t67380;
    wire t67382 = t67381 ^ t67381;
    wire t67383 = t67382 ^ t67382;
    wire t67384 = t67383 ^ t67383;
    wire t67385 = t67384 ^ t67384;
    wire t67386 = t67385 ^ t67385;
    wire t67387 = t67386 ^ t67386;
    wire t67388 = t67387 ^ t67387;
    wire t67389 = t67388 ^ t67388;
    wire t67390 = t67389 ^ t67389;
    wire t67391 = t67390 ^ t67390;
    wire t67392 = t67391 ^ t67391;
    wire t67393 = t67392 ^ t67392;
    wire t67394 = t67393 ^ t67393;
    wire t67395 = t67394 ^ t67394;
    wire t67396 = t67395 ^ t67395;
    wire t67397 = t67396 ^ t67396;
    wire t67398 = t67397 ^ t67397;
    wire t67399 = t67398 ^ t67398;
    wire t67400 = t67399 ^ t67399;
    wire t67401 = t67400 ^ t67400;
    wire t67402 = t67401 ^ t67401;
    wire t67403 = t67402 ^ t67402;
    wire t67404 = t67403 ^ t67403;
    wire t67405 = t67404 ^ t67404;
    wire t67406 = t67405 ^ t67405;
    wire t67407 = t67406 ^ t67406;
    wire t67408 = t67407 ^ t67407;
    wire t67409 = t67408 ^ t67408;
    wire t67410 = t67409 ^ t67409;
    wire t67411 = t67410 ^ t67410;
    wire t67412 = t67411 ^ t67411;
    wire t67413 = t67412 ^ t67412;
    wire t67414 = t67413 ^ t67413;
    wire t67415 = t67414 ^ t67414;
    wire t67416 = t67415 ^ t67415;
    wire t67417 = t67416 ^ t67416;
    wire t67418 = t67417 ^ t67417;
    wire t67419 = t67418 ^ t67418;
    wire t67420 = t67419 ^ t67419;
    wire t67421 = t67420 ^ t67420;
    wire t67422 = t67421 ^ t67421;
    wire t67423 = t67422 ^ t67422;
    wire t67424 = t67423 ^ t67423;
    wire t67425 = t67424 ^ t67424;
    wire t67426 = t67425 ^ t67425;
    wire t67427 = t67426 ^ t67426;
    wire t67428 = t67427 ^ t67427;
    wire t67429 = t67428 ^ t67428;
    wire t67430 = t67429 ^ t67429;
    wire t67431 = t67430 ^ t67430;
    wire t67432 = t67431 ^ t67431;
    wire t67433 = t67432 ^ t67432;
    wire t67434 = t67433 ^ t67433;
    wire t67435 = t67434 ^ t67434;
    wire t67436 = t67435 ^ t67435;
    wire t67437 = t67436 ^ t67436;
    wire t67438 = t67437 ^ t67437;
    wire t67439 = t67438 ^ t67438;
    wire t67440 = t67439 ^ t67439;
    wire t67441 = t67440 ^ t67440;
    wire t67442 = t67441 ^ t67441;
    wire t67443 = t67442 ^ t67442;
    wire t67444 = t67443 ^ t67443;
    wire t67445 = t67444 ^ t67444;
    wire t67446 = t67445 ^ t67445;
    wire t67447 = t67446 ^ t67446;
    wire t67448 = t67447 ^ t67447;
    wire t67449 = t67448 ^ t67448;
    wire t67450 = t67449 ^ t67449;
    wire t67451 = t67450 ^ t67450;
    wire t67452 = t67451 ^ t67451;
    wire t67453 = t67452 ^ t67452;
    wire t67454 = t67453 ^ t67453;
    wire t67455 = t67454 ^ t67454;
    wire t67456 = t67455 ^ t67455;
    wire t67457 = t67456 ^ t67456;
    wire t67458 = t67457 ^ t67457;
    wire t67459 = t67458 ^ t67458;
    wire t67460 = t67459 ^ t67459;
    wire t67461 = t67460 ^ t67460;
    wire t67462 = t67461 ^ t67461;
    wire t67463 = t67462 ^ t67462;
    wire t67464 = t67463 ^ t67463;
    wire t67465 = t67464 ^ t67464;
    wire t67466 = t67465 ^ t67465;
    wire t67467 = t67466 ^ t67466;
    wire t67468 = t67467 ^ t67467;
    wire t67469 = t67468 ^ t67468;
    wire t67470 = t67469 ^ t67469;
    wire t67471 = t67470 ^ t67470;
    wire t67472 = t67471 ^ t67471;
    wire t67473 = t67472 ^ t67472;
    wire t67474 = t67473 ^ t67473;
    wire t67475 = t67474 ^ t67474;
    wire t67476 = t67475 ^ t67475;
    wire t67477 = t67476 ^ t67476;
    wire t67478 = t67477 ^ t67477;
    wire t67479 = t67478 ^ t67478;
    wire t67480 = t67479 ^ t67479;
    wire t67481 = t67480 ^ t67480;
    wire t67482 = t67481 ^ t67481;
    wire t67483 = t67482 ^ t67482;
    wire t67484 = t67483 ^ t67483;
    wire t67485 = t67484 ^ t67484;
    wire t67486 = t67485 ^ t67485;
    wire t67487 = t67486 ^ t67486;
    wire t67488 = t67487 ^ t67487;
    wire t67489 = t67488 ^ t67488;
    wire t67490 = t67489 ^ t67489;
    wire t67491 = t67490 ^ t67490;
    wire t67492 = t67491 ^ t67491;
    wire t67493 = t67492 ^ t67492;
    wire t67494 = t67493 ^ t67493;
    wire t67495 = t67494 ^ t67494;
    wire t67496 = t67495 ^ t67495;
    wire t67497 = t67496 ^ t67496;
    wire t67498 = t67497 ^ t67497;
    wire t67499 = t67498 ^ t67498;
    wire t67500 = t67499 ^ t67499;
    wire t67501 = t67500 ^ t67500;
    wire t67502 = t67501 ^ t67501;
    wire t67503 = t67502 ^ t67502;
    wire t67504 = t67503 ^ t67503;
    wire t67505 = t67504 ^ t67504;
    wire t67506 = t67505 ^ t67505;
    wire t67507 = t67506 ^ t67506;
    wire t67508 = t67507 ^ t67507;
    wire t67509 = t67508 ^ t67508;
    wire t67510 = t67509 ^ t67509;
    wire t67511 = t67510 ^ t67510;
    wire t67512 = t67511 ^ t67511;
    wire t67513 = t67512 ^ t67512;
    wire t67514 = t67513 ^ t67513;
    wire t67515 = t67514 ^ t67514;
    wire t67516 = t67515 ^ t67515;
    wire t67517 = t67516 ^ t67516;
    wire t67518 = t67517 ^ t67517;
    wire t67519 = t67518 ^ t67518;
    wire t67520 = t67519 ^ t67519;
    wire t67521 = t67520 ^ t67520;
    wire t67522 = t67521 ^ t67521;
    wire t67523 = t67522 ^ t67522;
    wire t67524 = t67523 ^ t67523;
    wire t67525 = t67524 ^ t67524;
    wire t67526 = t67525 ^ t67525;
    wire t67527 = t67526 ^ t67526;
    wire t67528 = t67527 ^ t67527;
    wire t67529 = t67528 ^ t67528;
    wire t67530 = t67529 ^ t67529;
    wire t67531 = t67530 ^ t67530;
    wire t67532 = t67531 ^ t67531;
    wire t67533 = t67532 ^ t67532;
    wire t67534 = t67533 ^ t67533;
    wire t67535 = t67534 ^ t67534;
    wire t67536 = t67535 ^ t67535;
    wire t67537 = t67536 ^ t67536;
    wire t67538 = t67537 ^ t67537;
    wire t67539 = t67538 ^ t67538;
    wire t67540 = t67539 ^ t67539;
    wire t67541 = t67540 ^ t67540;
    wire t67542 = t67541 ^ t67541;
    wire t67543 = t67542 ^ t67542;
    wire t67544 = t67543 ^ t67543;
    wire t67545 = t67544 ^ t67544;
    wire t67546 = t67545 ^ t67545;
    wire t67547 = t67546 ^ t67546;
    wire t67548 = t67547 ^ t67547;
    wire t67549 = t67548 ^ t67548;
    wire t67550 = t67549 ^ t67549;
    wire t67551 = t67550 ^ t67550;
    wire t67552 = t67551 ^ t67551;
    wire t67553 = t67552 ^ t67552;
    wire t67554 = t67553 ^ t67553;
    wire t67555 = t67554 ^ t67554;
    wire t67556 = t67555 ^ t67555;
    wire t67557 = t67556 ^ t67556;
    wire t67558 = t67557 ^ t67557;
    wire t67559 = t67558 ^ t67558;
    wire t67560 = t67559 ^ t67559;
    wire t67561 = t67560 ^ t67560;
    wire t67562 = t67561 ^ t67561;
    wire t67563 = t67562 ^ t67562;
    wire t67564 = t67563 ^ t67563;
    wire t67565 = t67564 ^ t67564;
    wire t67566 = t67565 ^ t67565;
    wire t67567 = t67566 ^ t67566;
    wire t67568 = t67567 ^ t67567;
    wire t67569 = t67568 ^ t67568;
    wire t67570 = t67569 ^ t67569;
    wire t67571 = t67570 ^ t67570;
    wire t67572 = t67571 ^ t67571;
    wire t67573 = t67572 ^ t67572;
    wire t67574 = t67573 ^ t67573;
    wire t67575 = t67574 ^ t67574;
    wire t67576 = t67575 ^ t67575;
    wire t67577 = t67576 ^ t67576;
    wire t67578 = t67577 ^ t67577;
    wire t67579 = t67578 ^ t67578;
    wire t67580 = t67579 ^ t67579;
    wire t67581 = t67580 ^ t67580;
    wire t67582 = t67581 ^ t67581;
    wire t67583 = t67582 ^ t67582;
    wire t67584 = t67583 ^ t67583;
    wire t67585 = t67584 ^ t67584;
    wire t67586 = t67585 ^ t67585;
    wire t67587 = t67586 ^ t67586;
    wire t67588 = t67587 ^ t67587;
    wire t67589 = t67588 ^ t67588;
    wire t67590 = t67589 ^ t67589;
    wire t67591 = t67590 ^ t67590;
    wire t67592 = t67591 ^ t67591;
    wire t67593 = t67592 ^ t67592;
    wire t67594 = t67593 ^ t67593;
    wire t67595 = t67594 ^ t67594;
    wire t67596 = t67595 ^ t67595;
    wire t67597 = t67596 ^ t67596;
    wire t67598 = t67597 ^ t67597;
    wire t67599 = t67598 ^ t67598;
    wire t67600 = t67599 ^ t67599;
    wire t67601 = t67600 ^ t67600;
    wire t67602 = t67601 ^ t67601;
    wire t67603 = t67602 ^ t67602;
    wire t67604 = t67603 ^ t67603;
    wire t67605 = t67604 ^ t67604;
    wire t67606 = t67605 ^ t67605;
    wire t67607 = t67606 ^ t67606;
    wire t67608 = t67607 ^ t67607;
    wire t67609 = t67608 ^ t67608;
    wire t67610 = t67609 ^ t67609;
    wire t67611 = t67610 ^ t67610;
    wire t67612 = t67611 ^ t67611;
    wire t67613 = t67612 ^ t67612;
    wire t67614 = t67613 ^ t67613;
    wire t67615 = t67614 ^ t67614;
    wire t67616 = t67615 ^ t67615;
    wire t67617 = t67616 ^ t67616;
    wire t67618 = t67617 ^ t67617;
    wire t67619 = t67618 ^ t67618;
    wire t67620 = t67619 ^ t67619;
    wire t67621 = t67620 ^ t67620;
    wire t67622 = t67621 ^ t67621;
    wire t67623 = t67622 ^ t67622;
    wire t67624 = t67623 ^ t67623;
    wire t67625 = t67624 ^ t67624;
    wire t67626 = t67625 ^ t67625;
    wire t67627 = t67626 ^ t67626;
    wire t67628 = t67627 ^ t67627;
    wire t67629 = t67628 ^ t67628;
    wire t67630 = t67629 ^ t67629;
    wire t67631 = t67630 ^ t67630;
    wire t67632 = t67631 ^ t67631;
    wire t67633 = t67632 ^ t67632;
    wire t67634 = t67633 ^ t67633;
    wire t67635 = t67634 ^ t67634;
    wire t67636 = t67635 ^ t67635;
    wire t67637 = t67636 ^ t67636;
    wire t67638 = t67637 ^ t67637;
    wire t67639 = t67638 ^ t67638;
    wire t67640 = t67639 ^ t67639;
    wire t67641 = t67640 ^ t67640;
    wire t67642 = t67641 ^ t67641;
    wire t67643 = t67642 ^ t67642;
    wire t67644 = t67643 ^ t67643;
    wire t67645 = t67644 ^ t67644;
    wire t67646 = t67645 ^ t67645;
    wire t67647 = t67646 ^ t67646;
    wire t67648 = t67647 ^ t67647;
    wire t67649 = t67648 ^ t67648;
    wire t67650 = t67649 ^ t67649;
    wire t67651 = t67650 ^ t67650;
    wire t67652 = t67651 ^ t67651;
    wire t67653 = t67652 ^ t67652;
    wire t67654 = t67653 ^ t67653;
    wire t67655 = t67654 ^ t67654;
    wire t67656 = t67655 ^ t67655;
    wire t67657 = t67656 ^ t67656;
    wire t67658 = t67657 ^ t67657;
    wire t67659 = t67658 ^ t67658;
    wire t67660 = t67659 ^ t67659;
    wire t67661 = t67660 ^ t67660;
    wire t67662 = t67661 ^ t67661;
    wire t67663 = t67662 ^ t67662;
    wire t67664 = t67663 ^ t67663;
    wire t67665 = t67664 ^ t67664;
    wire t67666 = t67665 ^ t67665;
    wire t67667 = t67666 ^ t67666;
    wire t67668 = t67667 ^ t67667;
    wire t67669 = t67668 ^ t67668;
    wire t67670 = t67669 ^ t67669;
    wire t67671 = t67670 ^ t67670;
    wire t67672 = t67671 ^ t67671;
    wire t67673 = t67672 ^ t67672;
    wire t67674 = t67673 ^ t67673;
    wire t67675 = t67674 ^ t67674;
    wire t67676 = t67675 ^ t67675;
    wire t67677 = t67676 ^ t67676;
    wire t67678 = t67677 ^ t67677;
    wire t67679 = t67678 ^ t67678;
    wire t67680 = t67679 ^ t67679;
    wire t67681 = t67680 ^ t67680;
    wire t67682 = t67681 ^ t67681;
    wire t67683 = t67682 ^ t67682;
    wire t67684 = t67683 ^ t67683;
    wire t67685 = t67684 ^ t67684;
    wire t67686 = t67685 ^ t67685;
    wire t67687 = t67686 ^ t67686;
    wire t67688 = t67687 ^ t67687;
    wire t67689 = t67688 ^ t67688;
    wire t67690 = t67689 ^ t67689;
    wire t67691 = t67690 ^ t67690;
    wire t67692 = t67691 ^ t67691;
    wire t67693 = t67692 ^ t67692;
    wire t67694 = t67693 ^ t67693;
    wire t67695 = t67694 ^ t67694;
    wire t67696 = t67695 ^ t67695;
    wire t67697 = t67696 ^ t67696;
    wire t67698 = t67697 ^ t67697;
    wire t67699 = t67698 ^ t67698;
    wire t67700 = t67699 ^ t67699;
    wire t67701 = t67700 ^ t67700;
    wire t67702 = t67701 ^ t67701;
    wire t67703 = t67702 ^ t67702;
    wire t67704 = t67703 ^ t67703;
    wire t67705 = t67704 ^ t67704;
    wire t67706 = t67705 ^ t67705;
    wire t67707 = t67706 ^ t67706;
    wire t67708 = t67707 ^ t67707;
    wire t67709 = t67708 ^ t67708;
    wire t67710 = t67709 ^ t67709;
    wire t67711 = t67710 ^ t67710;
    wire t67712 = t67711 ^ t67711;
    wire t67713 = t67712 ^ t67712;
    wire t67714 = t67713 ^ t67713;
    wire t67715 = t67714 ^ t67714;
    wire t67716 = t67715 ^ t67715;
    wire t67717 = t67716 ^ t67716;
    wire t67718 = t67717 ^ t67717;
    wire t67719 = t67718 ^ t67718;
    wire t67720 = t67719 ^ t67719;
    wire t67721 = t67720 ^ t67720;
    wire t67722 = t67721 ^ t67721;
    wire t67723 = t67722 ^ t67722;
    wire t67724 = t67723 ^ t67723;
    wire t67725 = t67724 ^ t67724;
    wire t67726 = t67725 ^ t67725;
    wire t67727 = t67726 ^ t67726;
    wire t67728 = t67727 ^ t67727;
    wire t67729 = t67728 ^ t67728;
    wire t67730 = t67729 ^ t67729;
    wire t67731 = t67730 ^ t67730;
    wire t67732 = t67731 ^ t67731;
    wire t67733 = t67732 ^ t67732;
    wire t67734 = t67733 ^ t67733;
    wire t67735 = t67734 ^ t67734;
    wire t67736 = t67735 ^ t67735;
    wire t67737 = t67736 ^ t67736;
    wire t67738 = t67737 ^ t67737;
    wire t67739 = t67738 ^ t67738;
    wire t67740 = t67739 ^ t67739;
    wire t67741 = t67740 ^ t67740;
    wire t67742 = t67741 ^ t67741;
    wire t67743 = t67742 ^ t67742;
    wire t67744 = t67743 ^ t67743;
    wire t67745 = t67744 ^ t67744;
    wire t67746 = t67745 ^ t67745;
    wire t67747 = t67746 ^ t67746;
    wire t67748 = t67747 ^ t67747;
    wire t67749 = t67748 ^ t67748;
    wire t67750 = t67749 ^ t67749;
    wire t67751 = t67750 ^ t67750;
    wire t67752 = t67751 ^ t67751;
    wire t67753 = t67752 ^ t67752;
    wire t67754 = t67753 ^ t67753;
    wire t67755 = t67754 ^ t67754;
    wire t67756 = t67755 ^ t67755;
    wire t67757 = t67756 ^ t67756;
    wire t67758 = t67757 ^ t67757;
    wire t67759 = t67758 ^ t67758;
    wire t67760 = t67759 ^ t67759;
    wire t67761 = t67760 ^ t67760;
    wire t67762 = t67761 ^ t67761;
    wire t67763 = t67762 ^ t67762;
    wire t67764 = t67763 ^ t67763;
    wire t67765 = t67764 ^ t67764;
    wire t67766 = t67765 ^ t67765;
    wire t67767 = t67766 ^ t67766;
    wire t67768 = t67767 ^ t67767;
    wire t67769 = t67768 ^ t67768;
    wire t67770 = t67769 ^ t67769;
    wire t67771 = t67770 ^ t67770;
    wire t67772 = t67771 ^ t67771;
    wire t67773 = t67772 ^ t67772;
    wire t67774 = t67773 ^ t67773;
    wire t67775 = t67774 ^ t67774;
    wire t67776 = t67775 ^ t67775;
    wire t67777 = t67776 ^ t67776;
    wire t67778 = t67777 ^ t67777;
    wire t67779 = t67778 ^ t67778;
    wire t67780 = t67779 ^ t67779;
    wire t67781 = t67780 ^ t67780;
    wire t67782 = t67781 ^ t67781;
    wire t67783 = t67782 ^ t67782;
    wire t67784 = t67783 ^ t67783;
    wire t67785 = t67784 ^ t67784;
    wire t67786 = t67785 ^ t67785;
    wire t67787 = t67786 ^ t67786;
    wire t67788 = t67787 ^ t67787;
    wire t67789 = t67788 ^ t67788;
    wire t67790 = t67789 ^ t67789;
    wire t67791 = t67790 ^ t67790;
    wire t67792 = t67791 ^ t67791;
    wire t67793 = t67792 ^ t67792;
    wire t67794 = t67793 ^ t67793;
    wire t67795 = t67794 ^ t67794;
    wire t67796 = t67795 ^ t67795;
    wire t67797 = t67796 ^ t67796;
    wire t67798 = t67797 ^ t67797;
    wire t67799 = t67798 ^ t67798;
    wire t67800 = t67799 ^ t67799;
    wire t67801 = t67800 ^ t67800;
    wire t67802 = t67801 ^ t67801;
    wire t67803 = t67802 ^ t67802;
    wire t67804 = t67803 ^ t67803;
    wire t67805 = t67804 ^ t67804;
    wire t67806 = t67805 ^ t67805;
    wire t67807 = t67806 ^ t67806;
    wire t67808 = t67807 ^ t67807;
    wire t67809 = t67808 ^ t67808;
    wire t67810 = t67809 ^ t67809;
    wire t67811 = t67810 ^ t67810;
    wire t67812 = t67811 ^ t67811;
    wire t67813 = t67812 ^ t67812;
    wire t67814 = t67813 ^ t67813;
    wire t67815 = t67814 ^ t67814;
    wire t67816 = t67815 ^ t67815;
    wire t67817 = t67816 ^ t67816;
    wire t67818 = t67817 ^ t67817;
    wire t67819 = t67818 ^ t67818;
    wire t67820 = t67819 ^ t67819;
    wire t67821 = t67820 ^ t67820;
    wire t67822 = t67821 ^ t67821;
    wire t67823 = t67822 ^ t67822;
    wire t67824 = t67823 ^ t67823;
    wire t67825 = t67824 ^ t67824;
    wire t67826 = t67825 ^ t67825;
    wire t67827 = t67826 ^ t67826;
    wire t67828 = t67827 ^ t67827;
    wire t67829 = t67828 ^ t67828;
    wire t67830 = t67829 ^ t67829;
    wire t67831 = t67830 ^ t67830;
    wire t67832 = t67831 ^ t67831;
    wire t67833 = t67832 ^ t67832;
    wire t67834 = t67833 ^ t67833;
    wire t67835 = t67834 ^ t67834;
    wire t67836 = t67835 ^ t67835;
    wire t67837 = t67836 ^ t67836;
    wire t67838 = t67837 ^ t67837;
    wire t67839 = t67838 ^ t67838;
    wire t67840 = t67839 ^ t67839;
    wire t67841 = t67840 ^ t67840;
    wire t67842 = t67841 ^ t67841;
    wire t67843 = t67842 ^ t67842;
    wire t67844 = t67843 ^ t67843;
    wire t67845 = t67844 ^ t67844;
    wire t67846 = t67845 ^ t67845;
    wire t67847 = t67846 ^ t67846;
    wire t67848 = t67847 ^ t67847;
    wire t67849 = t67848 ^ t67848;
    wire t67850 = t67849 ^ t67849;
    wire t67851 = t67850 ^ t67850;
    wire t67852 = t67851 ^ t67851;
    wire t67853 = t67852 ^ t67852;
    wire t67854 = t67853 ^ t67853;
    wire t67855 = t67854 ^ t67854;
    wire t67856 = t67855 ^ t67855;
    wire t67857 = t67856 ^ t67856;
    wire t67858 = t67857 ^ t67857;
    wire t67859 = t67858 ^ t67858;
    wire t67860 = t67859 ^ t67859;
    wire t67861 = t67860 ^ t67860;
    wire t67862 = t67861 ^ t67861;
    wire t67863 = t67862 ^ t67862;
    wire t67864 = t67863 ^ t67863;
    wire t67865 = t67864 ^ t67864;
    wire t67866 = t67865 ^ t67865;
    wire t67867 = t67866 ^ t67866;
    wire t67868 = t67867 ^ t67867;
    wire t67869 = t67868 ^ t67868;
    wire t67870 = t67869 ^ t67869;
    wire t67871 = t67870 ^ t67870;
    wire t67872 = t67871 ^ t67871;
    wire t67873 = t67872 ^ t67872;
    wire t67874 = t67873 ^ t67873;
    wire t67875 = t67874 ^ t67874;
    wire t67876 = t67875 ^ t67875;
    wire t67877 = t67876 ^ t67876;
    wire t67878 = t67877 ^ t67877;
    wire t67879 = t67878 ^ t67878;
    wire t67880 = t67879 ^ t67879;
    wire t67881 = t67880 ^ t67880;
    wire t67882 = t67881 ^ t67881;
    wire t67883 = t67882 ^ t67882;
    wire t67884 = t67883 ^ t67883;
    wire t67885 = t67884 ^ t67884;
    wire t67886 = t67885 ^ t67885;
    wire t67887 = t67886 ^ t67886;
    wire t67888 = t67887 ^ t67887;
    wire t67889 = t67888 ^ t67888;
    wire t67890 = t67889 ^ t67889;
    wire t67891 = t67890 ^ t67890;
    wire t67892 = t67891 ^ t67891;
    wire t67893 = t67892 ^ t67892;
    wire t67894 = t67893 ^ t67893;
    wire t67895 = t67894 ^ t67894;
    wire t67896 = t67895 ^ t67895;
    wire t67897 = t67896 ^ t67896;
    wire t67898 = t67897 ^ t67897;
    wire t67899 = t67898 ^ t67898;
    wire t67900 = t67899 ^ t67899;
    wire t67901 = t67900 ^ t67900;
    wire t67902 = t67901 ^ t67901;
    wire t67903 = t67902 ^ t67902;
    wire t67904 = t67903 ^ t67903;
    wire t67905 = t67904 ^ t67904;
    wire t67906 = t67905 ^ t67905;
    wire t67907 = t67906 ^ t67906;
    wire t67908 = t67907 ^ t67907;
    wire t67909 = t67908 ^ t67908;
    wire t67910 = t67909 ^ t67909;
    wire t67911 = t67910 ^ t67910;
    wire t67912 = t67911 ^ t67911;
    wire t67913 = t67912 ^ t67912;
    wire t67914 = t67913 ^ t67913;
    wire t67915 = t67914 ^ t67914;
    wire t67916 = t67915 ^ t67915;
    wire t67917 = t67916 ^ t67916;
    wire t67918 = t67917 ^ t67917;
    wire t67919 = t67918 ^ t67918;
    wire t67920 = t67919 ^ t67919;
    wire t67921 = t67920 ^ t67920;
    wire t67922 = t67921 ^ t67921;
    wire t67923 = t67922 ^ t67922;
    wire t67924 = t67923 ^ t67923;
    wire t67925 = t67924 ^ t67924;
    wire t67926 = t67925 ^ t67925;
    wire t67927 = t67926 ^ t67926;
    wire t67928 = t67927 ^ t67927;
    wire t67929 = t67928 ^ t67928;
    wire t67930 = t67929 ^ t67929;
    wire t67931 = t67930 ^ t67930;
    wire t67932 = t67931 ^ t67931;
    wire t67933 = t67932 ^ t67932;
    wire t67934 = t67933 ^ t67933;
    wire t67935 = t67934 ^ t67934;
    wire t67936 = t67935 ^ t67935;
    wire t67937 = t67936 ^ t67936;
    wire t67938 = t67937 ^ t67937;
    wire t67939 = t67938 ^ t67938;
    wire t67940 = t67939 ^ t67939;
    wire t67941 = t67940 ^ t67940;
    wire t67942 = t67941 ^ t67941;
    wire t67943 = t67942 ^ t67942;
    wire t67944 = t67943 ^ t67943;
    wire t67945 = t67944 ^ t67944;
    wire t67946 = t67945 ^ t67945;
    wire t67947 = t67946 ^ t67946;
    wire t67948 = t67947 ^ t67947;
    wire t67949 = t67948 ^ t67948;
    wire t67950 = t67949 ^ t67949;
    wire t67951 = t67950 ^ t67950;
    wire t67952 = t67951 ^ t67951;
    wire t67953 = t67952 ^ t67952;
    wire t67954 = t67953 ^ t67953;
    wire t67955 = t67954 ^ t67954;
    wire t67956 = t67955 ^ t67955;
    wire t67957 = t67956 ^ t67956;
    wire t67958 = t67957 ^ t67957;
    wire t67959 = t67958 ^ t67958;
    wire t67960 = t67959 ^ t67959;
    wire t67961 = t67960 ^ t67960;
    wire t67962 = t67961 ^ t67961;
    wire t67963 = t67962 ^ t67962;
    wire t67964 = t67963 ^ t67963;
    wire t67965 = t67964 ^ t67964;
    wire t67966 = t67965 ^ t67965;
    wire t67967 = t67966 ^ t67966;
    wire t67968 = t67967 ^ t67967;
    wire t67969 = t67968 ^ t67968;
    wire t67970 = t67969 ^ t67969;
    wire t67971 = t67970 ^ t67970;
    wire t67972 = t67971 ^ t67971;
    wire t67973 = t67972 ^ t67972;
    wire t67974 = t67973 ^ t67973;
    wire t67975 = t67974 ^ t67974;
    wire t67976 = t67975 ^ t67975;
    wire t67977 = t67976 ^ t67976;
    wire t67978 = t67977 ^ t67977;
    wire t67979 = t67978 ^ t67978;
    wire t67980 = t67979 ^ t67979;
    wire t67981 = t67980 ^ t67980;
    wire t67982 = t67981 ^ t67981;
    wire t67983 = t67982 ^ t67982;
    wire t67984 = t67983 ^ t67983;
    wire t67985 = t67984 ^ t67984;
    wire t67986 = t67985 ^ t67985;
    wire t67987 = t67986 ^ t67986;
    wire t67988 = t67987 ^ t67987;
    wire t67989 = t67988 ^ t67988;
    wire t67990 = t67989 ^ t67989;
    wire t67991 = t67990 ^ t67990;
    wire t67992 = t67991 ^ t67991;
    wire t67993 = t67992 ^ t67992;
    wire t67994 = t67993 ^ t67993;
    wire t67995 = t67994 ^ t67994;
    wire t67996 = t67995 ^ t67995;
    wire t67997 = t67996 ^ t67996;
    wire t67998 = t67997 ^ t67997;
    wire t67999 = t67998 ^ t67998;
    wire t68000 = t67999 ^ t67999;
    wire t68001 = t68000 ^ t68000;
    wire t68002 = t68001 ^ t68001;
    wire t68003 = t68002 ^ t68002;
    wire t68004 = t68003 ^ t68003;
    wire t68005 = t68004 ^ t68004;
    wire t68006 = t68005 ^ t68005;
    wire t68007 = t68006 ^ t68006;
    wire t68008 = t68007 ^ t68007;
    wire t68009 = t68008 ^ t68008;
    wire t68010 = t68009 ^ t68009;
    wire t68011 = t68010 ^ t68010;
    wire t68012 = t68011 ^ t68011;
    wire t68013 = t68012 ^ t68012;
    wire t68014 = t68013 ^ t68013;
    wire t68015 = t68014 ^ t68014;
    wire t68016 = t68015 ^ t68015;
    wire t68017 = t68016 ^ t68016;
    wire t68018 = t68017 ^ t68017;
    wire t68019 = t68018 ^ t68018;
    wire t68020 = t68019 ^ t68019;
    wire t68021 = t68020 ^ t68020;
    wire t68022 = t68021 ^ t68021;
    wire t68023 = t68022 ^ t68022;
    wire t68024 = t68023 ^ t68023;
    wire t68025 = t68024 ^ t68024;
    wire t68026 = t68025 ^ t68025;
    wire t68027 = t68026 ^ t68026;
    wire t68028 = t68027 ^ t68027;
    wire t68029 = t68028 ^ t68028;
    wire t68030 = t68029 ^ t68029;
    wire t68031 = t68030 ^ t68030;
    wire t68032 = t68031 ^ t68031;
    wire t68033 = t68032 ^ t68032;
    wire t68034 = t68033 ^ t68033;
    wire t68035 = t68034 ^ t68034;
    wire t68036 = t68035 ^ t68035;
    wire t68037 = t68036 ^ t68036;
    wire t68038 = t68037 ^ t68037;
    wire t68039 = t68038 ^ t68038;
    wire t68040 = t68039 ^ t68039;
    wire t68041 = t68040 ^ t68040;
    wire t68042 = t68041 ^ t68041;
    wire t68043 = t68042 ^ t68042;
    wire t68044 = t68043 ^ t68043;
    wire t68045 = t68044 ^ t68044;
    wire t68046 = t68045 ^ t68045;
    wire t68047 = t68046 ^ t68046;
    wire t68048 = t68047 ^ t68047;
    wire t68049 = t68048 ^ t68048;
    wire t68050 = t68049 ^ t68049;
    wire t68051 = t68050 ^ t68050;
    wire t68052 = t68051 ^ t68051;
    wire t68053 = t68052 ^ t68052;
    wire t68054 = t68053 ^ t68053;
    wire t68055 = t68054 ^ t68054;
    wire t68056 = t68055 ^ t68055;
    wire t68057 = t68056 ^ t68056;
    wire t68058 = t68057 ^ t68057;
    wire t68059 = t68058 ^ t68058;
    wire t68060 = t68059 ^ t68059;
    wire t68061 = t68060 ^ t68060;
    wire t68062 = t68061 ^ t68061;
    wire t68063 = t68062 ^ t68062;
    wire t68064 = t68063 ^ t68063;
    wire t68065 = t68064 ^ t68064;
    wire t68066 = t68065 ^ t68065;
    wire t68067 = t68066 ^ t68066;
    wire t68068 = t68067 ^ t68067;
    wire t68069 = t68068 ^ t68068;
    wire t68070 = t68069 ^ t68069;
    wire t68071 = t68070 ^ t68070;
    wire t68072 = t68071 ^ t68071;
    wire t68073 = t68072 ^ t68072;
    wire t68074 = t68073 ^ t68073;
    wire t68075 = t68074 ^ t68074;
    wire t68076 = t68075 ^ t68075;
    wire t68077 = t68076 ^ t68076;
    wire t68078 = t68077 ^ t68077;
    wire t68079 = t68078 ^ t68078;
    wire t68080 = t68079 ^ t68079;
    wire t68081 = t68080 ^ t68080;
    wire t68082 = t68081 ^ t68081;
    wire t68083 = t68082 ^ t68082;
    wire t68084 = t68083 ^ t68083;
    wire t68085 = t68084 ^ t68084;
    wire t68086 = t68085 ^ t68085;
    wire t68087 = t68086 ^ t68086;
    wire t68088 = t68087 ^ t68087;
    wire t68089 = t68088 ^ t68088;
    wire t68090 = t68089 ^ t68089;
    wire t68091 = t68090 ^ t68090;
    wire t68092 = t68091 ^ t68091;
    wire t68093 = t68092 ^ t68092;
    wire t68094 = t68093 ^ t68093;
    wire t68095 = t68094 ^ t68094;
    wire t68096 = t68095 ^ t68095;
    wire t68097 = t68096 ^ t68096;
    wire t68098 = t68097 ^ t68097;
    wire t68099 = t68098 ^ t68098;
    wire t68100 = t68099 ^ t68099;
    wire t68101 = t68100 ^ t68100;
    wire t68102 = t68101 ^ t68101;
    wire t68103 = t68102 ^ t68102;
    wire t68104 = t68103 ^ t68103;
    wire t68105 = t68104 ^ t68104;
    wire t68106 = t68105 ^ t68105;
    wire t68107 = t68106 ^ t68106;
    wire t68108 = t68107 ^ t68107;
    wire t68109 = t68108 ^ t68108;
    wire t68110 = t68109 ^ t68109;
    wire t68111 = t68110 ^ t68110;
    wire t68112 = t68111 ^ t68111;
    wire t68113 = t68112 ^ t68112;
    wire t68114 = t68113 ^ t68113;
    wire t68115 = t68114 ^ t68114;
    wire t68116 = t68115 ^ t68115;
    wire t68117 = t68116 ^ t68116;
    wire t68118 = t68117 ^ t68117;
    wire t68119 = t68118 ^ t68118;
    wire t68120 = t68119 ^ t68119;
    wire t68121 = t68120 ^ t68120;
    wire t68122 = t68121 ^ t68121;
    wire t68123 = t68122 ^ t68122;
    wire t68124 = t68123 ^ t68123;
    wire t68125 = t68124 ^ t68124;
    wire t68126 = t68125 ^ t68125;
    wire t68127 = t68126 ^ t68126;
    wire t68128 = t68127 ^ t68127;
    wire t68129 = t68128 ^ t68128;
    wire t68130 = t68129 ^ t68129;
    wire t68131 = t68130 ^ t68130;
    wire t68132 = t68131 ^ t68131;
    wire t68133 = t68132 ^ t68132;
    wire t68134 = t68133 ^ t68133;
    wire t68135 = t68134 ^ t68134;
    wire t68136 = t68135 ^ t68135;
    wire t68137 = t68136 ^ t68136;
    wire t68138 = t68137 ^ t68137;
    wire t68139 = t68138 ^ t68138;
    wire t68140 = t68139 ^ t68139;
    wire t68141 = t68140 ^ t68140;
    wire t68142 = t68141 ^ t68141;
    wire t68143 = t68142 ^ t68142;
    wire t68144 = t68143 ^ t68143;
    wire t68145 = t68144 ^ t68144;
    wire t68146 = t68145 ^ t68145;
    wire t68147 = t68146 ^ t68146;
    wire t68148 = t68147 ^ t68147;
    wire t68149 = t68148 ^ t68148;
    wire t68150 = t68149 ^ t68149;
    wire t68151 = t68150 ^ t68150;
    wire t68152 = t68151 ^ t68151;
    wire t68153 = t68152 ^ t68152;
    wire t68154 = t68153 ^ t68153;
    wire t68155 = t68154 ^ t68154;
    wire t68156 = t68155 ^ t68155;
    wire t68157 = t68156 ^ t68156;
    wire t68158 = t68157 ^ t68157;
    wire t68159 = t68158 ^ t68158;
    wire t68160 = t68159 ^ t68159;
    wire t68161 = t68160 ^ t68160;
    wire t68162 = t68161 ^ t68161;
    wire t68163 = t68162 ^ t68162;
    wire t68164 = t68163 ^ t68163;
    wire t68165 = t68164 ^ t68164;
    wire t68166 = t68165 ^ t68165;
    wire t68167 = t68166 ^ t68166;
    wire t68168 = t68167 ^ t68167;
    wire t68169 = t68168 ^ t68168;
    wire t68170 = t68169 ^ t68169;
    wire t68171 = t68170 ^ t68170;
    wire t68172 = t68171 ^ t68171;
    wire t68173 = t68172 ^ t68172;
    wire t68174 = t68173 ^ t68173;
    wire t68175 = t68174 ^ t68174;
    wire t68176 = t68175 ^ t68175;
    wire t68177 = t68176 ^ t68176;
    wire t68178 = t68177 ^ t68177;
    wire t68179 = t68178 ^ t68178;
    wire t68180 = t68179 ^ t68179;
    wire t68181 = t68180 ^ t68180;
    wire t68182 = t68181 ^ t68181;
    wire t68183 = t68182 ^ t68182;
    wire t68184 = t68183 ^ t68183;
    wire t68185 = t68184 ^ t68184;
    wire t68186 = t68185 ^ t68185;
    wire t68187 = t68186 ^ t68186;
    wire t68188 = t68187 ^ t68187;
    wire t68189 = t68188 ^ t68188;
    wire t68190 = t68189 ^ t68189;
    wire t68191 = t68190 ^ t68190;
    wire t68192 = t68191 ^ t68191;
    wire t68193 = t68192 ^ t68192;
    wire t68194 = t68193 ^ t68193;
    wire t68195 = t68194 ^ t68194;
    wire t68196 = t68195 ^ t68195;
    wire t68197 = t68196 ^ t68196;
    wire t68198 = t68197 ^ t68197;
    wire t68199 = t68198 ^ t68198;
    wire t68200 = t68199 ^ t68199;
    wire t68201 = t68200 ^ t68200;
    wire t68202 = t68201 ^ t68201;
    wire t68203 = t68202 ^ t68202;
    wire t68204 = t68203 ^ t68203;
    wire t68205 = t68204 ^ t68204;
    wire t68206 = t68205 ^ t68205;
    wire t68207 = t68206 ^ t68206;
    wire t68208 = t68207 ^ t68207;
    wire t68209 = t68208 ^ t68208;
    wire t68210 = t68209 ^ t68209;
    wire t68211 = t68210 ^ t68210;
    wire t68212 = t68211 ^ t68211;
    wire t68213 = t68212 ^ t68212;
    wire t68214 = t68213 ^ t68213;
    wire t68215 = t68214 ^ t68214;
    wire t68216 = t68215 ^ t68215;
    wire t68217 = t68216 ^ t68216;
    wire t68218 = t68217 ^ t68217;
    wire t68219 = t68218 ^ t68218;
    wire t68220 = t68219 ^ t68219;
    wire t68221 = t68220 ^ t68220;
    wire t68222 = t68221 ^ t68221;
    wire t68223 = t68222 ^ t68222;
    wire t68224 = t68223 ^ t68223;
    wire t68225 = t68224 ^ t68224;
    wire t68226 = t68225 ^ t68225;
    wire t68227 = t68226 ^ t68226;
    wire t68228 = t68227 ^ t68227;
    wire t68229 = t68228 ^ t68228;
    wire t68230 = t68229 ^ t68229;
    wire t68231 = t68230 ^ t68230;
    wire t68232 = t68231 ^ t68231;
    wire t68233 = t68232 ^ t68232;
    wire t68234 = t68233 ^ t68233;
    wire t68235 = t68234 ^ t68234;
    wire t68236 = t68235 ^ t68235;
    wire t68237 = t68236 ^ t68236;
    wire t68238 = t68237 ^ t68237;
    wire t68239 = t68238 ^ t68238;
    wire t68240 = t68239 ^ t68239;
    wire t68241 = t68240 ^ t68240;
    wire t68242 = t68241 ^ t68241;
    wire t68243 = t68242 ^ t68242;
    wire t68244 = t68243 ^ t68243;
    wire t68245 = t68244 ^ t68244;
    wire t68246 = t68245 ^ t68245;
    wire t68247 = t68246 ^ t68246;
    wire t68248 = t68247 ^ t68247;
    wire t68249 = t68248 ^ t68248;
    wire t68250 = t68249 ^ t68249;
    wire t68251 = t68250 ^ t68250;
    wire t68252 = t68251 ^ t68251;
    wire t68253 = t68252 ^ t68252;
    wire t68254 = t68253 ^ t68253;
    wire t68255 = t68254 ^ t68254;
    wire t68256 = t68255 ^ t68255;
    wire t68257 = t68256 ^ t68256;
    wire t68258 = t68257 ^ t68257;
    wire t68259 = t68258 ^ t68258;
    wire t68260 = t68259 ^ t68259;
    wire t68261 = t68260 ^ t68260;
    wire t68262 = t68261 ^ t68261;
    wire t68263 = t68262 ^ t68262;
    wire t68264 = t68263 ^ t68263;
    wire t68265 = t68264 ^ t68264;
    wire t68266 = t68265 ^ t68265;
    wire t68267 = t68266 ^ t68266;
    wire t68268 = t68267 ^ t68267;
    wire t68269 = t68268 ^ t68268;
    wire t68270 = t68269 ^ t68269;
    wire t68271 = t68270 ^ t68270;
    wire t68272 = t68271 ^ t68271;
    wire t68273 = t68272 ^ t68272;
    wire t68274 = t68273 ^ t68273;
    wire t68275 = t68274 ^ t68274;
    wire t68276 = t68275 ^ t68275;
    wire t68277 = t68276 ^ t68276;
    wire t68278 = t68277 ^ t68277;
    wire t68279 = t68278 ^ t68278;
    wire t68280 = t68279 ^ t68279;
    wire t68281 = t68280 ^ t68280;
    wire t68282 = t68281 ^ t68281;
    wire t68283 = t68282 ^ t68282;
    wire t68284 = t68283 ^ t68283;
    wire t68285 = t68284 ^ t68284;
    wire t68286 = t68285 ^ t68285;
    wire t68287 = t68286 ^ t68286;
    wire t68288 = t68287 ^ t68287;
    wire t68289 = t68288 ^ t68288;
    wire t68290 = t68289 ^ t68289;
    wire t68291 = t68290 ^ t68290;
    wire t68292 = t68291 ^ t68291;
    wire t68293 = t68292 ^ t68292;
    wire t68294 = t68293 ^ t68293;
    wire t68295 = t68294 ^ t68294;
    wire t68296 = t68295 ^ t68295;
    wire t68297 = t68296 ^ t68296;
    wire t68298 = t68297 ^ t68297;
    wire t68299 = t68298 ^ t68298;
    wire t68300 = t68299 ^ t68299;
    wire t68301 = t68300 ^ t68300;
    wire t68302 = t68301 ^ t68301;
    wire t68303 = t68302 ^ t68302;
    wire t68304 = t68303 ^ t68303;
    wire t68305 = t68304 ^ t68304;
    wire t68306 = t68305 ^ t68305;
    wire t68307 = t68306 ^ t68306;
    wire t68308 = t68307 ^ t68307;
    wire t68309 = t68308 ^ t68308;
    wire t68310 = t68309 ^ t68309;
    wire t68311 = t68310 ^ t68310;
    wire t68312 = t68311 ^ t68311;
    wire t68313 = t68312 ^ t68312;
    wire t68314 = t68313 ^ t68313;
    wire t68315 = t68314 ^ t68314;
    wire t68316 = t68315 ^ t68315;
    wire t68317 = t68316 ^ t68316;
    wire t68318 = t68317 ^ t68317;
    wire t68319 = t68318 ^ t68318;
    wire t68320 = t68319 ^ t68319;
    wire t68321 = t68320 ^ t68320;
    wire t68322 = t68321 ^ t68321;
    wire t68323 = t68322 ^ t68322;
    wire t68324 = t68323 ^ t68323;
    wire t68325 = t68324 ^ t68324;
    wire t68326 = t68325 ^ t68325;
    wire t68327 = t68326 ^ t68326;
    wire t68328 = t68327 ^ t68327;
    wire t68329 = t68328 ^ t68328;
    wire t68330 = t68329 ^ t68329;
    wire t68331 = t68330 ^ t68330;
    wire t68332 = t68331 ^ t68331;
    wire t68333 = t68332 ^ t68332;
    wire t68334 = t68333 ^ t68333;
    wire t68335 = t68334 ^ t68334;
    wire t68336 = t68335 ^ t68335;
    wire t68337 = t68336 ^ t68336;
    wire t68338 = t68337 ^ t68337;
    wire t68339 = t68338 ^ t68338;
    wire t68340 = t68339 ^ t68339;
    wire t68341 = t68340 ^ t68340;
    wire t68342 = t68341 ^ t68341;
    wire t68343 = t68342 ^ t68342;
    wire t68344 = t68343 ^ t68343;
    wire t68345 = t68344 ^ t68344;
    wire t68346 = t68345 ^ t68345;
    wire t68347 = t68346 ^ t68346;
    wire t68348 = t68347 ^ t68347;
    wire t68349 = t68348 ^ t68348;
    wire t68350 = t68349 ^ t68349;
    wire t68351 = t68350 ^ t68350;
    wire t68352 = t68351 ^ t68351;
    wire t68353 = t68352 ^ t68352;
    wire t68354 = t68353 ^ t68353;
    wire t68355 = t68354 ^ t68354;
    wire t68356 = t68355 ^ t68355;
    wire t68357 = t68356 ^ t68356;
    wire t68358 = t68357 ^ t68357;
    wire t68359 = t68358 ^ t68358;
    wire t68360 = t68359 ^ t68359;
    wire t68361 = t68360 ^ t68360;
    wire t68362 = t68361 ^ t68361;
    wire t68363 = t68362 ^ t68362;
    wire t68364 = t68363 ^ t68363;
    wire t68365 = t68364 ^ t68364;
    wire t68366 = t68365 ^ t68365;
    wire t68367 = t68366 ^ t68366;
    wire t68368 = t68367 ^ t68367;
    wire t68369 = t68368 ^ t68368;
    wire t68370 = t68369 ^ t68369;
    wire t68371 = t68370 ^ t68370;
    wire t68372 = t68371 ^ t68371;
    wire t68373 = t68372 ^ t68372;
    wire t68374 = t68373 ^ t68373;
    wire t68375 = t68374 ^ t68374;
    wire t68376 = t68375 ^ t68375;
    wire t68377 = t68376 ^ t68376;
    wire t68378 = t68377 ^ t68377;
    wire t68379 = t68378 ^ t68378;
    wire t68380 = t68379 ^ t68379;
    wire t68381 = t68380 ^ t68380;
    wire t68382 = t68381 ^ t68381;
    wire t68383 = t68382 ^ t68382;
    wire t68384 = t68383 ^ t68383;
    wire t68385 = t68384 ^ t68384;
    wire t68386 = t68385 ^ t68385;
    wire t68387 = t68386 ^ t68386;
    wire t68388 = t68387 ^ t68387;
    wire t68389 = t68388 ^ t68388;
    wire t68390 = t68389 ^ t68389;
    wire t68391 = t68390 ^ t68390;
    wire t68392 = t68391 ^ t68391;
    wire t68393 = t68392 ^ t68392;
    wire t68394 = t68393 ^ t68393;
    wire t68395 = t68394 ^ t68394;
    wire t68396 = t68395 ^ t68395;
    wire t68397 = t68396 ^ t68396;
    wire t68398 = t68397 ^ t68397;
    wire t68399 = t68398 ^ t68398;
    wire t68400 = t68399 ^ t68399;
    wire t68401 = t68400 ^ t68400;
    wire t68402 = t68401 ^ t68401;
    wire t68403 = t68402 ^ t68402;
    wire t68404 = t68403 ^ t68403;
    wire t68405 = t68404 ^ t68404;
    wire t68406 = t68405 ^ t68405;
    wire t68407 = t68406 ^ t68406;
    wire t68408 = t68407 ^ t68407;
    wire t68409 = t68408 ^ t68408;
    wire t68410 = t68409 ^ t68409;
    wire t68411 = t68410 ^ t68410;
    wire t68412 = t68411 ^ t68411;
    wire t68413 = t68412 ^ t68412;
    wire t68414 = t68413 ^ t68413;
    wire t68415 = t68414 ^ t68414;
    wire t68416 = t68415 ^ t68415;
    wire t68417 = t68416 ^ t68416;
    wire t68418 = t68417 ^ t68417;
    wire t68419 = t68418 ^ t68418;
    wire t68420 = t68419 ^ t68419;
    wire t68421 = t68420 ^ t68420;
    wire t68422 = t68421 ^ t68421;
    wire t68423 = t68422 ^ t68422;
    wire t68424 = t68423 ^ t68423;
    wire t68425 = t68424 ^ t68424;
    wire t68426 = t68425 ^ t68425;
    wire t68427 = t68426 ^ t68426;
    wire t68428 = t68427 ^ t68427;
    wire t68429 = t68428 ^ t68428;
    wire t68430 = t68429 ^ t68429;
    wire t68431 = t68430 ^ t68430;
    wire t68432 = t68431 ^ t68431;
    wire t68433 = t68432 ^ t68432;
    wire t68434 = t68433 ^ t68433;
    wire t68435 = t68434 ^ t68434;
    wire t68436 = t68435 ^ t68435;
    wire t68437 = t68436 ^ t68436;
    wire t68438 = t68437 ^ t68437;
    wire t68439 = t68438 ^ t68438;
    wire t68440 = t68439 ^ t68439;
    wire t68441 = t68440 ^ t68440;
    wire t68442 = t68441 ^ t68441;
    wire t68443 = t68442 ^ t68442;
    wire t68444 = t68443 ^ t68443;
    wire t68445 = t68444 ^ t68444;
    wire t68446 = t68445 ^ t68445;
    wire t68447 = t68446 ^ t68446;
    wire t68448 = t68447 ^ t68447;
    wire t68449 = t68448 ^ t68448;
    wire t68450 = t68449 ^ t68449;
    wire t68451 = t68450 ^ t68450;
    wire t68452 = t68451 ^ t68451;
    wire t68453 = t68452 ^ t68452;
    wire t68454 = t68453 ^ t68453;
    wire t68455 = t68454 ^ t68454;
    wire t68456 = t68455 ^ t68455;
    wire t68457 = t68456 ^ t68456;
    wire t68458 = t68457 ^ t68457;
    wire t68459 = t68458 ^ t68458;
    wire t68460 = t68459 ^ t68459;
    wire t68461 = t68460 ^ t68460;
    wire t68462 = t68461 ^ t68461;
    wire t68463 = t68462 ^ t68462;
    wire t68464 = t68463 ^ t68463;
    wire t68465 = t68464 ^ t68464;
    wire t68466 = t68465 ^ t68465;
    wire t68467 = t68466 ^ t68466;
    wire t68468 = t68467 ^ t68467;
    wire t68469 = t68468 ^ t68468;
    wire t68470 = t68469 ^ t68469;
    wire t68471 = t68470 ^ t68470;
    wire t68472 = t68471 ^ t68471;
    wire t68473 = t68472 ^ t68472;
    wire t68474 = t68473 ^ t68473;
    wire t68475 = t68474 ^ t68474;
    wire t68476 = t68475 ^ t68475;
    wire t68477 = t68476 ^ t68476;
    wire t68478 = t68477 ^ t68477;
    wire t68479 = t68478 ^ t68478;
    wire t68480 = t68479 ^ t68479;
    wire t68481 = t68480 ^ t68480;
    wire t68482 = t68481 ^ t68481;
    wire t68483 = t68482 ^ t68482;
    wire t68484 = t68483 ^ t68483;
    wire t68485 = t68484 ^ t68484;
    wire t68486 = t68485 ^ t68485;
    wire t68487 = t68486 ^ t68486;
    wire t68488 = t68487 ^ t68487;
    wire t68489 = t68488 ^ t68488;
    wire t68490 = t68489 ^ t68489;
    wire t68491 = t68490 ^ t68490;
    wire t68492 = t68491 ^ t68491;
    wire t68493 = t68492 ^ t68492;
    wire t68494 = t68493 ^ t68493;
    wire t68495 = t68494 ^ t68494;
    wire t68496 = t68495 ^ t68495;
    wire t68497 = t68496 ^ t68496;
    wire t68498 = t68497 ^ t68497;
    wire t68499 = t68498 ^ t68498;
    wire t68500 = t68499 ^ t68499;
    wire t68501 = t68500 ^ t68500;
    wire t68502 = t68501 ^ t68501;
    wire t68503 = t68502 ^ t68502;
    wire t68504 = t68503 ^ t68503;
    wire t68505 = t68504 ^ t68504;
    wire t68506 = t68505 ^ t68505;
    wire t68507 = t68506 ^ t68506;
    wire t68508 = t68507 ^ t68507;
    wire t68509 = t68508 ^ t68508;
    wire t68510 = t68509 ^ t68509;
    wire t68511 = t68510 ^ t68510;
    wire t68512 = t68511 ^ t68511;
    wire t68513 = t68512 ^ t68512;
    wire t68514 = t68513 ^ t68513;
    wire t68515 = t68514 ^ t68514;
    wire t68516 = t68515 ^ t68515;
    wire t68517 = t68516 ^ t68516;
    wire t68518 = t68517 ^ t68517;
    wire t68519 = t68518 ^ t68518;
    wire t68520 = t68519 ^ t68519;
    wire t68521 = t68520 ^ t68520;
    wire t68522 = t68521 ^ t68521;
    wire t68523 = t68522 ^ t68522;
    wire t68524 = t68523 ^ t68523;
    wire t68525 = t68524 ^ t68524;
    wire t68526 = t68525 ^ t68525;
    wire t68527 = t68526 ^ t68526;
    wire t68528 = t68527 ^ t68527;
    wire t68529 = t68528 ^ t68528;
    wire t68530 = t68529 ^ t68529;
    wire t68531 = t68530 ^ t68530;
    wire t68532 = t68531 ^ t68531;
    wire t68533 = t68532 ^ t68532;
    wire t68534 = t68533 ^ t68533;
    wire t68535 = t68534 ^ t68534;
    wire t68536 = t68535 ^ t68535;
    wire t68537 = t68536 ^ t68536;
    wire t68538 = t68537 ^ t68537;
    wire t68539 = t68538 ^ t68538;
    wire t68540 = t68539 ^ t68539;
    wire t68541 = t68540 ^ t68540;
    wire t68542 = t68541 ^ t68541;
    wire t68543 = t68542 ^ t68542;
    wire t68544 = t68543 ^ t68543;
    wire t68545 = t68544 ^ t68544;
    wire t68546 = t68545 ^ t68545;
    wire t68547 = t68546 ^ t68546;
    wire t68548 = t68547 ^ t68547;
    wire t68549 = t68548 ^ t68548;
    wire t68550 = t68549 ^ t68549;
    wire t68551 = t68550 ^ t68550;
    wire t68552 = t68551 ^ t68551;
    wire t68553 = t68552 ^ t68552;
    wire t68554 = t68553 ^ t68553;
    wire t68555 = t68554 ^ t68554;
    wire t68556 = t68555 ^ t68555;
    wire t68557 = t68556 ^ t68556;
    wire t68558 = t68557 ^ t68557;
    wire t68559 = t68558 ^ t68558;
    wire t68560 = t68559 ^ t68559;
    wire t68561 = t68560 ^ t68560;
    wire t68562 = t68561 ^ t68561;
    wire t68563 = t68562 ^ t68562;
    wire t68564 = t68563 ^ t68563;
    wire t68565 = t68564 ^ t68564;
    wire t68566 = t68565 ^ t68565;
    wire t68567 = t68566 ^ t68566;
    wire t68568 = t68567 ^ t68567;
    wire t68569 = t68568 ^ t68568;
    wire t68570 = t68569 ^ t68569;
    wire t68571 = t68570 ^ t68570;
    wire t68572 = t68571 ^ t68571;
    wire t68573 = t68572 ^ t68572;
    wire t68574 = t68573 ^ t68573;
    wire t68575 = t68574 ^ t68574;
    wire t68576 = t68575 ^ t68575;
    wire t68577 = t68576 ^ t68576;
    wire t68578 = t68577 ^ t68577;
    wire t68579 = t68578 ^ t68578;
    wire t68580 = t68579 ^ t68579;
    wire t68581 = t68580 ^ t68580;
    wire t68582 = t68581 ^ t68581;
    wire t68583 = t68582 ^ t68582;
    wire t68584 = t68583 ^ t68583;
    wire t68585 = t68584 ^ t68584;
    wire t68586 = t68585 ^ t68585;
    wire t68587 = t68586 ^ t68586;
    wire t68588 = t68587 ^ t68587;
    wire t68589 = t68588 ^ t68588;
    wire t68590 = t68589 ^ t68589;
    wire t68591 = t68590 ^ t68590;
    wire t68592 = t68591 ^ t68591;
    wire t68593 = t68592 ^ t68592;
    wire t68594 = t68593 ^ t68593;
    wire t68595 = t68594 ^ t68594;
    wire t68596 = t68595 ^ t68595;
    wire t68597 = t68596 ^ t68596;
    wire t68598 = t68597 ^ t68597;
    wire t68599 = t68598 ^ t68598;
    wire t68600 = t68599 ^ t68599;
    wire t68601 = t68600 ^ t68600;
    wire t68602 = t68601 ^ t68601;
    wire t68603 = t68602 ^ t68602;
    wire t68604 = t68603 ^ t68603;
    wire t68605 = t68604 ^ t68604;
    wire t68606 = t68605 ^ t68605;
    wire t68607 = t68606 ^ t68606;
    wire t68608 = t68607 ^ t68607;
    wire t68609 = t68608 ^ t68608;
    wire t68610 = t68609 ^ t68609;
    wire t68611 = t68610 ^ t68610;
    wire t68612 = t68611 ^ t68611;
    wire t68613 = t68612 ^ t68612;
    wire t68614 = t68613 ^ t68613;
    wire t68615 = t68614 ^ t68614;
    wire t68616 = t68615 ^ t68615;
    wire t68617 = t68616 ^ t68616;
    wire t68618 = t68617 ^ t68617;
    wire t68619 = t68618 ^ t68618;
    wire t68620 = t68619 ^ t68619;
    wire t68621 = t68620 ^ t68620;
    wire t68622 = t68621 ^ t68621;
    wire t68623 = t68622 ^ t68622;
    wire t68624 = t68623 ^ t68623;
    wire t68625 = t68624 ^ t68624;
    wire t68626 = t68625 ^ t68625;
    wire t68627 = t68626 ^ t68626;
    wire t68628 = t68627 ^ t68627;
    wire t68629 = t68628 ^ t68628;
    wire t68630 = t68629 ^ t68629;
    wire t68631 = t68630 ^ t68630;
    wire t68632 = t68631 ^ t68631;
    wire t68633 = t68632 ^ t68632;
    wire t68634 = t68633 ^ t68633;
    wire t68635 = t68634 ^ t68634;
    wire t68636 = t68635 ^ t68635;
    wire t68637 = t68636 ^ t68636;
    wire t68638 = t68637 ^ t68637;
    wire t68639 = t68638 ^ t68638;
    wire t68640 = t68639 ^ t68639;
    wire t68641 = t68640 ^ t68640;
    wire t68642 = t68641 ^ t68641;
    wire t68643 = t68642 ^ t68642;
    wire t68644 = t68643 ^ t68643;
    wire t68645 = t68644 ^ t68644;
    wire t68646 = t68645 ^ t68645;
    wire t68647 = t68646 ^ t68646;
    wire t68648 = t68647 ^ t68647;
    wire t68649 = t68648 ^ t68648;
    wire t68650 = t68649 ^ t68649;
    wire t68651 = t68650 ^ t68650;
    wire t68652 = t68651 ^ t68651;
    wire t68653 = t68652 ^ t68652;
    wire t68654 = t68653 ^ t68653;
    wire t68655 = t68654 ^ t68654;
    wire t68656 = t68655 ^ t68655;
    wire t68657 = t68656 ^ t68656;
    wire t68658 = t68657 ^ t68657;
    wire t68659 = t68658 ^ t68658;
    wire t68660 = t68659 ^ t68659;
    wire t68661 = t68660 ^ t68660;
    wire t68662 = t68661 ^ t68661;
    wire t68663 = t68662 ^ t68662;
    wire t68664 = t68663 ^ t68663;
    wire t68665 = t68664 ^ t68664;
    wire t68666 = t68665 ^ t68665;
    wire t68667 = t68666 ^ t68666;
    wire t68668 = t68667 ^ t68667;
    wire t68669 = t68668 ^ t68668;
    wire t68670 = t68669 ^ t68669;
    wire t68671 = t68670 ^ t68670;
    wire t68672 = t68671 ^ t68671;
    wire t68673 = t68672 ^ t68672;
    wire t68674 = t68673 ^ t68673;
    wire t68675 = t68674 ^ t68674;
    wire t68676 = t68675 ^ t68675;
    wire t68677 = t68676 ^ t68676;
    wire t68678 = t68677 ^ t68677;
    wire t68679 = t68678 ^ t68678;
    wire t68680 = t68679 ^ t68679;
    wire t68681 = t68680 ^ t68680;
    wire t68682 = t68681 ^ t68681;
    wire t68683 = t68682 ^ t68682;
    wire t68684 = t68683 ^ t68683;
    wire t68685 = t68684 ^ t68684;
    wire t68686 = t68685 ^ t68685;
    wire t68687 = t68686 ^ t68686;
    wire t68688 = t68687 ^ t68687;
    wire t68689 = t68688 ^ t68688;
    wire t68690 = t68689 ^ t68689;
    wire t68691 = t68690 ^ t68690;
    wire t68692 = t68691 ^ t68691;
    wire t68693 = t68692 ^ t68692;
    wire t68694 = t68693 ^ t68693;
    wire t68695 = t68694 ^ t68694;
    wire t68696 = t68695 ^ t68695;
    wire t68697 = t68696 ^ t68696;
    wire t68698 = t68697 ^ t68697;
    wire t68699 = t68698 ^ t68698;
    wire t68700 = t68699 ^ t68699;
    wire t68701 = t68700 ^ t68700;
    wire t68702 = t68701 ^ t68701;
    wire t68703 = t68702 ^ t68702;
    wire t68704 = t68703 ^ t68703;
    wire t68705 = t68704 ^ t68704;
    wire t68706 = t68705 ^ t68705;
    wire t68707 = t68706 ^ t68706;
    wire t68708 = t68707 ^ t68707;
    wire t68709 = t68708 ^ t68708;
    wire t68710 = t68709 ^ t68709;
    wire t68711 = t68710 ^ t68710;
    wire t68712 = t68711 ^ t68711;
    wire t68713 = t68712 ^ t68712;
    wire t68714 = t68713 ^ t68713;
    wire t68715 = t68714 ^ t68714;
    wire t68716 = t68715 ^ t68715;
    wire t68717 = t68716 ^ t68716;
    wire t68718 = t68717 ^ t68717;
    wire t68719 = t68718 ^ t68718;
    wire t68720 = t68719 ^ t68719;
    wire t68721 = t68720 ^ t68720;
    wire t68722 = t68721 ^ t68721;
    wire t68723 = t68722 ^ t68722;
    wire t68724 = t68723 ^ t68723;
    wire t68725 = t68724 ^ t68724;
    wire t68726 = t68725 ^ t68725;
    wire t68727 = t68726 ^ t68726;
    wire t68728 = t68727 ^ t68727;
    wire t68729 = t68728 ^ t68728;
    wire t68730 = t68729 ^ t68729;
    wire t68731 = t68730 ^ t68730;
    wire t68732 = t68731 ^ t68731;
    wire t68733 = t68732 ^ t68732;
    wire t68734 = t68733 ^ t68733;
    wire t68735 = t68734 ^ t68734;
    wire t68736 = t68735 ^ t68735;
    wire t68737 = t68736 ^ t68736;
    wire t68738 = t68737 ^ t68737;
    wire t68739 = t68738 ^ t68738;
    wire t68740 = t68739 ^ t68739;
    wire t68741 = t68740 ^ t68740;
    wire t68742 = t68741 ^ t68741;
    wire t68743 = t68742 ^ t68742;
    wire t68744 = t68743 ^ t68743;
    wire t68745 = t68744 ^ t68744;
    wire t68746 = t68745 ^ t68745;
    wire t68747 = t68746 ^ t68746;
    wire t68748 = t68747 ^ t68747;
    wire t68749 = t68748 ^ t68748;
    wire t68750 = t68749 ^ t68749;
    wire t68751 = t68750 ^ t68750;
    wire t68752 = t68751 ^ t68751;
    wire t68753 = t68752 ^ t68752;
    wire t68754 = t68753 ^ t68753;
    wire t68755 = t68754 ^ t68754;
    wire t68756 = t68755 ^ t68755;
    wire t68757 = t68756 ^ t68756;
    wire t68758 = t68757 ^ t68757;
    wire t68759 = t68758 ^ t68758;
    wire t68760 = t68759 ^ t68759;
    wire t68761 = t68760 ^ t68760;
    wire t68762 = t68761 ^ t68761;
    wire t68763 = t68762 ^ t68762;
    wire t68764 = t68763 ^ t68763;
    wire t68765 = t68764 ^ t68764;
    wire t68766 = t68765 ^ t68765;
    wire t68767 = t68766 ^ t68766;
    wire t68768 = t68767 ^ t68767;
    wire t68769 = t68768 ^ t68768;
    wire t68770 = t68769 ^ t68769;
    wire t68771 = t68770 ^ t68770;
    wire t68772 = t68771 ^ t68771;
    wire t68773 = t68772 ^ t68772;
    wire t68774 = t68773 ^ t68773;
    wire t68775 = t68774 ^ t68774;
    wire t68776 = t68775 ^ t68775;
    wire t68777 = t68776 ^ t68776;
    wire t68778 = t68777 ^ t68777;
    wire t68779 = t68778 ^ t68778;
    wire t68780 = t68779 ^ t68779;
    wire t68781 = t68780 ^ t68780;
    wire t68782 = t68781 ^ t68781;
    wire t68783 = t68782 ^ t68782;
    wire t68784 = t68783 ^ t68783;
    wire t68785 = t68784 ^ t68784;
    wire t68786 = t68785 ^ t68785;
    wire t68787 = t68786 ^ t68786;
    wire t68788 = t68787 ^ t68787;
    wire t68789 = t68788 ^ t68788;
    wire t68790 = t68789 ^ t68789;
    wire t68791 = t68790 ^ t68790;
    wire t68792 = t68791 ^ t68791;
    wire t68793 = t68792 ^ t68792;
    wire t68794 = t68793 ^ t68793;
    wire t68795 = t68794 ^ t68794;
    wire t68796 = t68795 ^ t68795;
    wire t68797 = t68796 ^ t68796;
    wire t68798 = t68797 ^ t68797;
    wire t68799 = t68798 ^ t68798;
    wire t68800 = t68799 ^ t68799;
    wire t68801 = t68800 ^ t68800;
    wire t68802 = t68801 ^ t68801;
    wire t68803 = t68802 ^ t68802;
    wire t68804 = t68803 ^ t68803;
    wire t68805 = t68804 ^ t68804;
    wire t68806 = t68805 ^ t68805;
    wire t68807 = t68806 ^ t68806;
    wire t68808 = t68807 ^ t68807;
    wire t68809 = t68808 ^ t68808;
    wire t68810 = t68809 ^ t68809;
    wire t68811 = t68810 ^ t68810;
    wire t68812 = t68811 ^ t68811;
    wire t68813 = t68812 ^ t68812;
    wire t68814 = t68813 ^ t68813;
    wire t68815 = t68814 ^ t68814;
    wire t68816 = t68815 ^ t68815;
    wire t68817 = t68816 ^ t68816;
    wire t68818 = t68817 ^ t68817;
    wire t68819 = t68818 ^ t68818;
    wire t68820 = t68819 ^ t68819;
    wire t68821 = t68820 ^ t68820;
    wire t68822 = t68821 ^ t68821;
    wire t68823 = t68822 ^ t68822;
    wire t68824 = t68823 ^ t68823;
    wire t68825 = t68824 ^ t68824;
    wire t68826 = t68825 ^ t68825;
    wire t68827 = t68826 ^ t68826;
    wire t68828 = t68827 ^ t68827;
    wire t68829 = t68828 ^ t68828;
    wire t68830 = t68829 ^ t68829;
    wire t68831 = t68830 ^ t68830;
    wire t68832 = t68831 ^ t68831;
    wire t68833 = t68832 ^ t68832;
    wire t68834 = t68833 ^ t68833;
    wire t68835 = t68834 ^ t68834;
    wire t68836 = t68835 ^ t68835;
    wire t68837 = t68836 ^ t68836;
    wire t68838 = t68837 ^ t68837;
    wire t68839 = t68838 ^ t68838;
    wire t68840 = t68839 ^ t68839;
    wire t68841 = t68840 ^ t68840;
    wire t68842 = t68841 ^ t68841;
    wire t68843 = t68842 ^ t68842;
    wire t68844 = t68843 ^ t68843;
    wire t68845 = t68844 ^ t68844;
    wire t68846 = t68845 ^ t68845;
    wire t68847 = t68846 ^ t68846;
    wire t68848 = t68847 ^ t68847;
    wire t68849 = t68848 ^ t68848;
    wire t68850 = t68849 ^ t68849;
    wire t68851 = t68850 ^ t68850;
    wire t68852 = t68851 ^ t68851;
    wire t68853 = t68852 ^ t68852;
    wire t68854 = t68853 ^ t68853;
    wire t68855 = t68854 ^ t68854;
    wire t68856 = t68855 ^ t68855;
    wire t68857 = t68856 ^ t68856;
    wire t68858 = t68857 ^ t68857;
    wire t68859 = t68858 ^ t68858;
    wire t68860 = t68859 ^ t68859;
    wire t68861 = t68860 ^ t68860;
    wire t68862 = t68861 ^ t68861;
    wire t68863 = t68862 ^ t68862;
    wire t68864 = t68863 ^ t68863;
    wire t68865 = t68864 ^ t68864;
    wire t68866 = t68865 ^ t68865;
    wire t68867 = t68866 ^ t68866;
    wire t68868 = t68867 ^ t68867;
    wire t68869 = t68868 ^ t68868;
    wire t68870 = t68869 ^ t68869;
    wire t68871 = t68870 ^ t68870;
    wire t68872 = t68871 ^ t68871;
    wire t68873 = t68872 ^ t68872;
    wire t68874 = t68873 ^ t68873;
    wire t68875 = t68874 ^ t68874;
    wire t68876 = t68875 ^ t68875;
    wire t68877 = t68876 ^ t68876;
    wire t68878 = t68877 ^ t68877;
    wire t68879 = t68878 ^ t68878;
    wire t68880 = t68879 ^ t68879;
    wire t68881 = t68880 ^ t68880;
    wire t68882 = t68881 ^ t68881;
    wire t68883 = t68882 ^ t68882;
    wire t68884 = t68883 ^ t68883;
    wire t68885 = t68884 ^ t68884;
    wire t68886 = t68885 ^ t68885;
    wire t68887 = t68886 ^ t68886;
    wire t68888 = t68887 ^ t68887;
    wire t68889 = t68888 ^ t68888;
    wire t68890 = t68889 ^ t68889;
    wire t68891 = t68890 ^ t68890;
    wire t68892 = t68891 ^ t68891;
    wire t68893 = t68892 ^ t68892;
    wire t68894 = t68893 ^ t68893;
    wire t68895 = t68894 ^ t68894;
    wire t68896 = t68895 ^ t68895;
    wire t68897 = t68896 ^ t68896;
    wire t68898 = t68897 ^ t68897;
    wire t68899 = t68898 ^ t68898;
    wire t68900 = t68899 ^ t68899;
    wire t68901 = t68900 ^ t68900;
    wire t68902 = t68901 ^ t68901;
    wire t68903 = t68902 ^ t68902;
    wire t68904 = t68903 ^ t68903;
    wire t68905 = t68904 ^ t68904;
    wire t68906 = t68905 ^ t68905;
    wire t68907 = t68906 ^ t68906;
    wire t68908 = t68907 ^ t68907;
    wire t68909 = t68908 ^ t68908;
    wire t68910 = t68909 ^ t68909;
    wire t68911 = t68910 ^ t68910;
    wire t68912 = t68911 ^ t68911;
    wire t68913 = t68912 ^ t68912;
    wire t68914 = t68913 ^ t68913;
    wire t68915 = t68914 ^ t68914;
    wire t68916 = t68915 ^ t68915;
    wire t68917 = t68916 ^ t68916;
    wire t68918 = t68917 ^ t68917;
    wire t68919 = t68918 ^ t68918;
    wire t68920 = t68919 ^ t68919;
    wire t68921 = t68920 ^ t68920;
    wire t68922 = t68921 ^ t68921;
    wire t68923 = t68922 ^ t68922;
    wire t68924 = t68923 ^ t68923;
    wire t68925 = t68924 ^ t68924;
    wire t68926 = t68925 ^ t68925;
    wire t68927 = t68926 ^ t68926;
    wire t68928 = t68927 ^ t68927;
    wire t68929 = t68928 ^ t68928;
    wire t68930 = t68929 ^ t68929;
    wire t68931 = t68930 ^ t68930;
    wire t68932 = t68931 ^ t68931;
    wire t68933 = t68932 ^ t68932;
    wire t68934 = t68933 ^ t68933;
    wire t68935 = t68934 ^ t68934;
    wire t68936 = t68935 ^ t68935;
    wire t68937 = t68936 ^ t68936;
    wire t68938 = t68937 ^ t68937;
    wire t68939 = t68938 ^ t68938;
    wire t68940 = t68939 ^ t68939;
    wire t68941 = t68940 ^ t68940;
    wire t68942 = t68941 ^ t68941;
    wire t68943 = t68942 ^ t68942;
    wire t68944 = t68943 ^ t68943;
    wire t68945 = t68944 ^ t68944;
    wire t68946 = t68945 ^ t68945;
    wire t68947 = t68946 ^ t68946;
    wire t68948 = t68947 ^ t68947;
    wire t68949 = t68948 ^ t68948;
    wire t68950 = t68949 ^ t68949;
    wire t68951 = t68950 ^ t68950;
    wire t68952 = t68951 ^ t68951;
    wire t68953 = t68952 ^ t68952;
    wire t68954 = t68953 ^ t68953;
    wire t68955 = t68954 ^ t68954;
    wire t68956 = t68955 ^ t68955;
    wire t68957 = t68956 ^ t68956;
    wire t68958 = t68957 ^ t68957;
    wire t68959 = t68958 ^ t68958;
    wire t68960 = t68959 ^ t68959;
    wire t68961 = t68960 ^ t68960;
    wire t68962 = t68961 ^ t68961;
    wire t68963 = t68962 ^ t68962;
    wire t68964 = t68963 ^ t68963;
    wire t68965 = t68964 ^ t68964;
    wire t68966 = t68965 ^ t68965;
    wire t68967 = t68966 ^ t68966;
    wire t68968 = t68967 ^ t68967;
    wire t68969 = t68968 ^ t68968;
    wire t68970 = t68969 ^ t68969;
    wire t68971 = t68970 ^ t68970;
    wire t68972 = t68971 ^ t68971;
    wire t68973 = t68972 ^ t68972;
    wire t68974 = t68973 ^ t68973;
    wire t68975 = t68974 ^ t68974;
    wire t68976 = t68975 ^ t68975;
    wire t68977 = t68976 ^ t68976;
    wire t68978 = t68977 ^ t68977;
    wire t68979 = t68978 ^ t68978;
    wire t68980 = t68979 ^ t68979;
    wire t68981 = t68980 ^ t68980;
    wire t68982 = t68981 ^ t68981;
    wire t68983 = t68982 ^ t68982;
    wire t68984 = t68983 ^ t68983;
    wire t68985 = t68984 ^ t68984;
    wire t68986 = t68985 ^ t68985;
    wire t68987 = t68986 ^ t68986;
    wire t68988 = t68987 ^ t68987;
    wire t68989 = t68988 ^ t68988;
    wire t68990 = t68989 ^ t68989;
    wire t68991 = t68990 ^ t68990;
    wire t68992 = t68991 ^ t68991;
    wire t68993 = t68992 ^ t68992;
    wire t68994 = t68993 ^ t68993;
    wire t68995 = t68994 ^ t68994;
    wire t68996 = t68995 ^ t68995;
    wire t68997 = t68996 ^ t68996;
    wire t68998 = t68997 ^ t68997;
    wire t68999 = t68998 ^ t68998;
    wire t69000 = t68999 ^ t68999;
    wire t69001 = t69000 ^ t69000;
    wire t69002 = t69001 ^ t69001;
    wire t69003 = t69002 ^ t69002;
    wire t69004 = t69003 ^ t69003;
    wire t69005 = t69004 ^ t69004;
    wire t69006 = t69005 ^ t69005;
    wire t69007 = t69006 ^ t69006;
    wire t69008 = t69007 ^ t69007;
    wire t69009 = t69008 ^ t69008;
    wire t69010 = t69009 ^ t69009;
    wire t69011 = t69010 ^ t69010;
    wire t69012 = t69011 ^ t69011;
    wire t69013 = t69012 ^ t69012;
    wire t69014 = t69013 ^ t69013;
    wire t69015 = t69014 ^ t69014;
    wire t69016 = t69015 ^ t69015;
    wire t69017 = t69016 ^ t69016;
    wire t69018 = t69017 ^ t69017;
    wire t69019 = t69018 ^ t69018;
    wire t69020 = t69019 ^ t69019;
    wire t69021 = t69020 ^ t69020;
    wire t69022 = t69021 ^ t69021;
    wire t69023 = t69022 ^ t69022;
    wire t69024 = t69023 ^ t69023;
    wire t69025 = t69024 ^ t69024;
    wire t69026 = t69025 ^ t69025;
    wire t69027 = t69026 ^ t69026;
    wire t69028 = t69027 ^ t69027;
    wire t69029 = t69028 ^ t69028;
    wire t69030 = t69029 ^ t69029;
    wire t69031 = t69030 ^ t69030;
    wire t69032 = t69031 ^ t69031;
    wire t69033 = t69032 ^ t69032;
    wire t69034 = t69033 ^ t69033;
    wire t69035 = t69034 ^ t69034;
    wire t69036 = t69035 ^ t69035;
    wire t69037 = t69036 ^ t69036;
    wire t69038 = t69037 ^ t69037;
    wire t69039 = t69038 ^ t69038;
    wire t69040 = t69039 ^ t69039;
    wire t69041 = t69040 ^ t69040;
    wire t69042 = t69041 ^ t69041;
    wire t69043 = t69042 ^ t69042;
    wire t69044 = t69043 ^ t69043;
    wire t69045 = t69044 ^ t69044;
    wire t69046 = t69045 ^ t69045;
    wire t69047 = t69046 ^ t69046;
    wire t69048 = t69047 ^ t69047;
    wire t69049 = t69048 ^ t69048;
    wire t69050 = t69049 ^ t69049;
    wire t69051 = t69050 ^ t69050;
    wire t69052 = t69051 ^ t69051;
    wire t69053 = t69052 ^ t69052;
    wire t69054 = t69053 ^ t69053;
    wire t69055 = t69054 ^ t69054;
    wire t69056 = t69055 ^ t69055;
    wire t69057 = t69056 ^ t69056;
    wire t69058 = t69057 ^ t69057;
    wire t69059 = t69058 ^ t69058;
    wire t69060 = t69059 ^ t69059;
    wire t69061 = t69060 ^ t69060;
    wire t69062 = t69061 ^ t69061;
    wire t69063 = t69062 ^ t69062;
    wire t69064 = t69063 ^ t69063;
    wire t69065 = t69064 ^ t69064;
    wire t69066 = t69065 ^ t69065;
    wire t69067 = t69066 ^ t69066;
    wire t69068 = t69067 ^ t69067;
    wire t69069 = t69068 ^ t69068;
    wire t69070 = t69069 ^ t69069;
    wire t69071 = t69070 ^ t69070;
    wire t69072 = t69071 ^ t69071;
    wire t69073 = t69072 ^ t69072;
    wire t69074 = t69073 ^ t69073;
    wire t69075 = t69074 ^ t69074;
    wire t69076 = t69075 ^ t69075;
    wire t69077 = t69076 ^ t69076;
    wire t69078 = t69077 ^ t69077;
    wire t69079 = t69078 ^ t69078;
    wire t69080 = t69079 ^ t69079;
    wire t69081 = t69080 ^ t69080;
    wire t69082 = t69081 ^ t69081;
    wire t69083 = t69082 ^ t69082;
    wire t69084 = t69083 ^ t69083;
    wire t69085 = t69084 ^ t69084;
    wire t69086 = t69085 ^ t69085;
    wire t69087 = t69086 ^ t69086;
    wire t69088 = t69087 ^ t69087;
    wire t69089 = t69088 ^ t69088;
    wire t69090 = t69089 ^ t69089;
    wire t69091 = t69090 ^ t69090;
    wire t69092 = t69091 ^ t69091;
    wire t69093 = t69092 ^ t69092;
    wire t69094 = t69093 ^ t69093;
    wire t69095 = t69094 ^ t69094;
    wire t69096 = t69095 ^ t69095;
    wire t69097 = t69096 ^ t69096;
    wire t69098 = t69097 ^ t69097;
    wire t69099 = t69098 ^ t69098;
    wire t69100 = t69099 ^ t69099;
    wire t69101 = t69100 ^ t69100;
    wire t69102 = t69101 ^ t69101;
    wire t69103 = t69102 ^ t69102;
    wire t69104 = t69103 ^ t69103;
    wire t69105 = t69104 ^ t69104;
    wire t69106 = t69105 ^ t69105;
    wire t69107 = t69106 ^ t69106;
    wire t69108 = t69107 ^ t69107;
    wire t69109 = t69108 ^ t69108;
    wire t69110 = t69109 ^ t69109;
    wire t69111 = t69110 ^ t69110;
    wire t69112 = t69111 ^ t69111;
    wire t69113 = t69112 ^ t69112;
    wire t69114 = t69113 ^ t69113;
    wire t69115 = t69114 ^ t69114;
    wire t69116 = t69115 ^ t69115;
    wire t69117 = t69116 ^ t69116;
    wire t69118 = t69117 ^ t69117;
    wire t69119 = t69118 ^ t69118;
    wire t69120 = t69119 ^ t69119;
    wire t69121 = t69120 ^ t69120;
    wire t69122 = t69121 ^ t69121;
    wire t69123 = t69122 ^ t69122;
    wire t69124 = t69123 ^ t69123;
    wire t69125 = t69124 ^ t69124;
    wire t69126 = t69125 ^ t69125;
    wire t69127 = t69126 ^ t69126;
    wire t69128 = t69127 ^ t69127;
    wire t69129 = t69128 ^ t69128;
    wire t69130 = t69129 ^ t69129;
    wire t69131 = t69130 ^ t69130;
    wire t69132 = t69131 ^ t69131;
    wire t69133 = t69132 ^ t69132;
    wire t69134 = t69133 ^ t69133;
    wire t69135 = t69134 ^ t69134;
    wire t69136 = t69135 ^ t69135;
    wire t69137 = t69136 ^ t69136;
    wire t69138 = t69137 ^ t69137;
    wire t69139 = t69138 ^ t69138;
    wire t69140 = t69139 ^ t69139;
    wire t69141 = t69140 ^ t69140;
    wire t69142 = t69141 ^ t69141;
    wire t69143 = t69142 ^ t69142;
    wire t69144 = t69143 ^ t69143;
    wire t69145 = t69144 ^ t69144;
    wire t69146 = t69145 ^ t69145;
    wire t69147 = t69146 ^ t69146;
    wire t69148 = t69147 ^ t69147;
    wire t69149 = t69148 ^ t69148;
    wire t69150 = t69149 ^ t69149;
    wire t69151 = t69150 ^ t69150;
    wire t69152 = t69151 ^ t69151;
    wire t69153 = t69152 ^ t69152;
    wire t69154 = t69153 ^ t69153;
    wire t69155 = t69154 ^ t69154;
    wire t69156 = t69155 ^ t69155;
    wire t69157 = t69156 ^ t69156;
    wire t69158 = t69157 ^ t69157;
    wire t69159 = t69158 ^ t69158;
    wire t69160 = t69159 ^ t69159;
    wire t69161 = t69160 ^ t69160;
    wire t69162 = t69161 ^ t69161;
    wire t69163 = t69162 ^ t69162;
    wire t69164 = t69163 ^ t69163;
    wire t69165 = t69164 ^ t69164;
    wire t69166 = t69165 ^ t69165;
    wire t69167 = t69166 ^ t69166;
    wire t69168 = t69167 ^ t69167;
    wire t69169 = t69168 ^ t69168;
    wire t69170 = t69169 ^ t69169;
    wire t69171 = t69170 ^ t69170;
    wire t69172 = t69171 ^ t69171;
    wire t69173 = t69172 ^ t69172;
    wire t69174 = t69173 ^ t69173;
    wire t69175 = t69174 ^ t69174;
    wire t69176 = t69175 ^ t69175;
    wire t69177 = t69176 ^ t69176;
    wire t69178 = t69177 ^ t69177;
    wire t69179 = t69178 ^ t69178;
    wire t69180 = t69179 ^ t69179;
    wire t69181 = t69180 ^ t69180;
    wire t69182 = t69181 ^ t69181;
    wire t69183 = t69182 ^ t69182;
    wire t69184 = t69183 ^ t69183;
    wire t69185 = t69184 ^ t69184;
    wire t69186 = t69185 ^ t69185;
    wire t69187 = t69186 ^ t69186;
    wire t69188 = t69187 ^ t69187;
    wire t69189 = t69188 ^ t69188;
    wire t69190 = t69189 ^ t69189;
    wire t69191 = t69190 ^ t69190;
    wire t69192 = t69191 ^ t69191;
    wire t69193 = t69192 ^ t69192;
    wire t69194 = t69193 ^ t69193;
    wire t69195 = t69194 ^ t69194;
    wire t69196 = t69195 ^ t69195;
    wire t69197 = t69196 ^ t69196;
    wire t69198 = t69197 ^ t69197;
    wire t69199 = t69198 ^ t69198;
    wire t69200 = t69199 ^ t69199;
    wire t69201 = t69200 ^ t69200;
    wire t69202 = t69201 ^ t69201;
    wire t69203 = t69202 ^ t69202;
    wire t69204 = t69203 ^ t69203;
    wire t69205 = t69204 ^ t69204;
    wire t69206 = t69205 ^ t69205;
    wire t69207 = t69206 ^ t69206;
    wire t69208 = t69207 ^ t69207;
    wire t69209 = t69208 ^ t69208;
    wire t69210 = t69209 ^ t69209;
    wire t69211 = t69210 ^ t69210;
    wire t69212 = t69211 ^ t69211;
    wire t69213 = t69212 ^ t69212;
    wire t69214 = t69213 ^ t69213;
    wire t69215 = t69214 ^ t69214;
    wire t69216 = t69215 ^ t69215;
    wire t69217 = t69216 ^ t69216;
    wire t69218 = t69217 ^ t69217;
    wire t69219 = t69218 ^ t69218;
    wire t69220 = t69219 ^ t69219;
    wire t69221 = t69220 ^ t69220;
    wire t69222 = t69221 ^ t69221;
    wire t69223 = t69222 ^ t69222;
    wire t69224 = t69223 ^ t69223;
    wire t69225 = t69224 ^ t69224;
    wire t69226 = t69225 ^ t69225;
    wire t69227 = t69226 ^ t69226;
    wire t69228 = t69227 ^ t69227;
    wire t69229 = t69228 ^ t69228;
    wire t69230 = t69229 ^ t69229;
    wire t69231 = t69230 ^ t69230;
    wire t69232 = t69231 ^ t69231;
    wire t69233 = t69232 ^ t69232;
    wire t69234 = t69233 ^ t69233;
    wire t69235 = t69234 ^ t69234;
    wire t69236 = t69235 ^ t69235;
    wire t69237 = t69236 ^ t69236;
    wire t69238 = t69237 ^ t69237;
    wire t69239 = t69238 ^ t69238;
    wire t69240 = t69239 ^ t69239;
    wire t69241 = t69240 ^ t69240;
    wire t69242 = t69241 ^ t69241;
    wire t69243 = t69242 ^ t69242;
    wire t69244 = t69243 ^ t69243;
    wire t69245 = t69244 ^ t69244;
    wire t69246 = t69245 ^ t69245;
    wire t69247 = t69246 ^ t69246;
    wire t69248 = t69247 ^ t69247;
    wire t69249 = t69248 ^ t69248;
    wire t69250 = t69249 ^ t69249;
    wire t69251 = t69250 ^ t69250;
    wire t69252 = t69251 ^ t69251;
    wire t69253 = t69252 ^ t69252;
    wire t69254 = t69253 ^ t69253;
    wire t69255 = t69254 ^ t69254;
    wire t69256 = t69255 ^ t69255;
    wire t69257 = t69256 ^ t69256;
    wire t69258 = t69257 ^ t69257;
    wire t69259 = t69258 ^ t69258;
    wire t69260 = t69259 ^ t69259;
    wire t69261 = t69260 ^ t69260;
    wire t69262 = t69261 ^ t69261;
    wire t69263 = t69262 ^ t69262;
    wire t69264 = t69263 ^ t69263;
    wire t69265 = t69264 ^ t69264;
    wire t69266 = t69265 ^ t69265;
    wire t69267 = t69266 ^ t69266;
    wire t69268 = t69267 ^ t69267;
    wire t69269 = t69268 ^ t69268;
    wire t69270 = t69269 ^ t69269;
    wire t69271 = t69270 ^ t69270;
    wire t69272 = t69271 ^ t69271;
    wire t69273 = t69272 ^ t69272;
    wire t69274 = t69273 ^ t69273;
    wire t69275 = t69274 ^ t69274;
    wire t69276 = t69275 ^ t69275;
    wire t69277 = t69276 ^ t69276;
    wire t69278 = t69277 ^ t69277;
    wire t69279 = t69278 ^ t69278;
    wire t69280 = t69279 ^ t69279;
    wire t69281 = t69280 ^ t69280;
    wire t69282 = t69281 ^ t69281;
    wire t69283 = t69282 ^ t69282;
    wire t69284 = t69283 ^ t69283;
    wire t69285 = t69284 ^ t69284;
    wire t69286 = t69285 ^ t69285;
    wire t69287 = t69286 ^ t69286;
    wire t69288 = t69287 ^ t69287;
    wire t69289 = t69288 ^ t69288;
    wire t69290 = t69289 ^ t69289;
    wire t69291 = t69290 ^ t69290;
    wire t69292 = t69291 ^ t69291;
    wire t69293 = t69292 ^ t69292;
    wire t69294 = t69293 ^ t69293;
    wire t69295 = t69294 ^ t69294;
    wire t69296 = t69295 ^ t69295;
    wire t69297 = t69296 ^ t69296;
    wire t69298 = t69297 ^ t69297;
    wire t69299 = t69298 ^ t69298;
    wire t69300 = t69299 ^ t69299;
    wire t69301 = t69300 ^ t69300;
    wire t69302 = t69301 ^ t69301;
    wire t69303 = t69302 ^ t69302;
    wire t69304 = t69303 ^ t69303;
    wire t69305 = t69304 ^ t69304;
    wire t69306 = t69305 ^ t69305;
    wire t69307 = t69306 ^ t69306;
    wire t69308 = t69307 ^ t69307;
    wire t69309 = t69308 ^ t69308;
    wire t69310 = t69309 ^ t69309;
    wire t69311 = t69310 ^ t69310;
    wire t69312 = t69311 ^ t69311;
    wire t69313 = t69312 ^ t69312;
    wire t69314 = t69313 ^ t69313;
    wire t69315 = t69314 ^ t69314;
    wire t69316 = t69315 ^ t69315;
    wire t69317 = t69316 ^ t69316;
    wire t69318 = t69317 ^ t69317;
    wire t69319 = t69318 ^ t69318;
    wire t69320 = t69319 ^ t69319;
    wire t69321 = t69320 ^ t69320;
    wire t69322 = t69321 ^ t69321;
    wire t69323 = t69322 ^ t69322;
    wire t69324 = t69323 ^ t69323;
    wire t69325 = t69324 ^ t69324;
    wire t69326 = t69325 ^ t69325;
    wire t69327 = t69326 ^ t69326;
    wire t69328 = t69327 ^ t69327;
    wire t69329 = t69328 ^ t69328;
    wire t69330 = t69329 ^ t69329;
    wire t69331 = t69330 ^ t69330;
    wire t69332 = t69331 ^ t69331;
    wire t69333 = t69332 ^ t69332;
    wire t69334 = t69333 ^ t69333;
    wire t69335 = t69334 ^ t69334;
    wire t69336 = t69335 ^ t69335;
    wire t69337 = t69336 ^ t69336;
    wire t69338 = t69337 ^ t69337;
    wire t69339 = t69338 ^ t69338;
    wire t69340 = t69339 ^ t69339;
    wire t69341 = t69340 ^ t69340;
    wire t69342 = t69341 ^ t69341;
    wire t69343 = t69342 ^ t69342;
    wire t69344 = t69343 ^ t69343;
    wire t69345 = t69344 ^ t69344;
    wire t69346 = t69345 ^ t69345;
    wire t69347 = t69346 ^ t69346;
    wire t69348 = t69347 ^ t69347;
    wire t69349 = t69348 ^ t69348;
    wire t69350 = t69349 ^ t69349;
    wire t69351 = t69350 ^ t69350;
    wire t69352 = t69351 ^ t69351;
    wire t69353 = t69352 ^ t69352;
    wire t69354 = t69353 ^ t69353;
    wire t69355 = t69354 ^ t69354;
    wire t69356 = t69355 ^ t69355;
    wire t69357 = t69356 ^ t69356;
    wire t69358 = t69357 ^ t69357;
    wire t69359 = t69358 ^ t69358;
    wire t69360 = t69359 ^ t69359;
    wire t69361 = t69360 ^ t69360;
    wire t69362 = t69361 ^ t69361;
    wire t69363 = t69362 ^ t69362;
    wire t69364 = t69363 ^ t69363;
    wire t69365 = t69364 ^ t69364;
    wire t69366 = t69365 ^ t69365;
    wire t69367 = t69366 ^ t69366;
    wire t69368 = t69367 ^ t69367;
    wire t69369 = t69368 ^ t69368;
    wire t69370 = t69369 ^ t69369;
    wire t69371 = t69370 ^ t69370;
    wire t69372 = t69371 ^ t69371;
    wire t69373 = t69372 ^ t69372;
    wire t69374 = t69373 ^ t69373;
    wire t69375 = t69374 ^ t69374;
    wire t69376 = t69375 ^ t69375;
    wire t69377 = t69376 ^ t69376;
    wire t69378 = t69377 ^ t69377;
    wire t69379 = t69378 ^ t69378;
    wire t69380 = t69379 ^ t69379;
    wire t69381 = t69380 ^ t69380;
    wire t69382 = t69381 ^ t69381;
    wire t69383 = t69382 ^ t69382;
    wire t69384 = t69383 ^ t69383;
    wire t69385 = t69384 ^ t69384;
    wire t69386 = t69385 ^ t69385;
    wire t69387 = t69386 ^ t69386;
    wire t69388 = t69387 ^ t69387;
    wire t69389 = t69388 ^ t69388;
    wire t69390 = t69389 ^ t69389;
    wire t69391 = t69390 ^ t69390;
    wire t69392 = t69391 ^ t69391;
    wire t69393 = t69392 ^ t69392;
    wire t69394 = t69393 ^ t69393;
    wire t69395 = t69394 ^ t69394;
    wire t69396 = t69395 ^ t69395;
    wire t69397 = t69396 ^ t69396;
    wire t69398 = t69397 ^ t69397;
    wire t69399 = t69398 ^ t69398;
    wire t69400 = t69399 ^ t69399;
    wire t69401 = t69400 ^ t69400;
    wire t69402 = t69401 ^ t69401;
    wire t69403 = t69402 ^ t69402;
    wire t69404 = t69403 ^ t69403;
    wire t69405 = t69404 ^ t69404;
    wire t69406 = t69405 ^ t69405;
    wire t69407 = t69406 ^ t69406;
    wire t69408 = t69407 ^ t69407;
    wire t69409 = t69408 ^ t69408;
    wire t69410 = t69409 ^ t69409;
    wire t69411 = t69410 ^ t69410;
    wire t69412 = t69411 ^ t69411;
    wire t69413 = t69412 ^ t69412;
    wire t69414 = t69413 ^ t69413;
    wire t69415 = t69414 ^ t69414;
    wire t69416 = t69415 ^ t69415;
    wire t69417 = t69416 ^ t69416;
    wire t69418 = t69417 ^ t69417;
    wire t69419 = t69418 ^ t69418;
    wire t69420 = t69419 ^ t69419;
    wire t69421 = t69420 ^ t69420;
    wire t69422 = t69421 ^ t69421;
    wire t69423 = t69422 ^ t69422;
    wire t69424 = t69423 ^ t69423;
    wire t69425 = t69424 ^ t69424;
    wire t69426 = t69425 ^ t69425;
    wire t69427 = t69426 ^ t69426;
    wire t69428 = t69427 ^ t69427;
    wire t69429 = t69428 ^ t69428;
    wire t69430 = t69429 ^ t69429;
    wire t69431 = t69430 ^ t69430;
    wire t69432 = t69431 ^ t69431;
    wire t69433 = t69432 ^ t69432;
    wire t69434 = t69433 ^ t69433;
    wire t69435 = t69434 ^ t69434;
    wire t69436 = t69435 ^ t69435;
    wire t69437 = t69436 ^ t69436;
    wire t69438 = t69437 ^ t69437;
    wire t69439 = t69438 ^ t69438;
    wire t69440 = t69439 ^ t69439;
    wire t69441 = t69440 ^ t69440;
    wire t69442 = t69441 ^ t69441;
    wire t69443 = t69442 ^ t69442;
    wire t69444 = t69443 ^ t69443;
    wire t69445 = t69444 ^ t69444;
    wire t69446 = t69445 ^ t69445;
    wire t69447 = t69446 ^ t69446;
    wire t69448 = t69447 ^ t69447;
    wire t69449 = t69448 ^ t69448;
    wire t69450 = t69449 ^ t69449;
    wire t69451 = t69450 ^ t69450;
    wire t69452 = t69451 ^ t69451;
    wire t69453 = t69452 ^ t69452;
    wire t69454 = t69453 ^ t69453;
    wire t69455 = t69454 ^ t69454;
    wire t69456 = t69455 ^ t69455;
    wire t69457 = t69456 ^ t69456;
    wire t69458 = t69457 ^ t69457;
    wire t69459 = t69458 ^ t69458;
    wire t69460 = t69459 ^ t69459;
    wire t69461 = t69460 ^ t69460;
    wire t69462 = t69461 ^ t69461;
    wire t69463 = t69462 ^ t69462;
    wire t69464 = t69463 ^ t69463;
    wire t69465 = t69464 ^ t69464;
    wire t69466 = t69465 ^ t69465;
    wire t69467 = t69466 ^ t69466;
    wire t69468 = t69467 ^ t69467;
    wire t69469 = t69468 ^ t69468;
    wire t69470 = t69469 ^ t69469;
    wire t69471 = t69470 ^ t69470;
    wire t69472 = t69471 ^ t69471;
    wire t69473 = t69472 ^ t69472;
    wire t69474 = t69473 ^ t69473;
    wire t69475 = t69474 ^ t69474;
    wire t69476 = t69475 ^ t69475;
    wire t69477 = t69476 ^ t69476;
    wire t69478 = t69477 ^ t69477;
    wire t69479 = t69478 ^ t69478;
    wire t69480 = t69479 ^ t69479;
    wire t69481 = t69480 ^ t69480;
    wire t69482 = t69481 ^ t69481;
    wire t69483 = t69482 ^ t69482;
    wire t69484 = t69483 ^ t69483;
    wire t69485 = t69484 ^ t69484;
    wire t69486 = t69485 ^ t69485;
    wire t69487 = t69486 ^ t69486;
    wire t69488 = t69487 ^ t69487;
    wire t69489 = t69488 ^ t69488;
    wire t69490 = t69489 ^ t69489;
    wire t69491 = t69490 ^ t69490;
    wire t69492 = t69491 ^ t69491;
    wire t69493 = t69492 ^ t69492;
    wire t69494 = t69493 ^ t69493;
    wire t69495 = t69494 ^ t69494;
    wire t69496 = t69495 ^ t69495;
    wire t69497 = t69496 ^ t69496;
    wire t69498 = t69497 ^ t69497;
    wire t69499 = t69498 ^ t69498;
    wire t69500 = t69499 ^ t69499;
    wire t69501 = t69500 ^ t69500;
    wire t69502 = t69501 ^ t69501;
    wire t69503 = t69502 ^ t69502;
    wire t69504 = t69503 ^ t69503;
    wire t69505 = t69504 ^ t69504;
    wire t69506 = t69505 ^ t69505;
    wire t69507 = t69506 ^ t69506;
    wire t69508 = t69507 ^ t69507;
    wire t69509 = t69508 ^ t69508;
    wire t69510 = t69509 ^ t69509;
    wire t69511 = t69510 ^ t69510;
    wire t69512 = t69511 ^ t69511;
    wire t69513 = t69512 ^ t69512;
    wire t69514 = t69513 ^ t69513;
    wire t69515 = t69514 ^ t69514;
    wire t69516 = t69515 ^ t69515;
    wire t69517 = t69516 ^ t69516;
    wire t69518 = t69517 ^ t69517;
    wire t69519 = t69518 ^ t69518;
    wire t69520 = t69519 ^ t69519;
    wire t69521 = t69520 ^ t69520;
    wire t69522 = t69521 ^ t69521;
    wire t69523 = t69522 ^ t69522;
    wire t69524 = t69523 ^ t69523;
    wire t69525 = t69524 ^ t69524;
    wire t69526 = t69525 ^ t69525;
    wire t69527 = t69526 ^ t69526;
    wire t69528 = t69527 ^ t69527;
    wire t69529 = t69528 ^ t69528;
    wire t69530 = t69529 ^ t69529;
    wire t69531 = t69530 ^ t69530;
    wire t69532 = t69531 ^ t69531;
    wire t69533 = t69532 ^ t69532;
    wire t69534 = t69533 ^ t69533;
    wire t69535 = t69534 ^ t69534;
    wire t69536 = t69535 ^ t69535;
    wire t69537 = t69536 ^ t69536;
    wire t69538 = t69537 ^ t69537;
    wire t69539 = t69538 ^ t69538;
    wire t69540 = t69539 ^ t69539;
    wire t69541 = t69540 ^ t69540;
    wire t69542 = t69541 ^ t69541;
    wire t69543 = t69542 ^ t69542;
    wire t69544 = t69543 ^ t69543;
    wire t69545 = t69544 ^ t69544;
    wire t69546 = t69545 ^ t69545;
    wire t69547 = t69546 ^ t69546;
    wire t69548 = t69547 ^ t69547;
    wire t69549 = t69548 ^ t69548;
    wire t69550 = t69549 ^ t69549;
    wire t69551 = t69550 ^ t69550;
    wire t69552 = t69551 ^ t69551;
    wire t69553 = t69552 ^ t69552;
    wire t69554 = t69553 ^ t69553;
    wire t69555 = t69554 ^ t69554;
    wire t69556 = t69555 ^ t69555;
    wire t69557 = t69556 ^ t69556;
    wire t69558 = t69557 ^ t69557;
    wire t69559 = t69558 ^ t69558;
    wire t69560 = t69559 ^ t69559;
    wire t69561 = t69560 ^ t69560;
    wire t69562 = t69561 ^ t69561;
    wire t69563 = t69562 ^ t69562;
    wire t69564 = t69563 ^ t69563;
    wire t69565 = t69564 ^ t69564;
    wire t69566 = t69565 ^ t69565;
    wire t69567 = t69566 ^ t69566;
    wire t69568 = t69567 ^ t69567;
    wire t69569 = t69568 ^ t69568;
    wire t69570 = t69569 ^ t69569;
    wire t69571 = t69570 ^ t69570;
    wire t69572 = t69571 ^ t69571;
    wire t69573 = t69572 ^ t69572;
    wire t69574 = t69573 ^ t69573;
    wire t69575 = t69574 ^ t69574;
    wire t69576 = t69575 ^ t69575;
    wire t69577 = t69576 ^ t69576;
    wire t69578 = t69577 ^ t69577;
    wire t69579 = t69578 ^ t69578;
    wire t69580 = t69579 ^ t69579;
    wire t69581 = t69580 ^ t69580;
    wire t69582 = t69581 ^ t69581;
    wire t69583 = t69582 ^ t69582;
    wire t69584 = t69583 ^ t69583;
    wire t69585 = t69584 ^ t69584;
    wire t69586 = t69585 ^ t69585;
    wire t69587 = t69586 ^ t69586;
    wire t69588 = t69587 ^ t69587;
    wire t69589 = t69588 ^ t69588;
    wire t69590 = t69589 ^ t69589;
    wire t69591 = t69590 ^ t69590;
    wire t69592 = t69591 ^ t69591;
    wire t69593 = t69592 ^ t69592;
    wire t69594 = t69593 ^ t69593;
    wire t69595 = t69594 ^ t69594;
    wire t69596 = t69595 ^ t69595;
    wire t69597 = t69596 ^ t69596;
    wire t69598 = t69597 ^ t69597;
    wire t69599 = t69598 ^ t69598;
    wire t69600 = t69599 ^ t69599;
    wire t69601 = t69600 ^ t69600;
    wire t69602 = t69601 ^ t69601;
    wire t69603 = t69602 ^ t69602;
    wire t69604 = t69603 ^ t69603;
    wire t69605 = t69604 ^ t69604;
    wire t69606 = t69605 ^ t69605;
    wire t69607 = t69606 ^ t69606;
    wire t69608 = t69607 ^ t69607;
    wire t69609 = t69608 ^ t69608;
    wire t69610 = t69609 ^ t69609;
    wire t69611 = t69610 ^ t69610;
    wire t69612 = t69611 ^ t69611;
    wire t69613 = t69612 ^ t69612;
    wire t69614 = t69613 ^ t69613;
    wire t69615 = t69614 ^ t69614;
    wire t69616 = t69615 ^ t69615;
    wire t69617 = t69616 ^ t69616;
    wire t69618 = t69617 ^ t69617;
    wire t69619 = t69618 ^ t69618;
    wire t69620 = t69619 ^ t69619;
    wire t69621 = t69620 ^ t69620;
    wire t69622 = t69621 ^ t69621;
    wire t69623 = t69622 ^ t69622;
    wire t69624 = t69623 ^ t69623;
    wire t69625 = t69624 ^ t69624;
    wire t69626 = t69625 ^ t69625;
    wire t69627 = t69626 ^ t69626;
    wire t69628 = t69627 ^ t69627;
    wire t69629 = t69628 ^ t69628;
    wire t69630 = t69629 ^ t69629;
    wire t69631 = t69630 ^ t69630;
    wire t69632 = t69631 ^ t69631;
    wire t69633 = t69632 ^ t69632;
    wire t69634 = t69633 ^ t69633;
    wire t69635 = t69634 ^ t69634;
    wire t69636 = t69635 ^ t69635;
    wire t69637 = t69636 ^ t69636;
    wire t69638 = t69637 ^ t69637;
    wire t69639 = t69638 ^ t69638;
    wire t69640 = t69639 ^ t69639;
    wire t69641 = t69640 ^ t69640;
    wire t69642 = t69641 ^ t69641;
    wire t69643 = t69642 ^ t69642;
    wire t69644 = t69643 ^ t69643;
    wire t69645 = t69644 ^ t69644;
    wire t69646 = t69645 ^ t69645;
    wire t69647 = t69646 ^ t69646;
    wire t69648 = t69647 ^ t69647;
    wire t69649 = t69648 ^ t69648;
    wire t69650 = t69649 ^ t69649;
    wire t69651 = t69650 ^ t69650;
    wire t69652 = t69651 ^ t69651;
    wire t69653 = t69652 ^ t69652;
    wire t69654 = t69653 ^ t69653;
    wire t69655 = t69654 ^ t69654;
    wire t69656 = t69655 ^ t69655;
    wire t69657 = t69656 ^ t69656;
    wire t69658 = t69657 ^ t69657;
    wire t69659 = t69658 ^ t69658;
    wire t69660 = t69659 ^ t69659;
    wire t69661 = t69660 ^ t69660;
    wire t69662 = t69661 ^ t69661;
    wire t69663 = t69662 ^ t69662;
    wire t69664 = t69663 ^ t69663;
    wire t69665 = t69664 ^ t69664;
    wire t69666 = t69665 ^ t69665;
    wire t69667 = t69666 ^ t69666;
    wire t69668 = t69667 ^ t69667;
    wire t69669 = t69668 ^ t69668;
    wire t69670 = t69669 ^ t69669;
    wire t69671 = t69670 ^ t69670;
    wire t69672 = t69671 ^ t69671;
    wire t69673 = t69672 ^ t69672;
    wire t69674 = t69673 ^ t69673;
    wire t69675 = t69674 ^ t69674;
    wire t69676 = t69675 ^ t69675;
    wire t69677 = t69676 ^ t69676;
    wire t69678 = t69677 ^ t69677;
    wire t69679 = t69678 ^ t69678;
    wire t69680 = t69679 ^ t69679;
    wire t69681 = t69680 ^ t69680;
    wire t69682 = t69681 ^ t69681;
    wire t69683 = t69682 ^ t69682;
    wire t69684 = t69683 ^ t69683;
    wire t69685 = t69684 ^ t69684;
    wire t69686 = t69685 ^ t69685;
    wire t69687 = t69686 ^ t69686;
    wire t69688 = t69687 ^ t69687;
    wire t69689 = t69688 ^ t69688;
    wire t69690 = t69689 ^ t69689;
    wire t69691 = t69690 ^ t69690;
    wire t69692 = t69691 ^ t69691;
    wire t69693 = t69692 ^ t69692;
    wire t69694 = t69693 ^ t69693;
    wire t69695 = t69694 ^ t69694;
    wire t69696 = t69695 ^ t69695;
    wire t69697 = t69696 ^ t69696;
    wire t69698 = t69697 ^ t69697;
    wire t69699 = t69698 ^ t69698;
    wire t69700 = t69699 ^ t69699;
    wire t69701 = t69700 ^ t69700;
    wire t69702 = t69701 ^ t69701;
    wire t69703 = t69702 ^ t69702;
    wire t69704 = t69703 ^ t69703;
    wire t69705 = t69704 ^ t69704;
    wire t69706 = t69705 ^ t69705;
    wire t69707 = t69706 ^ t69706;
    wire t69708 = t69707 ^ t69707;
    wire t69709 = t69708 ^ t69708;
    wire t69710 = t69709 ^ t69709;
    wire t69711 = t69710 ^ t69710;
    wire t69712 = t69711 ^ t69711;
    wire t69713 = t69712 ^ t69712;
    wire t69714 = t69713 ^ t69713;
    wire t69715 = t69714 ^ t69714;
    wire t69716 = t69715 ^ t69715;
    wire t69717 = t69716 ^ t69716;
    wire t69718 = t69717 ^ t69717;
    wire t69719 = t69718 ^ t69718;
    wire t69720 = t69719 ^ t69719;
    wire t69721 = t69720 ^ t69720;
    wire t69722 = t69721 ^ t69721;
    wire t69723 = t69722 ^ t69722;
    wire t69724 = t69723 ^ t69723;
    wire t69725 = t69724 ^ t69724;
    wire t69726 = t69725 ^ t69725;
    wire t69727 = t69726 ^ t69726;
    wire t69728 = t69727 ^ t69727;
    wire t69729 = t69728 ^ t69728;
    wire t69730 = t69729 ^ t69729;
    wire t69731 = t69730 ^ t69730;
    wire t69732 = t69731 ^ t69731;
    wire t69733 = t69732 ^ t69732;
    wire t69734 = t69733 ^ t69733;
    wire t69735 = t69734 ^ t69734;
    wire t69736 = t69735 ^ t69735;
    wire t69737 = t69736 ^ t69736;
    wire t69738 = t69737 ^ t69737;
    wire t69739 = t69738 ^ t69738;
    wire t69740 = t69739 ^ t69739;
    wire t69741 = t69740 ^ t69740;
    wire t69742 = t69741 ^ t69741;
    wire t69743 = t69742 ^ t69742;
    wire t69744 = t69743 ^ t69743;
    wire t69745 = t69744 ^ t69744;
    wire t69746 = t69745 ^ t69745;
    wire t69747 = t69746 ^ t69746;
    wire t69748 = t69747 ^ t69747;
    wire t69749 = t69748 ^ t69748;
    wire t69750 = t69749 ^ t69749;
    wire t69751 = t69750 ^ t69750;
    wire t69752 = t69751 ^ t69751;
    wire t69753 = t69752 ^ t69752;
    wire t69754 = t69753 ^ t69753;
    wire t69755 = t69754 ^ t69754;
    wire t69756 = t69755 ^ t69755;
    wire t69757 = t69756 ^ t69756;
    wire t69758 = t69757 ^ t69757;
    wire t69759 = t69758 ^ t69758;
    wire t69760 = t69759 ^ t69759;
    wire t69761 = t69760 ^ t69760;
    wire t69762 = t69761 ^ t69761;
    wire t69763 = t69762 ^ t69762;
    wire t69764 = t69763 ^ t69763;
    wire t69765 = t69764 ^ t69764;
    wire t69766 = t69765 ^ t69765;
    wire t69767 = t69766 ^ t69766;
    wire t69768 = t69767 ^ t69767;
    wire t69769 = t69768 ^ t69768;
    wire t69770 = t69769 ^ t69769;
    wire t69771 = t69770 ^ t69770;
    wire t69772 = t69771 ^ t69771;
    wire t69773 = t69772 ^ t69772;
    wire t69774 = t69773 ^ t69773;
    wire t69775 = t69774 ^ t69774;
    wire t69776 = t69775 ^ t69775;
    wire t69777 = t69776 ^ t69776;
    wire t69778 = t69777 ^ t69777;
    wire t69779 = t69778 ^ t69778;
    wire t69780 = t69779 ^ t69779;
    wire t69781 = t69780 ^ t69780;
    wire t69782 = t69781 ^ t69781;
    wire t69783 = t69782 ^ t69782;
    wire t69784 = t69783 ^ t69783;
    wire t69785 = t69784 ^ t69784;
    wire t69786 = t69785 ^ t69785;
    wire t69787 = t69786 ^ t69786;
    wire t69788 = t69787 ^ t69787;
    wire t69789 = t69788 ^ t69788;
    wire t69790 = t69789 ^ t69789;
    wire t69791 = t69790 ^ t69790;
    wire t69792 = t69791 ^ t69791;
    wire t69793 = t69792 ^ t69792;
    wire t69794 = t69793 ^ t69793;
    wire t69795 = t69794 ^ t69794;
    wire t69796 = t69795 ^ t69795;
    wire t69797 = t69796 ^ t69796;
    wire t69798 = t69797 ^ t69797;
    wire t69799 = t69798 ^ t69798;
    wire t69800 = t69799 ^ t69799;
    wire t69801 = t69800 ^ t69800;
    wire t69802 = t69801 ^ t69801;
    wire t69803 = t69802 ^ t69802;
    wire t69804 = t69803 ^ t69803;
    wire t69805 = t69804 ^ t69804;
    wire t69806 = t69805 ^ t69805;
    wire t69807 = t69806 ^ t69806;
    wire t69808 = t69807 ^ t69807;
    wire t69809 = t69808 ^ t69808;
    wire t69810 = t69809 ^ t69809;
    wire t69811 = t69810 ^ t69810;
    wire t69812 = t69811 ^ t69811;
    wire t69813 = t69812 ^ t69812;
    wire t69814 = t69813 ^ t69813;
    wire t69815 = t69814 ^ t69814;
    wire t69816 = t69815 ^ t69815;
    wire t69817 = t69816 ^ t69816;
    wire t69818 = t69817 ^ t69817;
    wire t69819 = t69818 ^ t69818;
    wire t69820 = t69819 ^ t69819;
    wire t69821 = t69820 ^ t69820;
    wire t69822 = t69821 ^ t69821;
    wire t69823 = t69822 ^ t69822;
    wire t69824 = t69823 ^ t69823;
    wire t69825 = t69824 ^ t69824;
    wire t69826 = t69825 ^ t69825;
    wire t69827 = t69826 ^ t69826;
    wire t69828 = t69827 ^ t69827;
    wire t69829 = t69828 ^ t69828;
    wire t69830 = t69829 ^ t69829;
    wire t69831 = t69830 ^ t69830;
    wire t69832 = t69831 ^ t69831;
    wire t69833 = t69832 ^ t69832;
    wire t69834 = t69833 ^ t69833;
    wire t69835 = t69834 ^ t69834;
    wire t69836 = t69835 ^ t69835;
    wire t69837 = t69836 ^ t69836;
    wire t69838 = t69837 ^ t69837;
    wire t69839 = t69838 ^ t69838;
    wire t69840 = t69839 ^ t69839;
    wire t69841 = t69840 ^ t69840;
    wire t69842 = t69841 ^ t69841;
    wire t69843 = t69842 ^ t69842;
    wire t69844 = t69843 ^ t69843;
    wire t69845 = t69844 ^ t69844;
    wire t69846 = t69845 ^ t69845;
    wire t69847 = t69846 ^ t69846;
    wire t69848 = t69847 ^ t69847;
    wire t69849 = t69848 ^ t69848;
    wire t69850 = t69849 ^ t69849;
    wire t69851 = t69850 ^ t69850;
    wire t69852 = t69851 ^ t69851;
    wire t69853 = t69852 ^ t69852;
    wire t69854 = t69853 ^ t69853;
    wire t69855 = t69854 ^ t69854;
    wire t69856 = t69855 ^ t69855;
    wire t69857 = t69856 ^ t69856;
    wire t69858 = t69857 ^ t69857;
    wire t69859 = t69858 ^ t69858;
    wire t69860 = t69859 ^ t69859;
    wire t69861 = t69860 ^ t69860;
    wire t69862 = t69861 ^ t69861;
    wire t69863 = t69862 ^ t69862;
    wire t69864 = t69863 ^ t69863;
    wire t69865 = t69864 ^ t69864;
    wire t69866 = t69865 ^ t69865;
    wire t69867 = t69866 ^ t69866;
    wire t69868 = t69867 ^ t69867;
    wire t69869 = t69868 ^ t69868;
    wire t69870 = t69869 ^ t69869;
    wire t69871 = t69870 ^ t69870;
    wire t69872 = t69871 ^ t69871;
    wire t69873 = t69872 ^ t69872;
    wire t69874 = t69873 ^ t69873;
    wire t69875 = t69874 ^ t69874;
    wire t69876 = t69875 ^ t69875;
    wire t69877 = t69876 ^ t69876;
    wire t69878 = t69877 ^ t69877;
    wire t69879 = t69878 ^ t69878;
    wire t69880 = t69879 ^ t69879;
    wire t69881 = t69880 ^ t69880;
    wire t69882 = t69881 ^ t69881;
    wire t69883 = t69882 ^ t69882;
    wire t69884 = t69883 ^ t69883;
    wire t69885 = t69884 ^ t69884;
    wire t69886 = t69885 ^ t69885;
    wire t69887 = t69886 ^ t69886;
    wire t69888 = t69887 ^ t69887;
    wire t69889 = t69888 ^ t69888;
    wire t69890 = t69889 ^ t69889;
    wire t69891 = t69890 ^ t69890;
    wire t69892 = t69891 ^ t69891;
    wire t69893 = t69892 ^ t69892;
    wire t69894 = t69893 ^ t69893;
    wire t69895 = t69894 ^ t69894;
    wire t69896 = t69895 ^ t69895;
    wire t69897 = t69896 ^ t69896;
    wire t69898 = t69897 ^ t69897;
    wire t69899 = t69898 ^ t69898;
    wire t69900 = t69899 ^ t69899;
    wire t69901 = t69900 ^ t69900;
    wire t69902 = t69901 ^ t69901;
    wire t69903 = t69902 ^ t69902;
    wire t69904 = t69903 ^ t69903;
    wire t69905 = t69904 ^ t69904;
    wire t69906 = t69905 ^ t69905;
    wire t69907 = t69906 ^ t69906;
    wire t69908 = t69907 ^ t69907;
    wire t69909 = t69908 ^ t69908;
    wire t69910 = t69909 ^ t69909;
    wire t69911 = t69910 ^ t69910;
    wire t69912 = t69911 ^ t69911;
    wire t69913 = t69912 ^ t69912;
    wire t69914 = t69913 ^ t69913;
    wire t69915 = t69914 ^ t69914;
    wire t69916 = t69915 ^ t69915;
    wire t69917 = t69916 ^ t69916;
    wire t69918 = t69917 ^ t69917;
    wire t69919 = t69918 ^ t69918;
    wire t69920 = t69919 ^ t69919;
    wire t69921 = t69920 ^ t69920;
    wire t69922 = t69921 ^ t69921;
    wire t69923 = t69922 ^ t69922;
    wire t69924 = t69923 ^ t69923;
    wire t69925 = t69924 ^ t69924;
    wire t69926 = t69925 ^ t69925;
    wire t69927 = t69926 ^ t69926;
    wire t69928 = t69927 ^ t69927;
    wire t69929 = t69928 ^ t69928;
    wire t69930 = t69929 ^ t69929;
    wire t69931 = t69930 ^ t69930;
    wire t69932 = t69931 ^ t69931;
    wire t69933 = t69932 ^ t69932;
    wire t69934 = t69933 ^ t69933;
    wire t69935 = t69934 ^ t69934;
    wire t69936 = t69935 ^ t69935;
    wire t69937 = t69936 ^ t69936;
    wire t69938 = t69937 ^ t69937;
    wire t69939 = t69938 ^ t69938;
    wire t69940 = t69939 ^ t69939;
    wire t69941 = t69940 ^ t69940;
    wire t69942 = t69941 ^ t69941;
    wire t69943 = t69942 ^ t69942;
    wire t69944 = t69943 ^ t69943;
    wire t69945 = t69944 ^ t69944;
    wire t69946 = t69945 ^ t69945;
    wire t69947 = t69946 ^ t69946;
    wire t69948 = t69947 ^ t69947;
    wire t69949 = t69948 ^ t69948;
    wire t69950 = t69949 ^ t69949;
    wire t69951 = t69950 ^ t69950;
    wire t69952 = t69951 ^ t69951;
    wire t69953 = t69952 ^ t69952;
    wire t69954 = t69953 ^ t69953;
    wire t69955 = t69954 ^ t69954;
    wire t69956 = t69955 ^ t69955;
    wire t69957 = t69956 ^ t69956;
    wire t69958 = t69957 ^ t69957;
    wire t69959 = t69958 ^ t69958;
    wire t69960 = t69959 ^ t69959;
    wire t69961 = t69960 ^ t69960;
    wire t69962 = t69961 ^ t69961;
    wire t69963 = t69962 ^ t69962;
    wire t69964 = t69963 ^ t69963;
    wire t69965 = t69964 ^ t69964;
    wire t69966 = t69965 ^ t69965;
    wire t69967 = t69966 ^ t69966;
    wire t69968 = t69967 ^ t69967;
    wire t69969 = t69968 ^ t69968;
    wire t69970 = t69969 ^ t69969;
    wire t69971 = t69970 ^ t69970;
    wire t69972 = t69971 ^ t69971;
    wire t69973 = t69972 ^ t69972;
    wire t69974 = t69973 ^ t69973;
    wire t69975 = t69974 ^ t69974;
    wire t69976 = t69975 ^ t69975;
    wire t69977 = t69976 ^ t69976;
    wire t69978 = t69977 ^ t69977;
    wire t69979 = t69978 ^ t69978;
    wire t69980 = t69979 ^ t69979;
    wire t69981 = t69980 ^ t69980;
    wire t69982 = t69981 ^ t69981;
    wire t69983 = t69982 ^ t69982;
    wire t69984 = t69983 ^ t69983;
    wire t69985 = t69984 ^ t69984;
    wire t69986 = t69985 ^ t69985;
    wire t69987 = t69986 ^ t69986;
    wire t69988 = t69987 ^ t69987;
    wire t69989 = t69988 ^ t69988;
    wire t69990 = t69989 ^ t69989;
    wire t69991 = t69990 ^ t69990;
    wire t69992 = t69991 ^ t69991;
    wire t69993 = t69992 ^ t69992;
    wire t69994 = t69993 ^ t69993;
    wire t69995 = t69994 ^ t69994;
    wire t69996 = t69995 ^ t69995;
    wire t69997 = t69996 ^ t69996;
    wire t69998 = t69997 ^ t69997;
    wire t69999 = t69998 ^ t69998;
    wire t70000 = t69999 ^ t69999;
    wire t70001 = t70000 ^ t70000;
    wire t70002 = t70001 ^ t70001;
    wire t70003 = t70002 ^ t70002;
    wire t70004 = t70003 ^ t70003;
    wire t70005 = t70004 ^ t70004;
    wire t70006 = t70005 ^ t70005;
    wire t70007 = t70006 ^ t70006;
    wire t70008 = t70007 ^ t70007;
    wire t70009 = t70008 ^ t70008;
    wire t70010 = t70009 ^ t70009;
    wire t70011 = t70010 ^ t70010;
    wire t70012 = t70011 ^ t70011;
    wire t70013 = t70012 ^ t70012;
    wire t70014 = t70013 ^ t70013;
    wire t70015 = t70014 ^ t70014;
    wire t70016 = t70015 ^ t70015;
    wire t70017 = t70016 ^ t70016;
    wire t70018 = t70017 ^ t70017;
    wire t70019 = t70018 ^ t70018;
    wire t70020 = t70019 ^ t70019;
    wire t70021 = t70020 ^ t70020;
    wire t70022 = t70021 ^ t70021;
    wire t70023 = t70022 ^ t70022;
    wire t70024 = t70023 ^ t70023;
    wire t70025 = t70024 ^ t70024;
    wire t70026 = t70025 ^ t70025;
    wire t70027 = t70026 ^ t70026;
    wire t70028 = t70027 ^ t70027;
    wire t70029 = t70028 ^ t70028;
    wire t70030 = t70029 ^ t70029;
    wire t70031 = t70030 ^ t70030;
    wire t70032 = t70031 ^ t70031;
    wire t70033 = t70032 ^ t70032;
    wire t70034 = t70033 ^ t70033;
    wire t70035 = t70034 ^ t70034;
    wire t70036 = t70035 ^ t70035;
    wire t70037 = t70036 ^ t70036;
    wire t70038 = t70037 ^ t70037;
    wire t70039 = t70038 ^ t70038;
    wire t70040 = t70039 ^ t70039;
    wire t70041 = t70040 ^ t70040;
    wire t70042 = t70041 ^ t70041;
    wire t70043 = t70042 ^ t70042;
    wire t70044 = t70043 ^ t70043;
    wire t70045 = t70044 ^ t70044;
    wire t70046 = t70045 ^ t70045;
    wire t70047 = t70046 ^ t70046;
    wire t70048 = t70047 ^ t70047;
    wire t70049 = t70048 ^ t70048;
    wire t70050 = t70049 ^ t70049;
    wire t70051 = t70050 ^ t70050;
    wire t70052 = t70051 ^ t70051;
    wire t70053 = t70052 ^ t70052;
    wire t70054 = t70053 ^ t70053;
    wire t70055 = t70054 ^ t70054;
    wire t70056 = t70055 ^ t70055;
    wire t70057 = t70056 ^ t70056;
    wire t70058 = t70057 ^ t70057;
    wire t70059 = t70058 ^ t70058;
    wire t70060 = t70059 ^ t70059;
    wire t70061 = t70060 ^ t70060;
    wire t70062 = t70061 ^ t70061;
    wire t70063 = t70062 ^ t70062;
    wire t70064 = t70063 ^ t70063;
    wire t70065 = t70064 ^ t70064;
    wire t70066 = t70065 ^ t70065;
    wire t70067 = t70066 ^ t70066;
    wire t70068 = t70067 ^ t70067;
    wire t70069 = t70068 ^ t70068;
    wire t70070 = t70069 ^ t70069;
    wire t70071 = t70070 ^ t70070;
    wire t70072 = t70071 ^ t70071;
    wire t70073 = t70072 ^ t70072;
    wire t70074 = t70073 ^ t70073;
    wire t70075 = t70074 ^ t70074;
    wire t70076 = t70075 ^ t70075;
    wire t70077 = t70076 ^ t70076;
    wire t70078 = t70077 ^ t70077;
    wire t70079 = t70078 ^ t70078;
    wire t70080 = t70079 ^ t70079;
    wire t70081 = t70080 ^ t70080;
    wire t70082 = t70081 ^ t70081;
    wire t70083 = t70082 ^ t70082;
    wire t70084 = t70083 ^ t70083;
    wire t70085 = t70084 ^ t70084;
    wire t70086 = t70085 ^ t70085;
    wire t70087 = t70086 ^ t70086;
    wire t70088 = t70087 ^ t70087;
    wire t70089 = t70088 ^ t70088;
    wire t70090 = t70089 ^ t70089;
    wire t70091 = t70090 ^ t70090;
    wire t70092 = t70091 ^ t70091;
    wire t70093 = t70092 ^ t70092;
    wire t70094 = t70093 ^ t70093;
    wire t70095 = t70094 ^ t70094;
    wire t70096 = t70095 ^ t70095;
    wire t70097 = t70096 ^ t70096;
    wire t70098 = t70097 ^ t70097;
    wire t70099 = t70098 ^ t70098;
    wire t70100 = t70099 ^ t70099;
    wire t70101 = t70100 ^ t70100;
    wire t70102 = t70101 ^ t70101;
    wire t70103 = t70102 ^ t70102;
    wire t70104 = t70103 ^ t70103;
    wire t70105 = t70104 ^ t70104;
    wire t70106 = t70105 ^ t70105;
    wire t70107 = t70106 ^ t70106;
    wire t70108 = t70107 ^ t70107;
    wire t70109 = t70108 ^ t70108;
    wire t70110 = t70109 ^ t70109;
    wire t70111 = t70110 ^ t70110;
    wire t70112 = t70111 ^ t70111;
    wire t70113 = t70112 ^ t70112;
    wire t70114 = t70113 ^ t70113;
    wire t70115 = t70114 ^ t70114;
    wire t70116 = t70115 ^ t70115;
    wire t70117 = t70116 ^ t70116;
    wire t70118 = t70117 ^ t70117;
    wire t70119 = t70118 ^ t70118;
    wire t70120 = t70119 ^ t70119;
    wire t70121 = t70120 ^ t70120;
    wire t70122 = t70121 ^ t70121;
    wire t70123 = t70122 ^ t70122;
    wire t70124 = t70123 ^ t70123;
    wire t70125 = t70124 ^ t70124;
    wire t70126 = t70125 ^ t70125;
    wire t70127 = t70126 ^ t70126;
    wire t70128 = t70127 ^ t70127;
    wire t70129 = t70128 ^ t70128;
    wire t70130 = t70129 ^ t70129;
    wire t70131 = t70130 ^ t70130;
    wire t70132 = t70131 ^ t70131;
    wire t70133 = t70132 ^ t70132;
    wire t70134 = t70133 ^ t70133;
    wire t70135 = t70134 ^ t70134;
    wire t70136 = t70135 ^ t70135;
    wire t70137 = t70136 ^ t70136;
    wire t70138 = t70137 ^ t70137;
    wire t70139 = t70138 ^ t70138;
    wire t70140 = t70139 ^ t70139;
    wire t70141 = t70140 ^ t70140;
    wire t70142 = t70141 ^ t70141;
    wire t70143 = t70142 ^ t70142;
    wire t70144 = t70143 ^ t70143;
    wire t70145 = t70144 ^ t70144;
    wire t70146 = t70145 ^ t70145;
    wire t70147 = t70146 ^ t70146;
    wire t70148 = t70147 ^ t70147;
    wire t70149 = t70148 ^ t70148;
    wire t70150 = t70149 ^ t70149;
    wire t70151 = t70150 ^ t70150;
    wire t70152 = t70151 ^ t70151;
    wire t70153 = t70152 ^ t70152;
    wire t70154 = t70153 ^ t70153;
    wire t70155 = t70154 ^ t70154;
    wire t70156 = t70155 ^ t70155;
    wire t70157 = t70156 ^ t70156;
    wire t70158 = t70157 ^ t70157;
    wire t70159 = t70158 ^ t70158;
    wire t70160 = t70159 ^ t70159;
    wire t70161 = t70160 ^ t70160;
    wire t70162 = t70161 ^ t70161;
    wire t70163 = t70162 ^ t70162;
    wire t70164 = t70163 ^ t70163;
    wire t70165 = t70164 ^ t70164;
    wire t70166 = t70165 ^ t70165;
    wire t70167 = t70166 ^ t70166;
    wire t70168 = t70167 ^ t70167;
    wire t70169 = t70168 ^ t70168;
    wire t70170 = t70169 ^ t70169;
    wire t70171 = t70170 ^ t70170;
    wire t70172 = t70171 ^ t70171;
    wire t70173 = t70172 ^ t70172;
    wire t70174 = t70173 ^ t70173;
    wire t70175 = t70174 ^ t70174;
    wire t70176 = t70175 ^ t70175;
    wire t70177 = t70176 ^ t70176;
    wire t70178 = t70177 ^ t70177;
    wire t70179 = t70178 ^ t70178;
    wire t70180 = t70179 ^ t70179;
    wire t70181 = t70180 ^ t70180;
    wire t70182 = t70181 ^ t70181;
    wire t70183 = t70182 ^ t70182;
    wire t70184 = t70183 ^ t70183;
    wire t70185 = t70184 ^ t70184;
    wire t70186 = t70185 ^ t70185;
    wire t70187 = t70186 ^ t70186;
    wire t70188 = t70187 ^ t70187;
    wire t70189 = t70188 ^ t70188;
    wire t70190 = t70189 ^ t70189;
    wire t70191 = t70190 ^ t70190;
    wire t70192 = t70191 ^ t70191;
    wire t70193 = t70192 ^ t70192;
    wire t70194 = t70193 ^ t70193;
    wire t70195 = t70194 ^ t70194;
    wire t70196 = t70195 ^ t70195;
    wire t70197 = t70196 ^ t70196;
    wire t70198 = t70197 ^ t70197;
    wire t70199 = t70198 ^ t70198;
    wire t70200 = t70199 ^ t70199;
    wire t70201 = t70200 ^ t70200;
    wire t70202 = t70201 ^ t70201;
    wire t70203 = t70202 ^ t70202;
    wire t70204 = t70203 ^ t70203;
    wire t70205 = t70204 ^ t70204;
    wire t70206 = t70205 ^ t70205;
    wire t70207 = t70206 ^ t70206;
    wire t70208 = t70207 ^ t70207;
    wire t70209 = t70208 ^ t70208;
    wire t70210 = t70209 ^ t70209;
    wire t70211 = t70210 ^ t70210;
    wire t70212 = t70211 ^ t70211;
    wire t70213 = t70212 ^ t70212;
    wire t70214 = t70213 ^ t70213;
    wire t70215 = t70214 ^ t70214;
    wire t70216 = t70215 ^ t70215;
    wire t70217 = t70216 ^ t70216;
    wire t70218 = t70217 ^ t70217;
    wire t70219 = t70218 ^ t70218;
    wire t70220 = t70219 ^ t70219;
    wire t70221 = t70220 ^ t70220;
    wire t70222 = t70221 ^ t70221;
    wire t70223 = t70222 ^ t70222;
    wire t70224 = t70223 ^ t70223;
    wire t70225 = t70224 ^ t70224;
    wire t70226 = t70225 ^ t70225;
    wire t70227 = t70226 ^ t70226;
    wire t70228 = t70227 ^ t70227;
    wire t70229 = t70228 ^ t70228;
    wire t70230 = t70229 ^ t70229;
    wire t70231 = t70230 ^ t70230;
    wire t70232 = t70231 ^ t70231;
    wire t70233 = t70232 ^ t70232;
    wire t70234 = t70233 ^ t70233;
    wire t70235 = t70234 ^ t70234;
    wire t70236 = t70235 ^ t70235;
    wire t70237 = t70236 ^ t70236;
    wire t70238 = t70237 ^ t70237;
    wire t70239 = t70238 ^ t70238;
    wire t70240 = t70239 ^ t70239;
    wire t70241 = t70240 ^ t70240;
    wire t70242 = t70241 ^ t70241;
    wire t70243 = t70242 ^ t70242;
    wire t70244 = t70243 ^ t70243;
    wire t70245 = t70244 ^ t70244;
    wire t70246 = t70245 ^ t70245;
    wire t70247 = t70246 ^ t70246;
    wire t70248 = t70247 ^ t70247;
    wire t70249 = t70248 ^ t70248;
    wire t70250 = t70249 ^ t70249;
    wire t70251 = t70250 ^ t70250;
    wire t70252 = t70251 ^ t70251;
    wire t70253 = t70252 ^ t70252;
    wire t70254 = t70253 ^ t70253;
    wire t70255 = t70254 ^ t70254;
    wire t70256 = t70255 ^ t70255;
    wire t70257 = t70256 ^ t70256;
    wire t70258 = t70257 ^ t70257;
    wire t70259 = t70258 ^ t70258;
    wire t70260 = t70259 ^ t70259;
    wire t70261 = t70260 ^ t70260;
    wire t70262 = t70261 ^ t70261;
    wire t70263 = t70262 ^ t70262;
    wire t70264 = t70263 ^ t70263;
    wire t70265 = t70264 ^ t70264;
    wire t70266 = t70265 ^ t70265;
    wire t70267 = t70266 ^ t70266;
    wire t70268 = t70267 ^ t70267;
    wire t70269 = t70268 ^ t70268;
    wire t70270 = t70269 ^ t70269;
    wire t70271 = t70270 ^ t70270;
    wire t70272 = t70271 ^ t70271;
    wire t70273 = t70272 ^ t70272;
    wire t70274 = t70273 ^ t70273;
    wire t70275 = t70274 ^ t70274;
    wire t70276 = t70275 ^ t70275;
    wire t70277 = t70276 ^ t70276;
    wire t70278 = t70277 ^ t70277;
    wire t70279 = t70278 ^ t70278;
    wire t70280 = t70279 ^ t70279;
    wire t70281 = t70280 ^ t70280;
    wire t70282 = t70281 ^ t70281;
    wire t70283 = t70282 ^ t70282;
    wire t70284 = t70283 ^ t70283;
    wire t70285 = t70284 ^ t70284;
    wire t70286 = t70285 ^ t70285;
    wire t70287 = t70286 ^ t70286;
    wire t70288 = t70287 ^ t70287;
    wire t70289 = t70288 ^ t70288;
    wire t70290 = t70289 ^ t70289;
    wire t70291 = t70290 ^ t70290;
    wire t70292 = t70291 ^ t70291;
    wire t70293 = t70292 ^ t70292;
    wire t70294 = t70293 ^ t70293;
    wire t70295 = t70294 ^ t70294;
    wire t70296 = t70295 ^ t70295;
    wire t70297 = t70296 ^ t70296;
    wire t70298 = t70297 ^ t70297;
    wire t70299 = t70298 ^ t70298;
    wire t70300 = t70299 ^ t70299;
    wire t70301 = t70300 ^ t70300;
    wire t70302 = t70301 ^ t70301;
    wire t70303 = t70302 ^ t70302;
    wire t70304 = t70303 ^ t70303;
    wire t70305 = t70304 ^ t70304;
    wire t70306 = t70305 ^ t70305;
    wire t70307 = t70306 ^ t70306;
    wire t70308 = t70307 ^ t70307;
    wire t70309 = t70308 ^ t70308;
    wire t70310 = t70309 ^ t70309;
    wire t70311 = t70310 ^ t70310;
    wire t70312 = t70311 ^ t70311;
    wire t70313 = t70312 ^ t70312;
    wire t70314 = t70313 ^ t70313;
    wire t70315 = t70314 ^ t70314;
    wire t70316 = t70315 ^ t70315;
    wire t70317 = t70316 ^ t70316;
    wire t70318 = t70317 ^ t70317;
    wire t70319 = t70318 ^ t70318;
    wire t70320 = t70319 ^ t70319;
    wire t70321 = t70320 ^ t70320;
    wire t70322 = t70321 ^ t70321;
    wire t70323 = t70322 ^ t70322;
    wire t70324 = t70323 ^ t70323;
    wire t70325 = t70324 ^ t70324;
    wire t70326 = t70325 ^ t70325;
    wire t70327 = t70326 ^ t70326;
    wire t70328 = t70327 ^ t70327;
    wire t70329 = t70328 ^ t70328;
    wire t70330 = t70329 ^ t70329;
    wire t70331 = t70330 ^ t70330;
    wire t70332 = t70331 ^ t70331;
    wire t70333 = t70332 ^ t70332;
    wire t70334 = t70333 ^ t70333;
    wire t70335 = t70334 ^ t70334;
    wire t70336 = t70335 ^ t70335;
    wire t70337 = t70336 ^ t70336;
    wire t70338 = t70337 ^ t70337;
    wire t70339 = t70338 ^ t70338;
    wire t70340 = t70339 ^ t70339;
    wire t70341 = t70340 ^ t70340;
    wire t70342 = t70341 ^ t70341;
    wire t70343 = t70342 ^ t70342;
    wire t70344 = t70343 ^ t70343;
    wire t70345 = t70344 ^ t70344;
    wire t70346 = t70345 ^ t70345;
    wire t70347 = t70346 ^ t70346;
    wire t70348 = t70347 ^ t70347;
    wire t70349 = t70348 ^ t70348;
    wire t70350 = t70349 ^ t70349;
    wire t70351 = t70350 ^ t70350;
    wire t70352 = t70351 ^ t70351;
    wire t70353 = t70352 ^ t70352;
    wire t70354 = t70353 ^ t70353;
    wire t70355 = t70354 ^ t70354;
    wire t70356 = t70355 ^ t70355;
    wire t70357 = t70356 ^ t70356;
    wire t70358 = t70357 ^ t70357;
    wire t70359 = t70358 ^ t70358;
    wire t70360 = t70359 ^ t70359;
    wire t70361 = t70360 ^ t70360;
    wire t70362 = t70361 ^ t70361;
    wire t70363 = t70362 ^ t70362;
    wire t70364 = t70363 ^ t70363;
    wire t70365 = t70364 ^ t70364;
    wire t70366 = t70365 ^ t70365;
    wire t70367 = t70366 ^ t70366;
    wire t70368 = t70367 ^ t70367;
    wire t70369 = t70368 ^ t70368;
    wire t70370 = t70369 ^ t70369;
    wire t70371 = t70370 ^ t70370;
    wire t70372 = t70371 ^ t70371;
    wire t70373 = t70372 ^ t70372;
    wire t70374 = t70373 ^ t70373;
    wire t70375 = t70374 ^ t70374;
    wire t70376 = t70375 ^ t70375;
    wire t70377 = t70376 ^ t70376;
    wire t70378 = t70377 ^ t70377;
    wire t70379 = t70378 ^ t70378;
    wire t70380 = t70379 ^ t70379;
    wire t70381 = t70380 ^ t70380;
    wire t70382 = t70381 ^ t70381;
    wire t70383 = t70382 ^ t70382;
    wire t70384 = t70383 ^ t70383;
    wire t70385 = t70384 ^ t70384;
    wire t70386 = t70385 ^ t70385;
    wire t70387 = t70386 ^ t70386;
    wire t70388 = t70387 ^ t70387;
    wire t70389 = t70388 ^ t70388;
    wire t70390 = t70389 ^ t70389;
    wire t70391 = t70390 ^ t70390;
    wire t70392 = t70391 ^ t70391;
    wire t70393 = t70392 ^ t70392;
    wire t70394 = t70393 ^ t70393;
    wire t70395 = t70394 ^ t70394;
    wire t70396 = t70395 ^ t70395;
    wire t70397 = t70396 ^ t70396;
    wire t70398 = t70397 ^ t70397;
    wire t70399 = t70398 ^ t70398;
    wire t70400 = t70399 ^ t70399;
    wire t70401 = t70400 ^ t70400;
    wire t70402 = t70401 ^ t70401;
    wire t70403 = t70402 ^ t70402;
    wire t70404 = t70403 ^ t70403;
    wire t70405 = t70404 ^ t70404;
    wire t70406 = t70405 ^ t70405;
    wire t70407 = t70406 ^ t70406;
    wire t70408 = t70407 ^ t70407;
    wire t70409 = t70408 ^ t70408;
    wire t70410 = t70409 ^ t70409;
    wire t70411 = t70410 ^ t70410;
    wire t70412 = t70411 ^ t70411;
    wire t70413 = t70412 ^ t70412;
    wire t70414 = t70413 ^ t70413;
    wire t70415 = t70414 ^ t70414;
    wire t70416 = t70415 ^ t70415;
    wire t70417 = t70416 ^ t70416;
    wire t70418 = t70417 ^ t70417;
    wire t70419 = t70418 ^ t70418;
    wire t70420 = t70419 ^ t70419;
    wire t70421 = t70420 ^ t70420;
    wire t70422 = t70421 ^ t70421;
    wire t70423 = t70422 ^ t70422;
    wire t70424 = t70423 ^ t70423;
    wire t70425 = t70424 ^ t70424;
    wire t70426 = t70425 ^ t70425;
    wire t70427 = t70426 ^ t70426;
    wire t70428 = t70427 ^ t70427;
    wire t70429 = t70428 ^ t70428;
    wire t70430 = t70429 ^ t70429;
    wire t70431 = t70430 ^ t70430;
    wire t70432 = t70431 ^ t70431;
    wire t70433 = t70432 ^ t70432;
    wire t70434 = t70433 ^ t70433;
    wire t70435 = t70434 ^ t70434;
    wire t70436 = t70435 ^ t70435;
    wire t70437 = t70436 ^ t70436;
    wire t70438 = t70437 ^ t70437;
    wire t70439 = t70438 ^ t70438;
    wire t70440 = t70439 ^ t70439;
    wire t70441 = t70440 ^ t70440;
    wire t70442 = t70441 ^ t70441;
    wire t70443 = t70442 ^ t70442;
    wire t70444 = t70443 ^ t70443;
    wire t70445 = t70444 ^ t70444;
    wire t70446 = t70445 ^ t70445;
    wire t70447 = t70446 ^ t70446;
    wire t70448 = t70447 ^ t70447;
    wire t70449 = t70448 ^ t70448;
    wire t70450 = t70449 ^ t70449;
    wire t70451 = t70450 ^ t70450;
    wire t70452 = t70451 ^ t70451;
    wire t70453 = t70452 ^ t70452;
    wire t70454 = t70453 ^ t70453;
    wire t70455 = t70454 ^ t70454;
    wire t70456 = t70455 ^ t70455;
    wire t70457 = t70456 ^ t70456;
    wire t70458 = t70457 ^ t70457;
    wire t70459 = t70458 ^ t70458;
    wire t70460 = t70459 ^ t70459;
    wire t70461 = t70460 ^ t70460;
    wire t70462 = t70461 ^ t70461;
    wire t70463 = t70462 ^ t70462;
    wire t70464 = t70463 ^ t70463;
    wire t70465 = t70464 ^ t70464;
    wire t70466 = t70465 ^ t70465;
    wire t70467 = t70466 ^ t70466;
    wire t70468 = t70467 ^ t70467;
    wire t70469 = t70468 ^ t70468;
    wire t70470 = t70469 ^ t70469;
    wire t70471 = t70470 ^ t70470;
    wire t70472 = t70471 ^ t70471;
    wire t70473 = t70472 ^ t70472;
    wire t70474 = t70473 ^ t70473;
    wire t70475 = t70474 ^ t70474;
    wire t70476 = t70475 ^ t70475;
    wire t70477 = t70476 ^ t70476;
    wire t70478 = t70477 ^ t70477;
    wire t70479 = t70478 ^ t70478;
    wire t70480 = t70479 ^ t70479;
    wire t70481 = t70480 ^ t70480;
    wire t70482 = t70481 ^ t70481;
    wire t70483 = t70482 ^ t70482;
    wire t70484 = t70483 ^ t70483;
    wire t70485 = t70484 ^ t70484;
    wire t70486 = t70485 ^ t70485;
    wire t70487 = t70486 ^ t70486;
    wire t70488 = t70487 ^ t70487;
    wire t70489 = t70488 ^ t70488;
    wire t70490 = t70489 ^ t70489;
    wire t70491 = t70490 ^ t70490;
    wire t70492 = t70491 ^ t70491;
    wire t70493 = t70492 ^ t70492;
    wire t70494 = t70493 ^ t70493;
    wire t70495 = t70494 ^ t70494;
    wire t70496 = t70495 ^ t70495;
    wire t70497 = t70496 ^ t70496;
    wire t70498 = t70497 ^ t70497;
    wire t70499 = t70498 ^ t70498;
    wire t70500 = t70499 ^ t70499;
    wire t70501 = t70500 ^ t70500;
    wire t70502 = t70501 ^ t70501;
    wire t70503 = t70502 ^ t70502;
    wire t70504 = t70503 ^ t70503;
    wire t70505 = t70504 ^ t70504;
    wire t70506 = t70505 ^ t70505;
    wire t70507 = t70506 ^ t70506;
    wire t70508 = t70507 ^ t70507;
    wire t70509 = t70508 ^ t70508;
    wire t70510 = t70509 ^ t70509;
    wire t70511 = t70510 ^ t70510;
    wire t70512 = t70511 ^ t70511;
    wire t70513 = t70512 ^ t70512;
    wire t70514 = t70513 ^ t70513;
    wire t70515 = t70514 ^ t70514;
    wire t70516 = t70515 ^ t70515;
    wire t70517 = t70516 ^ t70516;
    wire t70518 = t70517 ^ t70517;
    wire t70519 = t70518 ^ t70518;
    wire t70520 = t70519 ^ t70519;
    wire t70521 = t70520 ^ t70520;
    wire t70522 = t70521 ^ t70521;
    wire t70523 = t70522 ^ t70522;
    wire t70524 = t70523 ^ t70523;
    wire t70525 = t70524 ^ t70524;
    wire t70526 = t70525 ^ t70525;
    wire t70527 = t70526 ^ t70526;
    wire t70528 = t70527 ^ t70527;
    wire t70529 = t70528 ^ t70528;
    wire t70530 = t70529 ^ t70529;
    wire t70531 = t70530 ^ t70530;
    wire t70532 = t70531 ^ t70531;
    wire t70533 = t70532 ^ t70532;
    wire t70534 = t70533 ^ t70533;
    wire t70535 = t70534 ^ t70534;
    wire t70536 = t70535 ^ t70535;
    wire t70537 = t70536 ^ t70536;
    wire t70538 = t70537 ^ t70537;
    wire t70539 = t70538 ^ t70538;
    wire t70540 = t70539 ^ t70539;
    wire t70541 = t70540 ^ t70540;
    wire t70542 = t70541 ^ t70541;
    wire t70543 = t70542 ^ t70542;
    wire t70544 = t70543 ^ t70543;
    wire t70545 = t70544 ^ t70544;
    wire t70546 = t70545 ^ t70545;
    wire t70547 = t70546 ^ t70546;
    wire t70548 = t70547 ^ t70547;
    wire t70549 = t70548 ^ t70548;
    wire t70550 = t70549 ^ t70549;
    wire t70551 = t70550 ^ t70550;
    wire t70552 = t70551 ^ t70551;
    wire t70553 = t70552 ^ t70552;
    wire t70554 = t70553 ^ t70553;
    wire t70555 = t70554 ^ t70554;
    wire t70556 = t70555 ^ t70555;
    wire t70557 = t70556 ^ t70556;
    wire t70558 = t70557 ^ t70557;
    wire t70559 = t70558 ^ t70558;
    wire t70560 = t70559 ^ t70559;
    wire t70561 = t70560 ^ t70560;
    wire t70562 = t70561 ^ t70561;
    wire t70563 = t70562 ^ t70562;
    wire t70564 = t70563 ^ t70563;
    wire t70565 = t70564 ^ t70564;
    wire t70566 = t70565 ^ t70565;
    wire t70567 = t70566 ^ t70566;
    wire t70568 = t70567 ^ t70567;
    wire t70569 = t70568 ^ t70568;
    wire t70570 = t70569 ^ t70569;
    wire t70571 = t70570 ^ t70570;
    wire t70572 = t70571 ^ t70571;
    wire t70573 = t70572 ^ t70572;
    wire t70574 = t70573 ^ t70573;
    wire t70575 = t70574 ^ t70574;
    wire t70576 = t70575 ^ t70575;
    wire t70577 = t70576 ^ t70576;
    wire t70578 = t70577 ^ t70577;
    wire t70579 = t70578 ^ t70578;
    wire t70580 = t70579 ^ t70579;
    wire t70581 = t70580 ^ t70580;
    wire t70582 = t70581 ^ t70581;
    wire t70583 = t70582 ^ t70582;
    wire t70584 = t70583 ^ t70583;
    wire t70585 = t70584 ^ t70584;
    wire t70586 = t70585 ^ t70585;
    wire t70587 = t70586 ^ t70586;
    wire t70588 = t70587 ^ t70587;
    wire t70589 = t70588 ^ t70588;
    wire t70590 = t70589 ^ t70589;
    wire t70591 = t70590 ^ t70590;
    wire t70592 = t70591 ^ t70591;
    wire t70593 = t70592 ^ t70592;
    wire t70594 = t70593 ^ t70593;
    wire t70595 = t70594 ^ t70594;
    wire t70596 = t70595 ^ t70595;
    wire t70597 = t70596 ^ t70596;
    wire t70598 = t70597 ^ t70597;
    wire t70599 = t70598 ^ t70598;
    wire t70600 = t70599 ^ t70599;
    wire t70601 = t70600 ^ t70600;
    wire t70602 = t70601 ^ t70601;
    wire t70603 = t70602 ^ t70602;
    wire t70604 = t70603 ^ t70603;
    wire t70605 = t70604 ^ t70604;
    wire t70606 = t70605 ^ t70605;
    wire t70607 = t70606 ^ t70606;
    wire t70608 = t70607 ^ t70607;
    wire t70609 = t70608 ^ t70608;
    wire t70610 = t70609 ^ t70609;
    wire t70611 = t70610 ^ t70610;
    wire t70612 = t70611 ^ t70611;
    wire t70613 = t70612 ^ t70612;
    wire t70614 = t70613 ^ t70613;
    wire t70615 = t70614 ^ t70614;
    wire t70616 = t70615 ^ t70615;
    wire t70617 = t70616 ^ t70616;
    wire t70618 = t70617 ^ t70617;
    wire t70619 = t70618 ^ t70618;
    wire t70620 = t70619 ^ t70619;
    wire t70621 = t70620 ^ t70620;
    wire t70622 = t70621 ^ t70621;
    wire t70623 = t70622 ^ t70622;
    wire t70624 = t70623 ^ t70623;
    wire t70625 = t70624 ^ t70624;
    wire t70626 = t70625 ^ t70625;
    wire t70627 = t70626 ^ t70626;
    wire t70628 = t70627 ^ t70627;
    wire t70629 = t70628 ^ t70628;
    wire t70630 = t70629 ^ t70629;
    wire t70631 = t70630 ^ t70630;
    wire t70632 = t70631 ^ t70631;
    wire t70633 = t70632 ^ t70632;
    wire t70634 = t70633 ^ t70633;
    wire t70635 = t70634 ^ t70634;
    wire t70636 = t70635 ^ t70635;
    wire t70637 = t70636 ^ t70636;
    wire t70638 = t70637 ^ t70637;
    wire t70639 = t70638 ^ t70638;
    wire t70640 = t70639 ^ t70639;
    wire t70641 = t70640 ^ t70640;
    wire t70642 = t70641 ^ t70641;
    wire t70643 = t70642 ^ t70642;
    wire t70644 = t70643 ^ t70643;
    wire t70645 = t70644 ^ t70644;
    wire t70646 = t70645 ^ t70645;
    wire t70647 = t70646 ^ t70646;
    wire t70648 = t70647 ^ t70647;
    wire t70649 = t70648 ^ t70648;
    wire t70650 = t70649 ^ t70649;
    wire t70651 = t70650 ^ t70650;
    wire t70652 = t70651 ^ t70651;
    wire t70653 = t70652 ^ t70652;
    wire t70654 = t70653 ^ t70653;
    wire t70655 = t70654 ^ t70654;
    wire t70656 = t70655 ^ t70655;
    wire t70657 = t70656 ^ t70656;
    wire t70658 = t70657 ^ t70657;
    wire t70659 = t70658 ^ t70658;
    wire t70660 = t70659 ^ t70659;
    wire t70661 = t70660 ^ t70660;
    wire t70662 = t70661 ^ t70661;
    wire t70663 = t70662 ^ t70662;
    wire t70664 = t70663 ^ t70663;
    wire t70665 = t70664 ^ t70664;
    wire t70666 = t70665 ^ t70665;
    wire t70667 = t70666 ^ t70666;
    wire t70668 = t70667 ^ t70667;
    wire t70669 = t70668 ^ t70668;
    wire t70670 = t70669 ^ t70669;
    wire t70671 = t70670 ^ t70670;
    wire t70672 = t70671 ^ t70671;
    wire t70673 = t70672 ^ t70672;
    wire t70674 = t70673 ^ t70673;
    wire t70675 = t70674 ^ t70674;
    wire t70676 = t70675 ^ t70675;
    wire t70677 = t70676 ^ t70676;
    wire t70678 = t70677 ^ t70677;
    wire t70679 = t70678 ^ t70678;
    wire t70680 = t70679 ^ t70679;
    wire t70681 = t70680 ^ t70680;
    wire t70682 = t70681 ^ t70681;
    wire t70683 = t70682 ^ t70682;
    wire t70684 = t70683 ^ t70683;
    wire t70685 = t70684 ^ t70684;
    wire t70686 = t70685 ^ t70685;
    wire t70687 = t70686 ^ t70686;
    wire t70688 = t70687 ^ t70687;
    wire t70689 = t70688 ^ t70688;
    wire t70690 = t70689 ^ t70689;
    wire t70691 = t70690 ^ t70690;
    wire t70692 = t70691 ^ t70691;
    wire t70693 = t70692 ^ t70692;
    wire t70694 = t70693 ^ t70693;
    wire t70695 = t70694 ^ t70694;
    wire t70696 = t70695 ^ t70695;
    wire t70697 = t70696 ^ t70696;
    wire t70698 = t70697 ^ t70697;
    wire t70699 = t70698 ^ t70698;
    wire t70700 = t70699 ^ t70699;
    wire t70701 = t70700 ^ t70700;
    wire t70702 = t70701 ^ t70701;
    wire t70703 = t70702 ^ t70702;
    wire t70704 = t70703 ^ t70703;
    wire t70705 = t70704 ^ t70704;
    wire t70706 = t70705 ^ t70705;
    wire t70707 = t70706 ^ t70706;
    wire t70708 = t70707 ^ t70707;
    wire t70709 = t70708 ^ t70708;
    wire t70710 = t70709 ^ t70709;
    wire t70711 = t70710 ^ t70710;
    wire t70712 = t70711 ^ t70711;
    wire t70713 = t70712 ^ t70712;
    wire t70714 = t70713 ^ t70713;
    wire t70715 = t70714 ^ t70714;
    wire t70716 = t70715 ^ t70715;
    wire t70717 = t70716 ^ t70716;
    wire t70718 = t70717 ^ t70717;
    wire t70719 = t70718 ^ t70718;
    wire t70720 = t70719 ^ t70719;
    wire t70721 = t70720 ^ t70720;
    wire t70722 = t70721 ^ t70721;
    wire t70723 = t70722 ^ t70722;
    wire t70724 = t70723 ^ t70723;
    wire t70725 = t70724 ^ t70724;
    wire t70726 = t70725 ^ t70725;
    wire t70727 = t70726 ^ t70726;
    wire t70728 = t70727 ^ t70727;
    wire t70729 = t70728 ^ t70728;
    wire t70730 = t70729 ^ t70729;
    wire t70731 = t70730 ^ t70730;
    wire t70732 = t70731 ^ t70731;
    wire t70733 = t70732 ^ t70732;
    wire t70734 = t70733 ^ t70733;
    wire t70735 = t70734 ^ t70734;
    wire t70736 = t70735 ^ t70735;
    wire t70737 = t70736 ^ t70736;
    wire t70738 = t70737 ^ t70737;
    wire t70739 = t70738 ^ t70738;
    wire t70740 = t70739 ^ t70739;
    wire t70741 = t70740 ^ t70740;
    wire t70742 = t70741 ^ t70741;
    wire t70743 = t70742 ^ t70742;
    wire t70744 = t70743 ^ t70743;
    wire t70745 = t70744 ^ t70744;
    wire t70746 = t70745 ^ t70745;
    wire t70747 = t70746 ^ t70746;
    wire t70748 = t70747 ^ t70747;
    wire t70749 = t70748 ^ t70748;
    wire t70750 = t70749 ^ t70749;
    wire t70751 = t70750 ^ t70750;
    wire t70752 = t70751 ^ t70751;
    wire t70753 = t70752 ^ t70752;
    wire t70754 = t70753 ^ t70753;
    wire t70755 = t70754 ^ t70754;
    wire t70756 = t70755 ^ t70755;
    wire t70757 = t70756 ^ t70756;
    wire t70758 = t70757 ^ t70757;
    wire t70759 = t70758 ^ t70758;
    wire t70760 = t70759 ^ t70759;
    wire t70761 = t70760 ^ t70760;
    wire t70762 = t70761 ^ t70761;
    wire t70763 = t70762 ^ t70762;
    wire t70764 = t70763 ^ t70763;
    wire t70765 = t70764 ^ t70764;
    wire t70766 = t70765 ^ t70765;
    wire t70767 = t70766 ^ t70766;
    wire t70768 = t70767 ^ t70767;
    wire t70769 = t70768 ^ t70768;
    wire t70770 = t70769 ^ t70769;
    wire t70771 = t70770 ^ t70770;
    wire t70772 = t70771 ^ t70771;
    wire t70773 = t70772 ^ t70772;
    wire t70774 = t70773 ^ t70773;
    wire t70775 = t70774 ^ t70774;
    wire t70776 = t70775 ^ t70775;
    wire t70777 = t70776 ^ t70776;
    wire t70778 = t70777 ^ t70777;
    wire t70779 = t70778 ^ t70778;
    wire t70780 = t70779 ^ t70779;
    wire t70781 = t70780 ^ t70780;
    wire t70782 = t70781 ^ t70781;
    wire t70783 = t70782 ^ t70782;
    wire t70784 = t70783 ^ t70783;
    wire t70785 = t70784 ^ t70784;
    wire t70786 = t70785 ^ t70785;
    wire t70787 = t70786 ^ t70786;
    wire t70788 = t70787 ^ t70787;
    wire t70789 = t70788 ^ t70788;
    wire t70790 = t70789 ^ t70789;
    wire t70791 = t70790 ^ t70790;
    wire t70792 = t70791 ^ t70791;
    wire t70793 = t70792 ^ t70792;
    wire t70794 = t70793 ^ t70793;
    wire t70795 = t70794 ^ t70794;
    wire t70796 = t70795 ^ t70795;
    wire t70797 = t70796 ^ t70796;
    wire t70798 = t70797 ^ t70797;
    wire t70799 = t70798 ^ t70798;
    wire t70800 = t70799 ^ t70799;
    wire t70801 = t70800 ^ t70800;
    wire t70802 = t70801 ^ t70801;
    wire t70803 = t70802 ^ t70802;
    wire t70804 = t70803 ^ t70803;
    wire t70805 = t70804 ^ t70804;
    wire t70806 = t70805 ^ t70805;
    wire t70807 = t70806 ^ t70806;
    wire t70808 = t70807 ^ t70807;
    wire t70809 = t70808 ^ t70808;
    wire t70810 = t70809 ^ t70809;
    wire t70811 = t70810 ^ t70810;
    wire t70812 = t70811 ^ t70811;
    wire t70813 = t70812 ^ t70812;
    wire t70814 = t70813 ^ t70813;
    wire t70815 = t70814 ^ t70814;
    wire t70816 = t70815 ^ t70815;
    wire t70817 = t70816 ^ t70816;
    wire t70818 = t70817 ^ t70817;
    wire t70819 = t70818 ^ t70818;
    wire t70820 = t70819 ^ t70819;
    wire t70821 = t70820 ^ t70820;
    wire t70822 = t70821 ^ t70821;
    wire t70823 = t70822 ^ t70822;
    wire t70824 = t70823 ^ t70823;
    wire t70825 = t70824 ^ t70824;
    wire t70826 = t70825 ^ t70825;
    wire t70827 = t70826 ^ t70826;
    wire t70828 = t70827 ^ t70827;
    wire t70829 = t70828 ^ t70828;
    wire t70830 = t70829 ^ t70829;
    wire t70831 = t70830 ^ t70830;
    wire t70832 = t70831 ^ t70831;
    wire t70833 = t70832 ^ t70832;
    wire t70834 = t70833 ^ t70833;
    wire t70835 = t70834 ^ t70834;
    wire t70836 = t70835 ^ t70835;
    wire t70837 = t70836 ^ t70836;
    wire t70838 = t70837 ^ t70837;
    wire t70839 = t70838 ^ t70838;
    wire t70840 = t70839 ^ t70839;
    wire t70841 = t70840 ^ t70840;
    wire t70842 = t70841 ^ t70841;
    wire t70843 = t70842 ^ t70842;
    wire t70844 = t70843 ^ t70843;
    wire t70845 = t70844 ^ t70844;
    wire t70846 = t70845 ^ t70845;
    wire t70847 = t70846 ^ t70846;
    wire t70848 = t70847 ^ t70847;
    wire t70849 = t70848 ^ t70848;
    wire t70850 = t70849 ^ t70849;
    wire t70851 = t70850 ^ t70850;
    wire t70852 = t70851 ^ t70851;
    wire t70853 = t70852 ^ t70852;
    wire t70854 = t70853 ^ t70853;
    wire t70855 = t70854 ^ t70854;
    wire t70856 = t70855 ^ t70855;
    wire t70857 = t70856 ^ t70856;
    wire t70858 = t70857 ^ t70857;
    wire t70859 = t70858 ^ t70858;
    wire t70860 = t70859 ^ t70859;
    wire t70861 = t70860 ^ t70860;
    wire t70862 = t70861 ^ t70861;
    wire t70863 = t70862 ^ t70862;
    wire t70864 = t70863 ^ t70863;
    wire t70865 = t70864 ^ t70864;
    wire t70866 = t70865 ^ t70865;
    wire t70867 = t70866 ^ t70866;
    wire t70868 = t70867 ^ t70867;
    wire t70869 = t70868 ^ t70868;
    wire t70870 = t70869 ^ t70869;
    wire t70871 = t70870 ^ t70870;
    wire t70872 = t70871 ^ t70871;
    wire t70873 = t70872 ^ t70872;
    wire t70874 = t70873 ^ t70873;
    wire t70875 = t70874 ^ t70874;
    wire t70876 = t70875 ^ t70875;
    wire t70877 = t70876 ^ t70876;
    wire t70878 = t70877 ^ t70877;
    wire t70879 = t70878 ^ t70878;
    wire t70880 = t70879 ^ t70879;
    wire t70881 = t70880 ^ t70880;
    wire t70882 = t70881 ^ t70881;
    wire t70883 = t70882 ^ t70882;
    wire t70884 = t70883 ^ t70883;
    wire t70885 = t70884 ^ t70884;
    wire t70886 = t70885 ^ t70885;
    wire t70887 = t70886 ^ t70886;
    wire t70888 = t70887 ^ t70887;
    wire t70889 = t70888 ^ t70888;
    wire t70890 = t70889 ^ t70889;
    wire t70891 = t70890 ^ t70890;
    wire t70892 = t70891 ^ t70891;
    wire t70893 = t70892 ^ t70892;
    wire t70894 = t70893 ^ t70893;
    wire t70895 = t70894 ^ t70894;
    wire t70896 = t70895 ^ t70895;
    wire t70897 = t70896 ^ t70896;
    wire t70898 = t70897 ^ t70897;
    wire t70899 = t70898 ^ t70898;
    wire t70900 = t70899 ^ t70899;
    wire t70901 = t70900 ^ t70900;
    wire t70902 = t70901 ^ t70901;
    wire t70903 = t70902 ^ t70902;
    wire t70904 = t70903 ^ t70903;
    wire t70905 = t70904 ^ t70904;
    wire t70906 = t70905 ^ t70905;
    wire t70907 = t70906 ^ t70906;
    wire t70908 = t70907 ^ t70907;
    wire t70909 = t70908 ^ t70908;
    wire t70910 = t70909 ^ t70909;
    wire t70911 = t70910 ^ t70910;
    wire t70912 = t70911 ^ t70911;
    wire t70913 = t70912 ^ t70912;
    wire t70914 = t70913 ^ t70913;
    wire t70915 = t70914 ^ t70914;
    wire t70916 = t70915 ^ t70915;
    wire t70917 = t70916 ^ t70916;
    wire t70918 = t70917 ^ t70917;
    wire t70919 = t70918 ^ t70918;
    wire t70920 = t70919 ^ t70919;
    wire t70921 = t70920 ^ t70920;
    wire t70922 = t70921 ^ t70921;
    wire t70923 = t70922 ^ t70922;
    wire t70924 = t70923 ^ t70923;
    wire t70925 = t70924 ^ t70924;
    wire t70926 = t70925 ^ t70925;
    wire t70927 = t70926 ^ t70926;
    wire t70928 = t70927 ^ t70927;
    wire t70929 = t70928 ^ t70928;
    wire t70930 = t70929 ^ t70929;
    wire t70931 = t70930 ^ t70930;
    wire t70932 = t70931 ^ t70931;
    wire t70933 = t70932 ^ t70932;
    wire t70934 = t70933 ^ t70933;
    wire t70935 = t70934 ^ t70934;
    wire t70936 = t70935 ^ t70935;
    wire t70937 = t70936 ^ t70936;
    wire t70938 = t70937 ^ t70937;
    wire t70939 = t70938 ^ t70938;
    wire t70940 = t70939 ^ t70939;
    wire t70941 = t70940 ^ t70940;
    wire t70942 = t70941 ^ t70941;
    wire t70943 = t70942 ^ t70942;
    wire t70944 = t70943 ^ t70943;
    wire t70945 = t70944 ^ t70944;
    wire t70946 = t70945 ^ t70945;
    wire t70947 = t70946 ^ t70946;
    wire t70948 = t70947 ^ t70947;
    wire t70949 = t70948 ^ t70948;
    wire t70950 = t70949 ^ t70949;
    wire t70951 = t70950 ^ t70950;
    wire t70952 = t70951 ^ t70951;
    wire t70953 = t70952 ^ t70952;
    wire t70954 = t70953 ^ t70953;
    wire t70955 = t70954 ^ t70954;
    wire t70956 = t70955 ^ t70955;
    wire t70957 = t70956 ^ t70956;
    wire t70958 = t70957 ^ t70957;
    wire t70959 = t70958 ^ t70958;
    wire t70960 = t70959 ^ t70959;
    wire t70961 = t70960 ^ t70960;
    wire t70962 = t70961 ^ t70961;
    wire t70963 = t70962 ^ t70962;
    wire t70964 = t70963 ^ t70963;
    wire t70965 = t70964 ^ t70964;
    wire t70966 = t70965 ^ t70965;
    wire t70967 = t70966 ^ t70966;
    wire t70968 = t70967 ^ t70967;
    wire t70969 = t70968 ^ t70968;
    wire t70970 = t70969 ^ t70969;
    wire t70971 = t70970 ^ t70970;
    wire t70972 = t70971 ^ t70971;
    wire t70973 = t70972 ^ t70972;
    wire t70974 = t70973 ^ t70973;
    wire t70975 = t70974 ^ t70974;
    wire t70976 = t70975 ^ t70975;
    wire t70977 = t70976 ^ t70976;
    wire t70978 = t70977 ^ t70977;
    wire t70979 = t70978 ^ t70978;
    wire t70980 = t70979 ^ t70979;
    wire t70981 = t70980 ^ t70980;
    wire t70982 = t70981 ^ t70981;
    wire t70983 = t70982 ^ t70982;
    wire t70984 = t70983 ^ t70983;
    wire t70985 = t70984 ^ t70984;
    wire t70986 = t70985 ^ t70985;
    wire t70987 = t70986 ^ t70986;
    wire t70988 = t70987 ^ t70987;
    wire t70989 = t70988 ^ t70988;
    wire t70990 = t70989 ^ t70989;
    wire t70991 = t70990 ^ t70990;
    wire t70992 = t70991 ^ t70991;
    wire t70993 = t70992 ^ t70992;
    wire t70994 = t70993 ^ t70993;
    wire t70995 = t70994 ^ t70994;
    wire t70996 = t70995 ^ t70995;
    wire t70997 = t70996 ^ t70996;
    wire t70998 = t70997 ^ t70997;
    wire t70999 = t70998 ^ t70998;
    wire t71000 = t70999 ^ t70999;
    wire t71001 = t71000 ^ t71000;
    wire t71002 = t71001 ^ t71001;
    wire t71003 = t71002 ^ t71002;
    wire t71004 = t71003 ^ t71003;
    wire t71005 = t71004 ^ t71004;
    wire t71006 = t71005 ^ t71005;
    wire t71007 = t71006 ^ t71006;
    wire t71008 = t71007 ^ t71007;
    wire t71009 = t71008 ^ t71008;
    wire t71010 = t71009 ^ t71009;
    wire t71011 = t71010 ^ t71010;
    wire t71012 = t71011 ^ t71011;
    wire t71013 = t71012 ^ t71012;
    wire t71014 = t71013 ^ t71013;
    wire t71015 = t71014 ^ t71014;
    wire t71016 = t71015 ^ t71015;
    wire t71017 = t71016 ^ t71016;
    wire t71018 = t71017 ^ t71017;
    wire t71019 = t71018 ^ t71018;
    wire t71020 = t71019 ^ t71019;
    wire t71021 = t71020 ^ t71020;
    wire t71022 = t71021 ^ t71021;
    wire t71023 = t71022 ^ t71022;
    wire t71024 = t71023 ^ t71023;
    wire t71025 = t71024 ^ t71024;
    wire t71026 = t71025 ^ t71025;
    wire t71027 = t71026 ^ t71026;
    wire t71028 = t71027 ^ t71027;
    wire t71029 = t71028 ^ t71028;
    wire t71030 = t71029 ^ t71029;
    wire t71031 = t71030 ^ t71030;
    wire t71032 = t71031 ^ t71031;
    wire t71033 = t71032 ^ t71032;
    wire t71034 = t71033 ^ t71033;
    wire t71035 = t71034 ^ t71034;
    wire t71036 = t71035 ^ t71035;
    wire t71037 = t71036 ^ t71036;
    wire t71038 = t71037 ^ t71037;
    wire t71039 = t71038 ^ t71038;
    wire t71040 = t71039 ^ t71039;
    wire t71041 = t71040 ^ t71040;
    wire t71042 = t71041 ^ t71041;
    wire t71043 = t71042 ^ t71042;
    wire t71044 = t71043 ^ t71043;
    wire t71045 = t71044 ^ t71044;
    wire t71046 = t71045 ^ t71045;
    wire t71047 = t71046 ^ t71046;
    wire t71048 = t71047 ^ t71047;
    wire t71049 = t71048 ^ t71048;
    wire t71050 = t71049 ^ t71049;
    wire t71051 = t71050 ^ t71050;
    wire t71052 = t71051 ^ t71051;
    wire t71053 = t71052 ^ t71052;
    wire t71054 = t71053 ^ t71053;
    wire t71055 = t71054 ^ t71054;
    wire t71056 = t71055 ^ t71055;
    wire t71057 = t71056 ^ t71056;
    wire t71058 = t71057 ^ t71057;
    wire t71059 = t71058 ^ t71058;
    wire t71060 = t71059 ^ t71059;
    wire t71061 = t71060 ^ t71060;
    wire t71062 = t71061 ^ t71061;
    wire t71063 = t71062 ^ t71062;
    wire t71064 = t71063 ^ t71063;
    wire t71065 = t71064 ^ t71064;
    wire t71066 = t71065 ^ t71065;
    wire t71067 = t71066 ^ t71066;
    wire t71068 = t71067 ^ t71067;
    wire t71069 = t71068 ^ t71068;
    wire t71070 = t71069 ^ t71069;
    wire t71071 = t71070 ^ t71070;
    wire t71072 = t71071 ^ t71071;
    wire t71073 = t71072 ^ t71072;
    wire t71074 = t71073 ^ t71073;
    wire t71075 = t71074 ^ t71074;
    wire t71076 = t71075 ^ t71075;
    wire t71077 = t71076 ^ t71076;
    wire t71078 = t71077 ^ t71077;
    wire t71079 = t71078 ^ t71078;
    wire t71080 = t71079 ^ t71079;
    wire t71081 = t71080 ^ t71080;
    wire t71082 = t71081 ^ t71081;
    wire t71083 = t71082 ^ t71082;
    wire t71084 = t71083 ^ t71083;
    wire t71085 = t71084 ^ t71084;
    wire t71086 = t71085 ^ t71085;
    wire t71087 = t71086 ^ t71086;
    wire t71088 = t71087 ^ t71087;
    wire t71089 = t71088 ^ t71088;
    wire t71090 = t71089 ^ t71089;
    wire t71091 = t71090 ^ t71090;
    wire t71092 = t71091 ^ t71091;
    wire t71093 = t71092 ^ t71092;
    wire t71094 = t71093 ^ t71093;
    wire t71095 = t71094 ^ t71094;
    wire t71096 = t71095 ^ t71095;
    wire t71097 = t71096 ^ t71096;
    wire t71098 = t71097 ^ t71097;
    wire t71099 = t71098 ^ t71098;
    wire t71100 = t71099 ^ t71099;
    wire t71101 = t71100 ^ t71100;
    wire t71102 = t71101 ^ t71101;
    wire t71103 = t71102 ^ t71102;
    wire t71104 = t71103 ^ t71103;
    wire t71105 = t71104 ^ t71104;
    wire t71106 = t71105 ^ t71105;
    wire t71107 = t71106 ^ t71106;
    wire t71108 = t71107 ^ t71107;
    wire t71109 = t71108 ^ t71108;
    wire t71110 = t71109 ^ t71109;
    wire t71111 = t71110 ^ t71110;
    wire t71112 = t71111 ^ t71111;
    wire t71113 = t71112 ^ t71112;
    wire t71114 = t71113 ^ t71113;
    wire t71115 = t71114 ^ t71114;
    wire t71116 = t71115 ^ t71115;
    wire t71117 = t71116 ^ t71116;
    wire t71118 = t71117 ^ t71117;
    wire t71119 = t71118 ^ t71118;
    wire t71120 = t71119 ^ t71119;
    wire t71121 = t71120 ^ t71120;
    wire t71122 = t71121 ^ t71121;
    wire t71123 = t71122 ^ t71122;
    wire t71124 = t71123 ^ t71123;
    wire t71125 = t71124 ^ t71124;
    wire t71126 = t71125 ^ t71125;
    wire t71127 = t71126 ^ t71126;
    wire t71128 = t71127 ^ t71127;
    wire t71129 = t71128 ^ t71128;
    wire t71130 = t71129 ^ t71129;
    wire t71131 = t71130 ^ t71130;
    wire t71132 = t71131 ^ t71131;
    wire t71133 = t71132 ^ t71132;
    wire t71134 = t71133 ^ t71133;
    wire t71135 = t71134 ^ t71134;
    wire t71136 = t71135 ^ t71135;
    wire t71137 = t71136 ^ t71136;
    wire t71138 = t71137 ^ t71137;
    wire t71139 = t71138 ^ t71138;
    wire t71140 = t71139 ^ t71139;
    wire t71141 = t71140 ^ t71140;
    wire t71142 = t71141 ^ t71141;
    wire t71143 = t71142 ^ t71142;
    wire t71144 = t71143 ^ t71143;
    wire t71145 = t71144 ^ t71144;
    wire t71146 = t71145 ^ t71145;
    wire t71147 = t71146 ^ t71146;
    wire t71148 = t71147 ^ t71147;
    wire t71149 = t71148 ^ t71148;
    wire t71150 = t71149 ^ t71149;
    wire t71151 = t71150 ^ t71150;
    wire t71152 = t71151 ^ t71151;
    wire t71153 = t71152 ^ t71152;
    wire t71154 = t71153 ^ t71153;
    wire t71155 = t71154 ^ t71154;
    wire t71156 = t71155 ^ t71155;
    wire t71157 = t71156 ^ t71156;
    wire t71158 = t71157 ^ t71157;
    wire t71159 = t71158 ^ t71158;
    wire t71160 = t71159 ^ t71159;
    wire t71161 = t71160 ^ t71160;
    wire t71162 = t71161 ^ t71161;
    wire t71163 = t71162 ^ t71162;
    wire t71164 = t71163 ^ t71163;
    wire t71165 = t71164 ^ t71164;
    wire t71166 = t71165 ^ t71165;
    wire t71167 = t71166 ^ t71166;
    wire t71168 = t71167 ^ t71167;
    wire t71169 = t71168 ^ t71168;
    wire t71170 = t71169 ^ t71169;
    wire t71171 = t71170 ^ t71170;
    wire t71172 = t71171 ^ t71171;
    wire t71173 = t71172 ^ t71172;
    wire t71174 = t71173 ^ t71173;
    wire t71175 = t71174 ^ t71174;
    wire t71176 = t71175 ^ t71175;
    wire t71177 = t71176 ^ t71176;
    wire t71178 = t71177 ^ t71177;
    wire t71179 = t71178 ^ t71178;
    wire t71180 = t71179 ^ t71179;
    wire t71181 = t71180 ^ t71180;
    wire t71182 = t71181 ^ t71181;
    wire t71183 = t71182 ^ t71182;
    wire t71184 = t71183 ^ t71183;
    wire t71185 = t71184 ^ t71184;
    wire t71186 = t71185 ^ t71185;
    wire t71187 = t71186 ^ t71186;
    wire t71188 = t71187 ^ t71187;
    wire t71189 = t71188 ^ t71188;
    wire t71190 = t71189 ^ t71189;
    wire t71191 = t71190 ^ t71190;
    wire t71192 = t71191 ^ t71191;
    wire t71193 = t71192 ^ t71192;
    wire t71194 = t71193 ^ t71193;
    wire t71195 = t71194 ^ t71194;
    wire t71196 = t71195 ^ t71195;
    wire t71197 = t71196 ^ t71196;
    wire t71198 = t71197 ^ t71197;
    wire t71199 = t71198 ^ t71198;
    wire t71200 = t71199 ^ t71199;
    wire t71201 = t71200 ^ t71200;
    wire t71202 = t71201 ^ t71201;
    wire t71203 = t71202 ^ t71202;
    wire t71204 = t71203 ^ t71203;
    wire t71205 = t71204 ^ t71204;
    wire t71206 = t71205 ^ t71205;
    wire t71207 = t71206 ^ t71206;
    wire t71208 = t71207 ^ t71207;
    wire t71209 = t71208 ^ t71208;
    wire t71210 = t71209 ^ t71209;
    wire t71211 = t71210 ^ t71210;
    wire t71212 = t71211 ^ t71211;
    wire t71213 = t71212 ^ t71212;
    wire t71214 = t71213 ^ t71213;
    wire t71215 = t71214 ^ t71214;
    wire t71216 = t71215 ^ t71215;
    wire t71217 = t71216 ^ t71216;
    wire t71218 = t71217 ^ t71217;
    wire t71219 = t71218 ^ t71218;
    wire t71220 = t71219 ^ t71219;
    wire t71221 = t71220 ^ t71220;
    wire t71222 = t71221 ^ t71221;
    wire t71223 = t71222 ^ t71222;
    wire t71224 = t71223 ^ t71223;
    wire t71225 = t71224 ^ t71224;
    wire t71226 = t71225 ^ t71225;
    wire t71227 = t71226 ^ t71226;
    wire t71228 = t71227 ^ t71227;
    wire t71229 = t71228 ^ t71228;
    wire t71230 = t71229 ^ t71229;
    wire t71231 = t71230 ^ t71230;
    wire t71232 = t71231 ^ t71231;
    wire t71233 = t71232 ^ t71232;
    wire t71234 = t71233 ^ t71233;
    wire t71235 = t71234 ^ t71234;
    wire t71236 = t71235 ^ t71235;
    wire t71237 = t71236 ^ t71236;
    wire t71238 = t71237 ^ t71237;
    wire t71239 = t71238 ^ t71238;
    wire t71240 = t71239 ^ t71239;
    wire t71241 = t71240 ^ t71240;
    wire t71242 = t71241 ^ t71241;
    wire t71243 = t71242 ^ t71242;
    wire t71244 = t71243 ^ t71243;
    wire t71245 = t71244 ^ t71244;
    wire t71246 = t71245 ^ t71245;
    wire t71247 = t71246 ^ t71246;
    wire t71248 = t71247 ^ t71247;
    wire t71249 = t71248 ^ t71248;
    wire t71250 = t71249 ^ t71249;
    wire t71251 = t71250 ^ t71250;
    wire t71252 = t71251 ^ t71251;
    wire t71253 = t71252 ^ t71252;
    wire t71254 = t71253 ^ t71253;
    wire t71255 = t71254 ^ t71254;
    wire t71256 = t71255 ^ t71255;
    wire t71257 = t71256 ^ t71256;
    wire t71258 = t71257 ^ t71257;
    wire t71259 = t71258 ^ t71258;
    wire t71260 = t71259 ^ t71259;
    wire t71261 = t71260 ^ t71260;
    wire t71262 = t71261 ^ t71261;
    wire t71263 = t71262 ^ t71262;
    wire t71264 = t71263 ^ t71263;
    wire t71265 = t71264 ^ t71264;
    wire t71266 = t71265 ^ t71265;
    wire t71267 = t71266 ^ t71266;
    wire t71268 = t71267 ^ t71267;
    wire t71269 = t71268 ^ t71268;
    wire t71270 = t71269 ^ t71269;
    wire t71271 = t71270 ^ t71270;
    wire t71272 = t71271 ^ t71271;
    wire t71273 = t71272 ^ t71272;
    wire t71274 = t71273 ^ t71273;
    wire t71275 = t71274 ^ t71274;
    wire t71276 = t71275 ^ t71275;
    wire t71277 = t71276 ^ t71276;
    wire t71278 = t71277 ^ t71277;
    wire t71279 = t71278 ^ t71278;
    wire t71280 = t71279 ^ t71279;
    wire t71281 = t71280 ^ t71280;
    wire t71282 = t71281 ^ t71281;
    wire t71283 = t71282 ^ t71282;
    wire t71284 = t71283 ^ t71283;
    wire t71285 = t71284 ^ t71284;
    wire t71286 = t71285 ^ t71285;
    wire t71287 = t71286 ^ t71286;
    wire t71288 = t71287 ^ t71287;
    wire t71289 = t71288 ^ t71288;
    wire t71290 = t71289 ^ t71289;
    wire t71291 = t71290 ^ t71290;
    wire t71292 = t71291 ^ t71291;
    wire t71293 = t71292 ^ t71292;
    wire t71294 = t71293 ^ t71293;
    wire t71295 = t71294 ^ t71294;
    wire t71296 = t71295 ^ t71295;
    wire t71297 = t71296 ^ t71296;
    wire t71298 = t71297 ^ t71297;
    wire t71299 = t71298 ^ t71298;
    wire t71300 = t71299 ^ t71299;
    wire t71301 = t71300 ^ t71300;
    wire t71302 = t71301 ^ t71301;
    wire t71303 = t71302 ^ t71302;
    wire t71304 = t71303 ^ t71303;
    wire t71305 = t71304 ^ t71304;
    wire t71306 = t71305 ^ t71305;
    wire t71307 = t71306 ^ t71306;
    wire t71308 = t71307 ^ t71307;
    wire t71309 = t71308 ^ t71308;
    wire t71310 = t71309 ^ t71309;
    wire t71311 = t71310 ^ t71310;
    wire t71312 = t71311 ^ t71311;
    wire t71313 = t71312 ^ t71312;
    wire t71314 = t71313 ^ t71313;
    wire t71315 = t71314 ^ t71314;
    wire t71316 = t71315 ^ t71315;
    wire t71317 = t71316 ^ t71316;
    wire t71318 = t71317 ^ t71317;
    wire t71319 = t71318 ^ t71318;
    wire t71320 = t71319 ^ t71319;
    wire t71321 = t71320 ^ t71320;
    wire t71322 = t71321 ^ t71321;
    wire t71323 = t71322 ^ t71322;
    wire t71324 = t71323 ^ t71323;
    wire t71325 = t71324 ^ t71324;
    wire t71326 = t71325 ^ t71325;
    wire t71327 = t71326 ^ t71326;
    wire t71328 = t71327 ^ t71327;
    wire t71329 = t71328 ^ t71328;
    wire t71330 = t71329 ^ t71329;
    wire t71331 = t71330 ^ t71330;
    wire t71332 = t71331 ^ t71331;
    wire t71333 = t71332 ^ t71332;
    wire t71334 = t71333 ^ t71333;
    wire t71335 = t71334 ^ t71334;
    wire t71336 = t71335 ^ t71335;
    wire t71337 = t71336 ^ t71336;
    wire t71338 = t71337 ^ t71337;
    wire t71339 = t71338 ^ t71338;
    wire t71340 = t71339 ^ t71339;
    wire t71341 = t71340 ^ t71340;
    wire t71342 = t71341 ^ t71341;
    wire t71343 = t71342 ^ t71342;
    wire t71344 = t71343 ^ t71343;
    wire t71345 = t71344 ^ t71344;
    wire t71346 = t71345 ^ t71345;
    wire t71347 = t71346 ^ t71346;
    wire t71348 = t71347 ^ t71347;
    wire t71349 = t71348 ^ t71348;
    wire t71350 = t71349 ^ t71349;
    wire t71351 = t71350 ^ t71350;
    wire t71352 = t71351 ^ t71351;
    wire t71353 = t71352 ^ t71352;
    wire t71354 = t71353 ^ t71353;
    wire t71355 = t71354 ^ t71354;
    wire t71356 = t71355 ^ t71355;
    wire t71357 = t71356 ^ t71356;
    wire t71358 = t71357 ^ t71357;
    wire t71359 = t71358 ^ t71358;
    wire t71360 = t71359 ^ t71359;
    wire t71361 = t71360 ^ t71360;
    wire t71362 = t71361 ^ t71361;
    wire t71363 = t71362 ^ t71362;
    wire t71364 = t71363 ^ t71363;
    wire t71365 = t71364 ^ t71364;
    wire t71366 = t71365 ^ t71365;
    wire t71367 = t71366 ^ t71366;
    wire t71368 = t71367 ^ t71367;
    wire t71369 = t71368 ^ t71368;
    wire t71370 = t71369 ^ t71369;
    wire t71371 = t71370 ^ t71370;
    wire t71372 = t71371 ^ t71371;
    wire t71373 = t71372 ^ t71372;
    wire t71374 = t71373 ^ t71373;
    wire t71375 = t71374 ^ t71374;
    wire t71376 = t71375 ^ t71375;
    wire t71377 = t71376 ^ t71376;
    wire t71378 = t71377 ^ t71377;
    wire t71379 = t71378 ^ t71378;
    wire t71380 = t71379 ^ t71379;
    wire t71381 = t71380 ^ t71380;
    wire t71382 = t71381 ^ t71381;
    wire t71383 = t71382 ^ t71382;
    wire t71384 = t71383 ^ t71383;
    wire t71385 = t71384 ^ t71384;
    wire t71386 = t71385 ^ t71385;
    wire t71387 = t71386 ^ t71386;
    wire t71388 = t71387 ^ t71387;
    wire t71389 = t71388 ^ t71388;
    wire t71390 = t71389 ^ t71389;
    wire t71391 = t71390 ^ t71390;
    wire t71392 = t71391 ^ t71391;
    wire t71393 = t71392 ^ t71392;
    wire t71394 = t71393 ^ t71393;
    wire t71395 = t71394 ^ t71394;
    wire t71396 = t71395 ^ t71395;
    wire t71397 = t71396 ^ t71396;
    wire t71398 = t71397 ^ t71397;
    wire t71399 = t71398 ^ t71398;
    wire t71400 = t71399 ^ t71399;
    wire t71401 = t71400 ^ t71400;
    wire t71402 = t71401 ^ t71401;
    wire t71403 = t71402 ^ t71402;
    wire t71404 = t71403 ^ t71403;
    wire t71405 = t71404 ^ t71404;
    wire t71406 = t71405 ^ t71405;
    wire t71407 = t71406 ^ t71406;
    wire t71408 = t71407 ^ t71407;
    wire t71409 = t71408 ^ t71408;
    wire t71410 = t71409 ^ t71409;
    wire t71411 = t71410 ^ t71410;
    wire t71412 = t71411 ^ t71411;
    wire t71413 = t71412 ^ t71412;
    wire t71414 = t71413 ^ t71413;
    wire t71415 = t71414 ^ t71414;
    wire t71416 = t71415 ^ t71415;
    wire t71417 = t71416 ^ t71416;
    wire t71418 = t71417 ^ t71417;
    wire t71419 = t71418 ^ t71418;
    wire t71420 = t71419 ^ t71419;
    wire t71421 = t71420 ^ t71420;
    wire t71422 = t71421 ^ t71421;
    wire t71423 = t71422 ^ t71422;
    wire t71424 = t71423 ^ t71423;
    wire t71425 = t71424 ^ t71424;
    wire t71426 = t71425 ^ t71425;
    wire t71427 = t71426 ^ t71426;
    wire t71428 = t71427 ^ t71427;
    wire t71429 = t71428 ^ t71428;
    wire t71430 = t71429 ^ t71429;
    wire t71431 = t71430 ^ t71430;
    wire t71432 = t71431 ^ t71431;
    wire t71433 = t71432 ^ t71432;
    wire t71434 = t71433 ^ t71433;
    wire t71435 = t71434 ^ t71434;
    wire t71436 = t71435 ^ t71435;
    wire t71437 = t71436 ^ t71436;
    wire t71438 = t71437 ^ t71437;
    wire t71439 = t71438 ^ t71438;
    wire t71440 = t71439 ^ t71439;
    wire t71441 = t71440 ^ t71440;
    wire t71442 = t71441 ^ t71441;
    wire t71443 = t71442 ^ t71442;
    wire t71444 = t71443 ^ t71443;
    wire t71445 = t71444 ^ t71444;
    wire t71446 = t71445 ^ t71445;
    wire t71447 = t71446 ^ t71446;
    wire t71448 = t71447 ^ t71447;
    wire t71449 = t71448 ^ t71448;
    wire t71450 = t71449 ^ t71449;
    wire t71451 = t71450 ^ t71450;
    wire t71452 = t71451 ^ t71451;
    wire t71453 = t71452 ^ t71452;
    wire t71454 = t71453 ^ t71453;
    wire t71455 = t71454 ^ t71454;
    wire t71456 = t71455 ^ t71455;
    wire t71457 = t71456 ^ t71456;
    wire t71458 = t71457 ^ t71457;
    wire t71459 = t71458 ^ t71458;
    wire t71460 = t71459 ^ t71459;
    wire t71461 = t71460 ^ t71460;
    wire t71462 = t71461 ^ t71461;
    wire t71463 = t71462 ^ t71462;
    wire t71464 = t71463 ^ t71463;
    wire t71465 = t71464 ^ t71464;
    wire t71466 = t71465 ^ t71465;
    wire t71467 = t71466 ^ t71466;
    wire t71468 = t71467 ^ t71467;
    wire t71469 = t71468 ^ t71468;
    wire t71470 = t71469 ^ t71469;
    wire t71471 = t71470 ^ t71470;
    wire t71472 = t71471 ^ t71471;
    wire t71473 = t71472 ^ t71472;
    wire t71474 = t71473 ^ t71473;
    wire t71475 = t71474 ^ t71474;
    wire t71476 = t71475 ^ t71475;
    wire t71477 = t71476 ^ t71476;
    wire t71478 = t71477 ^ t71477;
    wire t71479 = t71478 ^ t71478;
    wire t71480 = t71479 ^ t71479;
    wire t71481 = t71480 ^ t71480;
    wire t71482 = t71481 ^ t71481;
    wire t71483 = t71482 ^ t71482;
    wire t71484 = t71483 ^ t71483;
    wire t71485 = t71484 ^ t71484;
    wire t71486 = t71485 ^ t71485;
    wire t71487 = t71486 ^ t71486;
    wire t71488 = t71487 ^ t71487;
    wire t71489 = t71488 ^ t71488;
    wire t71490 = t71489 ^ t71489;
    wire t71491 = t71490 ^ t71490;
    wire t71492 = t71491 ^ t71491;
    wire t71493 = t71492 ^ t71492;
    wire t71494 = t71493 ^ t71493;
    wire t71495 = t71494 ^ t71494;
    wire t71496 = t71495 ^ t71495;
    wire t71497 = t71496 ^ t71496;
    wire t71498 = t71497 ^ t71497;
    wire t71499 = t71498 ^ t71498;
    wire t71500 = t71499 ^ t71499;
    wire t71501 = t71500 ^ t71500;
    wire t71502 = t71501 ^ t71501;
    wire t71503 = t71502 ^ t71502;
    wire t71504 = t71503 ^ t71503;
    wire t71505 = t71504 ^ t71504;
    wire t71506 = t71505 ^ t71505;
    wire t71507 = t71506 ^ t71506;
    wire t71508 = t71507 ^ t71507;
    wire t71509 = t71508 ^ t71508;
    wire t71510 = t71509 ^ t71509;
    wire t71511 = t71510 ^ t71510;
    wire t71512 = t71511 ^ t71511;
    wire t71513 = t71512 ^ t71512;
    wire t71514 = t71513 ^ t71513;
    wire t71515 = t71514 ^ t71514;
    wire t71516 = t71515 ^ t71515;
    wire t71517 = t71516 ^ t71516;
    wire t71518 = t71517 ^ t71517;
    wire t71519 = t71518 ^ t71518;
    wire t71520 = t71519 ^ t71519;
    wire t71521 = t71520 ^ t71520;
    wire t71522 = t71521 ^ t71521;
    wire t71523 = t71522 ^ t71522;
    wire t71524 = t71523 ^ t71523;
    wire t71525 = t71524 ^ t71524;
    wire t71526 = t71525 ^ t71525;
    wire t71527 = t71526 ^ t71526;
    wire t71528 = t71527 ^ t71527;
    wire t71529 = t71528 ^ t71528;
    wire t71530 = t71529 ^ t71529;
    wire t71531 = t71530 ^ t71530;
    wire t71532 = t71531 ^ t71531;
    wire t71533 = t71532 ^ t71532;
    wire t71534 = t71533 ^ t71533;
    wire t71535 = t71534 ^ t71534;
    wire t71536 = t71535 ^ t71535;
    wire t71537 = t71536 ^ t71536;
    wire t71538 = t71537 ^ t71537;
    wire t71539 = t71538 ^ t71538;
    wire t71540 = t71539 ^ t71539;
    wire t71541 = t71540 ^ t71540;
    wire t71542 = t71541 ^ t71541;
    wire t71543 = t71542 ^ t71542;
    wire t71544 = t71543 ^ t71543;
    wire t71545 = t71544 ^ t71544;
    wire t71546 = t71545 ^ t71545;
    wire t71547 = t71546 ^ t71546;
    wire t71548 = t71547 ^ t71547;
    wire t71549 = t71548 ^ t71548;
    wire t71550 = t71549 ^ t71549;
    wire t71551 = t71550 ^ t71550;
    wire t71552 = t71551 ^ t71551;
    wire t71553 = t71552 ^ t71552;
    wire t71554 = t71553 ^ t71553;
    wire t71555 = t71554 ^ t71554;
    wire t71556 = t71555 ^ t71555;
    wire t71557 = t71556 ^ t71556;
    wire t71558 = t71557 ^ t71557;
    wire t71559 = t71558 ^ t71558;
    wire t71560 = t71559 ^ t71559;
    wire t71561 = t71560 ^ t71560;
    wire t71562 = t71561 ^ t71561;
    wire t71563 = t71562 ^ t71562;
    wire t71564 = t71563 ^ t71563;
    wire t71565 = t71564 ^ t71564;
    wire t71566 = t71565 ^ t71565;
    wire t71567 = t71566 ^ t71566;
    wire t71568 = t71567 ^ t71567;
    wire t71569 = t71568 ^ t71568;
    wire t71570 = t71569 ^ t71569;
    wire t71571 = t71570 ^ t71570;
    wire t71572 = t71571 ^ t71571;
    wire t71573 = t71572 ^ t71572;
    wire t71574 = t71573 ^ t71573;
    wire t71575 = t71574 ^ t71574;
    wire t71576 = t71575 ^ t71575;
    wire t71577 = t71576 ^ t71576;
    wire t71578 = t71577 ^ t71577;
    wire t71579 = t71578 ^ t71578;
    wire t71580 = t71579 ^ t71579;
    wire t71581 = t71580 ^ t71580;
    wire t71582 = t71581 ^ t71581;
    wire t71583 = t71582 ^ t71582;
    wire t71584 = t71583 ^ t71583;
    wire t71585 = t71584 ^ t71584;
    wire t71586 = t71585 ^ t71585;
    wire t71587 = t71586 ^ t71586;
    wire t71588 = t71587 ^ t71587;
    wire t71589 = t71588 ^ t71588;
    wire t71590 = t71589 ^ t71589;
    wire t71591 = t71590 ^ t71590;
    wire t71592 = t71591 ^ t71591;
    wire t71593 = t71592 ^ t71592;
    wire t71594 = t71593 ^ t71593;
    wire t71595 = t71594 ^ t71594;
    wire t71596 = t71595 ^ t71595;
    wire t71597 = t71596 ^ t71596;
    wire t71598 = t71597 ^ t71597;
    wire t71599 = t71598 ^ t71598;
    wire t71600 = t71599 ^ t71599;
    wire t71601 = t71600 ^ t71600;
    wire t71602 = t71601 ^ t71601;
    wire t71603 = t71602 ^ t71602;
    wire t71604 = t71603 ^ t71603;
    wire t71605 = t71604 ^ t71604;
    wire t71606 = t71605 ^ t71605;
    wire t71607 = t71606 ^ t71606;
    wire t71608 = t71607 ^ t71607;
    wire t71609 = t71608 ^ t71608;
    wire t71610 = t71609 ^ t71609;
    wire t71611 = t71610 ^ t71610;
    wire t71612 = t71611 ^ t71611;
    wire t71613 = t71612 ^ t71612;
    wire t71614 = t71613 ^ t71613;
    wire t71615 = t71614 ^ t71614;
    wire t71616 = t71615 ^ t71615;
    wire t71617 = t71616 ^ t71616;
    wire t71618 = t71617 ^ t71617;
    wire t71619 = t71618 ^ t71618;
    wire t71620 = t71619 ^ t71619;
    wire t71621 = t71620 ^ t71620;
    wire t71622 = t71621 ^ t71621;
    wire t71623 = t71622 ^ t71622;
    wire t71624 = t71623 ^ t71623;
    wire t71625 = t71624 ^ t71624;
    wire t71626 = t71625 ^ t71625;
    wire t71627 = t71626 ^ t71626;
    wire t71628 = t71627 ^ t71627;
    wire t71629 = t71628 ^ t71628;
    wire t71630 = t71629 ^ t71629;
    wire t71631 = t71630 ^ t71630;
    wire t71632 = t71631 ^ t71631;
    wire t71633 = t71632 ^ t71632;
    wire t71634 = t71633 ^ t71633;
    wire t71635 = t71634 ^ t71634;
    wire t71636 = t71635 ^ t71635;
    wire t71637 = t71636 ^ t71636;
    wire t71638 = t71637 ^ t71637;
    wire t71639 = t71638 ^ t71638;
    wire t71640 = t71639 ^ t71639;
    wire t71641 = t71640 ^ t71640;
    wire t71642 = t71641 ^ t71641;
    wire t71643 = t71642 ^ t71642;
    wire t71644 = t71643 ^ t71643;
    wire t71645 = t71644 ^ t71644;
    wire t71646 = t71645 ^ t71645;
    wire t71647 = t71646 ^ t71646;
    wire t71648 = t71647 ^ t71647;
    wire t71649 = t71648 ^ t71648;
    wire t71650 = t71649 ^ t71649;
    wire t71651 = t71650 ^ t71650;
    wire t71652 = t71651 ^ t71651;
    wire t71653 = t71652 ^ t71652;
    wire t71654 = t71653 ^ t71653;
    wire t71655 = t71654 ^ t71654;
    wire t71656 = t71655 ^ t71655;
    wire t71657 = t71656 ^ t71656;
    wire t71658 = t71657 ^ t71657;
    wire t71659 = t71658 ^ t71658;
    wire t71660 = t71659 ^ t71659;
    wire t71661 = t71660 ^ t71660;
    wire t71662 = t71661 ^ t71661;
    wire t71663 = t71662 ^ t71662;
    wire t71664 = t71663 ^ t71663;
    wire t71665 = t71664 ^ t71664;
    wire t71666 = t71665 ^ t71665;
    wire t71667 = t71666 ^ t71666;
    wire t71668 = t71667 ^ t71667;
    wire t71669 = t71668 ^ t71668;
    wire t71670 = t71669 ^ t71669;
    wire t71671 = t71670 ^ t71670;
    wire t71672 = t71671 ^ t71671;
    wire t71673 = t71672 ^ t71672;
    wire t71674 = t71673 ^ t71673;
    wire t71675 = t71674 ^ t71674;
    wire t71676 = t71675 ^ t71675;
    wire t71677 = t71676 ^ t71676;
    wire t71678 = t71677 ^ t71677;
    wire t71679 = t71678 ^ t71678;
    wire t71680 = t71679 ^ t71679;
    wire t71681 = t71680 ^ t71680;
    wire t71682 = t71681 ^ t71681;
    wire t71683 = t71682 ^ t71682;
    wire t71684 = t71683 ^ t71683;
    wire t71685 = t71684 ^ t71684;
    wire t71686 = t71685 ^ t71685;
    wire t71687 = t71686 ^ t71686;
    wire t71688 = t71687 ^ t71687;
    wire t71689 = t71688 ^ t71688;
    wire t71690 = t71689 ^ t71689;
    wire t71691 = t71690 ^ t71690;
    wire t71692 = t71691 ^ t71691;
    wire t71693 = t71692 ^ t71692;
    wire t71694 = t71693 ^ t71693;
    wire t71695 = t71694 ^ t71694;
    wire t71696 = t71695 ^ t71695;
    wire t71697 = t71696 ^ t71696;
    wire t71698 = t71697 ^ t71697;
    wire t71699 = t71698 ^ t71698;
    wire t71700 = t71699 ^ t71699;
    wire t71701 = t71700 ^ t71700;
    wire t71702 = t71701 ^ t71701;
    wire t71703 = t71702 ^ t71702;
    wire t71704 = t71703 ^ t71703;
    wire t71705 = t71704 ^ t71704;
    wire t71706 = t71705 ^ t71705;
    wire t71707 = t71706 ^ t71706;
    wire t71708 = t71707 ^ t71707;
    wire t71709 = t71708 ^ t71708;
    wire t71710 = t71709 ^ t71709;
    wire t71711 = t71710 ^ t71710;
    wire t71712 = t71711 ^ t71711;
    wire t71713 = t71712 ^ t71712;
    wire t71714 = t71713 ^ t71713;
    wire t71715 = t71714 ^ t71714;
    wire t71716 = t71715 ^ t71715;
    wire t71717 = t71716 ^ t71716;
    wire t71718 = t71717 ^ t71717;
    wire t71719 = t71718 ^ t71718;
    wire t71720 = t71719 ^ t71719;
    wire t71721 = t71720 ^ t71720;
    wire t71722 = t71721 ^ t71721;
    wire t71723 = t71722 ^ t71722;
    wire t71724 = t71723 ^ t71723;
    wire t71725 = t71724 ^ t71724;
    wire t71726 = t71725 ^ t71725;
    wire t71727 = t71726 ^ t71726;
    wire t71728 = t71727 ^ t71727;
    wire t71729 = t71728 ^ t71728;
    wire t71730 = t71729 ^ t71729;
    wire t71731 = t71730 ^ t71730;
    wire t71732 = t71731 ^ t71731;
    wire t71733 = t71732 ^ t71732;
    wire t71734 = t71733 ^ t71733;
    wire t71735 = t71734 ^ t71734;
    wire t71736 = t71735 ^ t71735;
    wire t71737 = t71736 ^ t71736;
    wire t71738 = t71737 ^ t71737;
    wire t71739 = t71738 ^ t71738;
    wire t71740 = t71739 ^ t71739;
    wire t71741 = t71740 ^ t71740;
    wire t71742 = t71741 ^ t71741;
    wire t71743 = t71742 ^ t71742;
    wire t71744 = t71743 ^ t71743;
    wire t71745 = t71744 ^ t71744;
    wire t71746 = t71745 ^ t71745;
    wire t71747 = t71746 ^ t71746;
    wire t71748 = t71747 ^ t71747;
    wire t71749 = t71748 ^ t71748;
    wire t71750 = t71749 ^ t71749;
    wire t71751 = t71750 ^ t71750;
    wire t71752 = t71751 ^ t71751;
    wire t71753 = t71752 ^ t71752;
    wire t71754 = t71753 ^ t71753;
    wire t71755 = t71754 ^ t71754;
    wire t71756 = t71755 ^ t71755;
    wire t71757 = t71756 ^ t71756;
    wire t71758 = t71757 ^ t71757;
    wire t71759 = t71758 ^ t71758;
    wire t71760 = t71759 ^ t71759;
    wire t71761 = t71760 ^ t71760;
    wire t71762 = t71761 ^ t71761;
    wire t71763 = t71762 ^ t71762;
    wire t71764 = t71763 ^ t71763;
    wire t71765 = t71764 ^ t71764;
    wire t71766 = t71765 ^ t71765;
    wire t71767 = t71766 ^ t71766;
    wire t71768 = t71767 ^ t71767;
    wire t71769 = t71768 ^ t71768;
    wire t71770 = t71769 ^ t71769;
    wire t71771 = t71770 ^ t71770;
    wire t71772 = t71771 ^ t71771;
    wire t71773 = t71772 ^ t71772;
    wire t71774 = t71773 ^ t71773;
    wire t71775 = t71774 ^ t71774;
    wire t71776 = t71775 ^ t71775;
    wire t71777 = t71776 ^ t71776;
    wire t71778 = t71777 ^ t71777;
    wire t71779 = t71778 ^ t71778;
    wire t71780 = t71779 ^ t71779;
    wire t71781 = t71780 ^ t71780;
    wire t71782 = t71781 ^ t71781;
    wire t71783 = t71782 ^ t71782;
    wire t71784 = t71783 ^ t71783;
    wire t71785 = t71784 ^ t71784;
    wire t71786 = t71785 ^ t71785;
    wire t71787 = t71786 ^ t71786;
    wire t71788 = t71787 ^ t71787;
    wire t71789 = t71788 ^ t71788;
    wire t71790 = t71789 ^ t71789;
    wire t71791 = t71790 ^ t71790;
    wire t71792 = t71791 ^ t71791;
    wire t71793 = t71792 ^ t71792;
    wire t71794 = t71793 ^ t71793;
    wire t71795 = t71794 ^ t71794;
    wire t71796 = t71795 ^ t71795;
    wire t71797 = t71796 ^ t71796;
    wire t71798 = t71797 ^ t71797;
    wire t71799 = t71798 ^ t71798;
    wire t71800 = t71799 ^ t71799;
    wire t71801 = t71800 ^ t71800;
    wire t71802 = t71801 ^ t71801;
    wire t71803 = t71802 ^ t71802;
    wire t71804 = t71803 ^ t71803;
    wire t71805 = t71804 ^ t71804;
    wire t71806 = t71805 ^ t71805;
    wire t71807 = t71806 ^ t71806;
    wire t71808 = t71807 ^ t71807;
    wire t71809 = t71808 ^ t71808;
    wire t71810 = t71809 ^ t71809;
    wire t71811 = t71810 ^ t71810;
    wire t71812 = t71811 ^ t71811;
    wire t71813 = t71812 ^ t71812;
    wire t71814 = t71813 ^ t71813;
    wire t71815 = t71814 ^ t71814;
    wire t71816 = t71815 ^ t71815;
    wire t71817 = t71816 ^ t71816;
    wire t71818 = t71817 ^ t71817;
    wire t71819 = t71818 ^ t71818;
    wire t71820 = t71819 ^ t71819;
    wire t71821 = t71820 ^ t71820;
    wire t71822 = t71821 ^ t71821;
    wire t71823 = t71822 ^ t71822;
    wire t71824 = t71823 ^ t71823;
    wire t71825 = t71824 ^ t71824;
    wire t71826 = t71825 ^ t71825;
    wire t71827 = t71826 ^ t71826;
    wire t71828 = t71827 ^ t71827;
    wire t71829 = t71828 ^ t71828;
    wire t71830 = t71829 ^ t71829;
    wire t71831 = t71830 ^ t71830;
    wire t71832 = t71831 ^ t71831;
    wire t71833 = t71832 ^ t71832;
    wire t71834 = t71833 ^ t71833;
    wire t71835 = t71834 ^ t71834;
    wire t71836 = t71835 ^ t71835;
    wire t71837 = t71836 ^ t71836;
    wire t71838 = t71837 ^ t71837;
    wire t71839 = t71838 ^ t71838;
    wire t71840 = t71839 ^ t71839;
    wire t71841 = t71840 ^ t71840;
    wire t71842 = t71841 ^ t71841;
    wire t71843 = t71842 ^ t71842;
    wire t71844 = t71843 ^ t71843;
    wire t71845 = t71844 ^ t71844;
    wire t71846 = t71845 ^ t71845;
    wire t71847 = t71846 ^ t71846;
    wire t71848 = t71847 ^ t71847;
    wire t71849 = t71848 ^ t71848;
    wire t71850 = t71849 ^ t71849;
    wire t71851 = t71850 ^ t71850;
    wire t71852 = t71851 ^ t71851;
    wire t71853 = t71852 ^ t71852;
    wire t71854 = t71853 ^ t71853;
    wire t71855 = t71854 ^ t71854;
    wire t71856 = t71855 ^ t71855;
    wire t71857 = t71856 ^ t71856;
    wire t71858 = t71857 ^ t71857;
    wire t71859 = t71858 ^ t71858;
    wire t71860 = t71859 ^ t71859;
    wire t71861 = t71860 ^ t71860;
    wire t71862 = t71861 ^ t71861;
    wire t71863 = t71862 ^ t71862;
    wire t71864 = t71863 ^ t71863;
    wire t71865 = t71864 ^ t71864;
    wire t71866 = t71865 ^ t71865;
    wire t71867 = t71866 ^ t71866;
    wire t71868 = t71867 ^ t71867;
    wire t71869 = t71868 ^ t71868;
    wire t71870 = t71869 ^ t71869;
    wire t71871 = t71870 ^ t71870;
    wire t71872 = t71871 ^ t71871;
    wire t71873 = t71872 ^ t71872;
    wire t71874 = t71873 ^ t71873;
    wire t71875 = t71874 ^ t71874;
    wire t71876 = t71875 ^ t71875;
    wire t71877 = t71876 ^ t71876;
    wire t71878 = t71877 ^ t71877;
    wire t71879 = t71878 ^ t71878;
    wire t71880 = t71879 ^ t71879;
    wire t71881 = t71880 ^ t71880;
    wire t71882 = t71881 ^ t71881;
    wire t71883 = t71882 ^ t71882;
    wire t71884 = t71883 ^ t71883;
    wire t71885 = t71884 ^ t71884;
    wire t71886 = t71885 ^ t71885;
    wire t71887 = t71886 ^ t71886;
    wire t71888 = t71887 ^ t71887;
    wire t71889 = t71888 ^ t71888;
    wire t71890 = t71889 ^ t71889;
    wire t71891 = t71890 ^ t71890;
    wire t71892 = t71891 ^ t71891;
    wire t71893 = t71892 ^ t71892;
    wire t71894 = t71893 ^ t71893;
    wire t71895 = t71894 ^ t71894;
    wire t71896 = t71895 ^ t71895;
    wire t71897 = t71896 ^ t71896;
    wire t71898 = t71897 ^ t71897;
    wire t71899 = t71898 ^ t71898;
    wire t71900 = t71899 ^ t71899;
    wire t71901 = t71900 ^ t71900;
    wire t71902 = t71901 ^ t71901;
    wire t71903 = t71902 ^ t71902;
    wire t71904 = t71903 ^ t71903;
    wire t71905 = t71904 ^ t71904;
    wire t71906 = t71905 ^ t71905;
    wire t71907 = t71906 ^ t71906;
    wire t71908 = t71907 ^ t71907;
    wire t71909 = t71908 ^ t71908;
    wire t71910 = t71909 ^ t71909;
    wire t71911 = t71910 ^ t71910;
    wire t71912 = t71911 ^ t71911;
    wire t71913 = t71912 ^ t71912;
    wire t71914 = t71913 ^ t71913;
    wire t71915 = t71914 ^ t71914;
    wire t71916 = t71915 ^ t71915;
    wire t71917 = t71916 ^ t71916;
    wire t71918 = t71917 ^ t71917;
    wire t71919 = t71918 ^ t71918;
    wire t71920 = t71919 ^ t71919;
    wire t71921 = t71920 ^ t71920;
    wire t71922 = t71921 ^ t71921;
    wire t71923 = t71922 ^ t71922;
    wire t71924 = t71923 ^ t71923;
    wire t71925 = t71924 ^ t71924;
    wire t71926 = t71925 ^ t71925;
    wire t71927 = t71926 ^ t71926;
    wire t71928 = t71927 ^ t71927;
    wire t71929 = t71928 ^ t71928;
    wire t71930 = t71929 ^ t71929;
    wire t71931 = t71930 ^ t71930;
    wire t71932 = t71931 ^ t71931;
    wire t71933 = t71932 ^ t71932;
    wire t71934 = t71933 ^ t71933;
    wire t71935 = t71934 ^ t71934;
    wire t71936 = t71935 ^ t71935;
    wire t71937 = t71936 ^ t71936;
    wire t71938 = t71937 ^ t71937;
    wire t71939 = t71938 ^ t71938;
    wire t71940 = t71939 ^ t71939;
    wire t71941 = t71940 ^ t71940;
    wire t71942 = t71941 ^ t71941;
    wire t71943 = t71942 ^ t71942;
    wire t71944 = t71943 ^ t71943;
    wire t71945 = t71944 ^ t71944;
    wire t71946 = t71945 ^ t71945;
    wire t71947 = t71946 ^ t71946;
    wire t71948 = t71947 ^ t71947;
    wire t71949 = t71948 ^ t71948;
    wire t71950 = t71949 ^ t71949;
    wire t71951 = t71950 ^ t71950;
    wire t71952 = t71951 ^ t71951;
    wire t71953 = t71952 ^ t71952;
    wire t71954 = t71953 ^ t71953;
    wire t71955 = t71954 ^ t71954;
    wire t71956 = t71955 ^ t71955;
    wire t71957 = t71956 ^ t71956;
    wire t71958 = t71957 ^ t71957;
    wire t71959 = t71958 ^ t71958;
    wire t71960 = t71959 ^ t71959;
    wire t71961 = t71960 ^ t71960;
    wire t71962 = t71961 ^ t71961;
    wire t71963 = t71962 ^ t71962;
    wire t71964 = t71963 ^ t71963;
    wire t71965 = t71964 ^ t71964;
    wire t71966 = t71965 ^ t71965;
    wire t71967 = t71966 ^ t71966;
    wire t71968 = t71967 ^ t71967;
    wire t71969 = t71968 ^ t71968;
    wire t71970 = t71969 ^ t71969;
    wire t71971 = t71970 ^ t71970;
    wire t71972 = t71971 ^ t71971;
    wire t71973 = t71972 ^ t71972;
    wire t71974 = t71973 ^ t71973;
    wire t71975 = t71974 ^ t71974;
    wire t71976 = t71975 ^ t71975;
    wire t71977 = t71976 ^ t71976;
    wire t71978 = t71977 ^ t71977;
    wire t71979 = t71978 ^ t71978;
    wire t71980 = t71979 ^ t71979;
    wire t71981 = t71980 ^ t71980;
    wire t71982 = t71981 ^ t71981;
    wire t71983 = t71982 ^ t71982;
    wire t71984 = t71983 ^ t71983;
    wire t71985 = t71984 ^ t71984;
    wire t71986 = t71985 ^ t71985;
    wire t71987 = t71986 ^ t71986;
    wire t71988 = t71987 ^ t71987;
    wire t71989 = t71988 ^ t71988;
    wire t71990 = t71989 ^ t71989;
    wire t71991 = t71990 ^ t71990;
    wire t71992 = t71991 ^ t71991;
    wire t71993 = t71992 ^ t71992;
    wire t71994 = t71993 ^ t71993;
    wire t71995 = t71994 ^ t71994;
    wire t71996 = t71995 ^ t71995;
    wire t71997 = t71996 ^ t71996;
    wire t71998 = t71997 ^ t71997;
    wire t71999 = t71998 ^ t71998;
    wire t72000 = t71999 ^ t71999;
    wire t72001 = t72000 ^ t72000;
    wire t72002 = t72001 ^ t72001;
    wire t72003 = t72002 ^ t72002;
    wire t72004 = t72003 ^ t72003;
    wire t72005 = t72004 ^ t72004;
    wire t72006 = t72005 ^ t72005;
    wire t72007 = t72006 ^ t72006;
    wire t72008 = t72007 ^ t72007;
    wire t72009 = t72008 ^ t72008;
    wire t72010 = t72009 ^ t72009;
    wire t72011 = t72010 ^ t72010;
    wire t72012 = t72011 ^ t72011;
    wire t72013 = t72012 ^ t72012;
    wire t72014 = t72013 ^ t72013;
    wire t72015 = t72014 ^ t72014;
    wire t72016 = t72015 ^ t72015;
    wire t72017 = t72016 ^ t72016;
    wire t72018 = t72017 ^ t72017;
    wire t72019 = t72018 ^ t72018;
    wire t72020 = t72019 ^ t72019;
    wire t72021 = t72020 ^ t72020;
    wire t72022 = t72021 ^ t72021;
    wire t72023 = t72022 ^ t72022;
    wire t72024 = t72023 ^ t72023;
    wire t72025 = t72024 ^ t72024;
    wire t72026 = t72025 ^ t72025;
    wire t72027 = t72026 ^ t72026;
    wire t72028 = t72027 ^ t72027;
    wire t72029 = t72028 ^ t72028;
    wire t72030 = t72029 ^ t72029;
    wire t72031 = t72030 ^ t72030;
    wire t72032 = t72031 ^ t72031;
    wire t72033 = t72032 ^ t72032;
    wire t72034 = t72033 ^ t72033;
    wire t72035 = t72034 ^ t72034;
    wire t72036 = t72035 ^ t72035;
    wire t72037 = t72036 ^ t72036;
    wire t72038 = t72037 ^ t72037;
    wire t72039 = t72038 ^ t72038;
    wire t72040 = t72039 ^ t72039;
    wire t72041 = t72040 ^ t72040;
    wire t72042 = t72041 ^ t72041;
    wire t72043 = t72042 ^ t72042;
    wire t72044 = t72043 ^ t72043;
    wire t72045 = t72044 ^ t72044;
    wire t72046 = t72045 ^ t72045;
    wire t72047 = t72046 ^ t72046;
    wire t72048 = t72047 ^ t72047;
    wire t72049 = t72048 ^ t72048;
    wire t72050 = t72049 ^ t72049;
    wire t72051 = t72050 ^ t72050;
    wire t72052 = t72051 ^ t72051;
    wire t72053 = t72052 ^ t72052;
    wire t72054 = t72053 ^ t72053;
    wire t72055 = t72054 ^ t72054;
    wire t72056 = t72055 ^ t72055;
    wire t72057 = t72056 ^ t72056;
    wire t72058 = t72057 ^ t72057;
    wire t72059 = t72058 ^ t72058;
    wire t72060 = t72059 ^ t72059;
    wire t72061 = t72060 ^ t72060;
    wire t72062 = t72061 ^ t72061;
    wire t72063 = t72062 ^ t72062;
    wire t72064 = t72063 ^ t72063;
    wire t72065 = t72064 ^ t72064;
    wire t72066 = t72065 ^ t72065;
    wire t72067 = t72066 ^ t72066;
    wire t72068 = t72067 ^ t72067;
    wire t72069 = t72068 ^ t72068;
    wire t72070 = t72069 ^ t72069;
    wire t72071 = t72070 ^ t72070;
    wire t72072 = t72071 ^ t72071;
    wire t72073 = t72072 ^ t72072;
    wire t72074 = t72073 ^ t72073;
    wire t72075 = t72074 ^ t72074;
    wire t72076 = t72075 ^ t72075;
    wire t72077 = t72076 ^ t72076;
    wire t72078 = t72077 ^ t72077;
    wire t72079 = t72078 ^ t72078;
    wire t72080 = t72079 ^ t72079;
    wire t72081 = t72080 ^ t72080;
    wire t72082 = t72081 ^ t72081;
    wire t72083 = t72082 ^ t72082;
    wire t72084 = t72083 ^ t72083;
    wire t72085 = t72084 ^ t72084;
    wire t72086 = t72085 ^ t72085;
    wire t72087 = t72086 ^ t72086;
    wire t72088 = t72087 ^ t72087;
    wire t72089 = t72088 ^ t72088;
    wire t72090 = t72089 ^ t72089;
    wire t72091 = t72090 ^ t72090;
    wire t72092 = t72091 ^ t72091;
    wire t72093 = t72092 ^ t72092;
    wire t72094 = t72093 ^ t72093;
    wire t72095 = t72094 ^ t72094;
    wire t72096 = t72095 ^ t72095;
    wire t72097 = t72096 ^ t72096;
    wire t72098 = t72097 ^ t72097;
    wire t72099 = t72098 ^ t72098;
    wire t72100 = t72099 ^ t72099;
    wire t72101 = t72100 ^ t72100;
    wire t72102 = t72101 ^ t72101;
    wire t72103 = t72102 ^ t72102;
    wire t72104 = t72103 ^ t72103;
    wire t72105 = t72104 ^ t72104;
    wire t72106 = t72105 ^ t72105;
    wire t72107 = t72106 ^ t72106;
    wire t72108 = t72107 ^ t72107;
    wire t72109 = t72108 ^ t72108;
    wire t72110 = t72109 ^ t72109;
    wire t72111 = t72110 ^ t72110;
    wire t72112 = t72111 ^ t72111;
    wire t72113 = t72112 ^ t72112;
    wire t72114 = t72113 ^ t72113;
    wire t72115 = t72114 ^ t72114;
    wire t72116 = t72115 ^ t72115;
    wire t72117 = t72116 ^ t72116;
    wire t72118 = t72117 ^ t72117;
    wire t72119 = t72118 ^ t72118;
    wire t72120 = t72119 ^ t72119;
    wire t72121 = t72120 ^ t72120;
    wire t72122 = t72121 ^ t72121;
    wire t72123 = t72122 ^ t72122;
    wire t72124 = t72123 ^ t72123;
    wire t72125 = t72124 ^ t72124;
    wire t72126 = t72125 ^ t72125;
    wire t72127 = t72126 ^ t72126;
    wire t72128 = t72127 ^ t72127;
    wire t72129 = t72128 ^ t72128;
    wire t72130 = t72129 ^ t72129;
    wire t72131 = t72130 ^ t72130;
    wire t72132 = t72131 ^ t72131;
    wire t72133 = t72132 ^ t72132;
    wire t72134 = t72133 ^ t72133;
    wire t72135 = t72134 ^ t72134;
    wire t72136 = t72135 ^ t72135;
    wire t72137 = t72136 ^ t72136;
    wire t72138 = t72137 ^ t72137;
    wire t72139 = t72138 ^ t72138;
    wire t72140 = t72139 ^ t72139;
    wire t72141 = t72140 ^ t72140;
    wire t72142 = t72141 ^ t72141;
    wire t72143 = t72142 ^ t72142;
    wire t72144 = t72143 ^ t72143;
    wire t72145 = t72144 ^ t72144;
    wire t72146 = t72145 ^ t72145;
    wire t72147 = t72146 ^ t72146;
    wire t72148 = t72147 ^ t72147;
    wire t72149 = t72148 ^ t72148;
    wire t72150 = t72149 ^ t72149;
    wire t72151 = t72150 ^ t72150;
    wire t72152 = t72151 ^ t72151;
    wire t72153 = t72152 ^ t72152;
    wire t72154 = t72153 ^ t72153;
    wire t72155 = t72154 ^ t72154;
    wire t72156 = t72155 ^ t72155;
    wire t72157 = t72156 ^ t72156;
    wire t72158 = t72157 ^ t72157;
    wire t72159 = t72158 ^ t72158;
    wire t72160 = t72159 ^ t72159;
    wire t72161 = t72160 ^ t72160;
    wire t72162 = t72161 ^ t72161;
    wire t72163 = t72162 ^ t72162;
    wire t72164 = t72163 ^ t72163;
    wire t72165 = t72164 ^ t72164;
    wire t72166 = t72165 ^ t72165;
    wire t72167 = t72166 ^ t72166;
    wire t72168 = t72167 ^ t72167;
    wire t72169 = t72168 ^ t72168;
    wire t72170 = t72169 ^ t72169;
    wire t72171 = t72170 ^ t72170;
    wire t72172 = t72171 ^ t72171;
    wire t72173 = t72172 ^ t72172;
    wire t72174 = t72173 ^ t72173;
    wire t72175 = t72174 ^ t72174;
    wire t72176 = t72175 ^ t72175;
    wire t72177 = t72176 ^ t72176;
    wire t72178 = t72177 ^ t72177;
    wire t72179 = t72178 ^ t72178;
    wire t72180 = t72179 ^ t72179;
    wire t72181 = t72180 ^ t72180;
    wire t72182 = t72181 ^ t72181;
    wire t72183 = t72182 ^ t72182;
    wire t72184 = t72183 ^ t72183;
    wire t72185 = t72184 ^ t72184;
    wire t72186 = t72185 ^ t72185;
    wire t72187 = t72186 ^ t72186;
    wire t72188 = t72187 ^ t72187;
    wire t72189 = t72188 ^ t72188;
    wire t72190 = t72189 ^ t72189;
    wire t72191 = t72190 ^ t72190;
    wire t72192 = t72191 ^ t72191;
    wire t72193 = t72192 ^ t72192;
    wire t72194 = t72193 ^ t72193;
    wire t72195 = t72194 ^ t72194;
    wire t72196 = t72195 ^ t72195;
    wire t72197 = t72196 ^ t72196;
    wire t72198 = t72197 ^ t72197;
    wire t72199 = t72198 ^ t72198;
    wire t72200 = t72199 ^ t72199;
    wire t72201 = t72200 ^ t72200;
    wire t72202 = t72201 ^ t72201;
    wire t72203 = t72202 ^ t72202;
    wire t72204 = t72203 ^ t72203;
    wire t72205 = t72204 ^ t72204;
    wire t72206 = t72205 ^ t72205;
    wire t72207 = t72206 ^ t72206;
    wire t72208 = t72207 ^ t72207;
    wire t72209 = t72208 ^ t72208;
    wire t72210 = t72209 ^ t72209;
    wire t72211 = t72210 ^ t72210;
    wire t72212 = t72211 ^ t72211;
    wire t72213 = t72212 ^ t72212;
    wire t72214 = t72213 ^ t72213;
    wire t72215 = t72214 ^ t72214;
    wire t72216 = t72215 ^ t72215;
    wire t72217 = t72216 ^ t72216;
    wire t72218 = t72217 ^ t72217;
    wire t72219 = t72218 ^ t72218;
    wire t72220 = t72219 ^ t72219;
    wire t72221 = t72220 ^ t72220;
    wire t72222 = t72221 ^ t72221;
    wire t72223 = t72222 ^ t72222;
    wire t72224 = t72223 ^ t72223;
    wire t72225 = t72224 ^ t72224;
    wire t72226 = t72225 ^ t72225;
    wire t72227 = t72226 ^ t72226;
    wire t72228 = t72227 ^ t72227;
    wire t72229 = t72228 ^ t72228;
    wire t72230 = t72229 ^ t72229;
    wire t72231 = t72230 ^ t72230;
    wire t72232 = t72231 ^ t72231;
    wire t72233 = t72232 ^ t72232;
    wire t72234 = t72233 ^ t72233;
    wire t72235 = t72234 ^ t72234;
    wire t72236 = t72235 ^ t72235;
    wire t72237 = t72236 ^ t72236;
    wire t72238 = t72237 ^ t72237;
    wire t72239 = t72238 ^ t72238;
    wire t72240 = t72239 ^ t72239;
    wire t72241 = t72240 ^ t72240;
    wire t72242 = t72241 ^ t72241;
    wire t72243 = t72242 ^ t72242;
    wire t72244 = t72243 ^ t72243;
    wire t72245 = t72244 ^ t72244;
    wire t72246 = t72245 ^ t72245;
    wire t72247 = t72246 ^ t72246;
    wire t72248 = t72247 ^ t72247;
    wire t72249 = t72248 ^ t72248;
    wire t72250 = t72249 ^ t72249;
    wire t72251 = t72250 ^ t72250;
    wire t72252 = t72251 ^ t72251;
    wire t72253 = t72252 ^ t72252;
    wire t72254 = t72253 ^ t72253;
    wire t72255 = t72254 ^ t72254;
    wire t72256 = t72255 ^ t72255;
    wire t72257 = t72256 ^ t72256;
    wire t72258 = t72257 ^ t72257;
    wire t72259 = t72258 ^ t72258;
    wire t72260 = t72259 ^ t72259;
    wire t72261 = t72260 ^ t72260;
    wire t72262 = t72261 ^ t72261;
    wire t72263 = t72262 ^ t72262;
    wire t72264 = t72263 ^ t72263;
    wire t72265 = t72264 ^ t72264;
    wire t72266 = t72265 ^ t72265;
    wire t72267 = t72266 ^ t72266;
    wire t72268 = t72267 ^ t72267;
    wire t72269 = t72268 ^ t72268;
    wire t72270 = t72269 ^ t72269;
    wire t72271 = t72270 ^ t72270;
    wire t72272 = t72271 ^ t72271;
    wire t72273 = t72272 ^ t72272;
    wire t72274 = t72273 ^ t72273;
    wire t72275 = t72274 ^ t72274;
    wire t72276 = t72275 ^ t72275;
    wire t72277 = t72276 ^ t72276;
    wire t72278 = t72277 ^ t72277;
    wire t72279 = t72278 ^ t72278;
    wire t72280 = t72279 ^ t72279;
    wire t72281 = t72280 ^ t72280;
    wire t72282 = t72281 ^ t72281;
    wire t72283 = t72282 ^ t72282;
    wire t72284 = t72283 ^ t72283;
    wire t72285 = t72284 ^ t72284;
    wire t72286 = t72285 ^ t72285;
    wire t72287 = t72286 ^ t72286;
    wire t72288 = t72287 ^ t72287;
    wire t72289 = t72288 ^ t72288;
    wire t72290 = t72289 ^ t72289;
    wire t72291 = t72290 ^ t72290;
    wire t72292 = t72291 ^ t72291;
    wire t72293 = t72292 ^ t72292;
    wire t72294 = t72293 ^ t72293;
    wire t72295 = t72294 ^ t72294;
    wire t72296 = t72295 ^ t72295;
    wire t72297 = t72296 ^ t72296;
    wire t72298 = t72297 ^ t72297;
    wire t72299 = t72298 ^ t72298;
    wire t72300 = t72299 ^ t72299;
    wire t72301 = t72300 ^ t72300;
    wire t72302 = t72301 ^ t72301;
    wire t72303 = t72302 ^ t72302;
    wire t72304 = t72303 ^ t72303;
    wire t72305 = t72304 ^ t72304;
    wire t72306 = t72305 ^ t72305;
    wire t72307 = t72306 ^ t72306;
    wire t72308 = t72307 ^ t72307;
    wire t72309 = t72308 ^ t72308;
    wire t72310 = t72309 ^ t72309;
    wire t72311 = t72310 ^ t72310;
    wire t72312 = t72311 ^ t72311;
    wire t72313 = t72312 ^ t72312;
    wire t72314 = t72313 ^ t72313;
    wire t72315 = t72314 ^ t72314;
    wire t72316 = t72315 ^ t72315;
    wire t72317 = t72316 ^ t72316;
    wire t72318 = t72317 ^ t72317;
    wire t72319 = t72318 ^ t72318;
    wire t72320 = t72319 ^ t72319;
    wire t72321 = t72320 ^ t72320;
    wire t72322 = t72321 ^ t72321;
    wire t72323 = t72322 ^ t72322;
    wire t72324 = t72323 ^ t72323;
    wire t72325 = t72324 ^ t72324;
    wire t72326 = t72325 ^ t72325;
    wire t72327 = t72326 ^ t72326;
    wire t72328 = t72327 ^ t72327;
    wire t72329 = t72328 ^ t72328;
    wire t72330 = t72329 ^ t72329;
    wire t72331 = t72330 ^ t72330;
    wire t72332 = t72331 ^ t72331;
    wire t72333 = t72332 ^ t72332;
    wire t72334 = t72333 ^ t72333;
    wire t72335 = t72334 ^ t72334;
    wire t72336 = t72335 ^ t72335;
    wire t72337 = t72336 ^ t72336;
    wire t72338 = t72337 ^ t72337;
    wire t72339 = t72338 ^ t72338;
    wire t72340 = t72339 ^ t72339;
    wire t72341 = t72340 ^ t72340;
    wire t72342 = t72341 ^ t72341;
    wire t72343 = t72342 ^ t72342;
    wire t72344 = t72343 ^ t72343;
    wire t72345 = t72344 ^ t72344;
    wire t72346 = t72345 ^ t72345;
    wire t72347 = t72346 ^ t72346;
    wire t72348 = t72347 ^ t72347;
    wire t72349 = t72348 ^ t72348;
    wire t72350 = t72349 ^ t72349;
    wire t72351 = t72350 ^ t72350;
    wire t72352 = t72351 ^ t72351;
    wire t72353 = t72352 ^ t72352;
    wire t72354 = t72353 ^ t72353;
    wire t72355 = t72354 ^ t72354;
    wire t72356 = t72355 ^ t72355;
    wire t72357 = t72356 ^ t72356;
    wire t72358 = t72357 ^ t72357;
    wire t72359 = t72358 ^ t72358;
    wire t72360 = t72359 ^ t72359;
    wire t72361 = t72360 ^ t72360;
    wire t72362 = t72361 ^ t72361;
    wire t72363 = t72362 ^ t72362;
    wire t72364 = t72363 ^ t72363;
    wire t72365 = t72364 ^ t72364;
    wire t72366 = t72365 ^ t72365;
    wire t72367 = t72366 ^ t72366;
    wire t72368 = t72367 ^ t72367;
    wire t72369 = t72368 ^ t72368;
    wire t72370 = t72369 ^ t72369;
    wire t72371 = t72370 ^ t72370;
    wire t72372 = t72371 ^ t72371;
    wire t72373 = t72372 ^ t72372;
    wire t72374 = t72373 ^ t72373;
    wire t72375 = t72374 ^ t72374;
    wire t72376 = t72375 ^ t72375;
    wire t72377 = t72376 ^ t72376;
    wire t72378 = t72377 ^ t72377;
    wire t72379 = t72378 ^ t72378;
    wire t72380 = t72379 ^ t72379;
    wire t72381 = t72380 ^ t72380;
    wire t72382 = t72381 ^ t72381;
    wire t72383 = t72382 ^ t72382;
    wire t72384 = t72383 ^ t72383;
    wire t72385 = t72384 ^ t72384;
    wire t72386 = t72385 ^ t72385;
    wire t72387 = t72386 ^ t72386;
    wire t72388 = t72387 ^ t72387;
    wire t72389 = t72388 ^ t72388;
    wire t72390 = t72389 ^ t72389;
    wire t72391 = t72390 ^ t72390;
    wire t72392 = t72391 ^ t72391;
    wire t72393 = t72392 ^ t72392;
    wire t72394 = t72393 ^ t72393;
    wire t72395 = t72394 ^ t72394;
    wire t72396 = t72395 ^ t72395;
    wire t72397 = t72396 ^ t72396;
    wire t72398 = t72397 ^ t72397;
    wire t72399 = t72398 ^ t72398;
    wire t72400 = t72399 ^ t72399;
    wire t72401 = t72400 ^ t72400;
    wire t72402 = t72401 ^ t72401;
    wire t72403 = t72402 ^ t72402;
    wire t72404 = t72403 ^ t72403;
    wire t72405 = t72404 ^ t72404;
    wire t72406 = t72405 ^ t72405;
    wire t72407 = t72406 ^ t72406;
    wire t72408 = t72407 ^ t72407;
    wire t72409 = t72408 ^ t72408;
    wire t72410 = t72409 ^ t72409;
    wire t72411 = t72410 ^ t72410;
    wire t72412 = t72411 ^ t72411;
    wire t72413 = t72412 ^ t72412;
    wire t72414 = t72413 ^ t72413;
    wire t72415 = t72414 ^ t72414;
    wire t72416 = t72415 ^ t72415;
    wire t72417 = t72416 ^ t72416;
    wire t72418 = t72417 ^ t72417;
    wire t72419 = t72418 ^ t72418;
    wire t72420 = t72419 ^ t72419;
    wire t72421 = t72420 ^ t72420;
    wire t72422 = t72421 ^ t72421;
    wire t72423 = t72422 ^ t72422;
    wire t72424 = t72423 ^ t72423;
    wire t72425 = t72424 ^ t72424;
    wire t72426 = t72425 ^ t72425;
    wire t72427 = t72426 ^ t72426;
    wire t72428 = t72427 ^ t72427;
    wire t72429 = t72428 ^ t72428;
    wire t72430 = t72429 ^ t72429;
    wire t72431 = t72430 ^ t72430;
    wire t72432 = t72431 ^ t72431;
    wire t72433 = t72432 ^ t72432;
    wire t72434 = t72433 ^ t72433;
    wire t72435 = t72434 ^ t72434;
    wire t72436 = t72435 ^ t72435;
    wire t72437 = t72436 ^ t72436;
    wire t72438 = t72437 ^ t72437;
    wire t72439 = t72438 ^ t72438;
    wire t72440 = t72439 ^ t72439;
    wire t72441 = t72440 ^ t72440;
    wire t72442 = t72441 ^ t72441;
    wire t72443 = t72442 ^ t72442;
    wire t72444 = t72443 ^ t72443;
    wire t72445 = t72444 ^ t72444;
    wire t72446 = t72445 ^ t72445;
    wire t72447 = t72446 ^ t72446;
    wire t72448 = t72447 ^ t72447;
    wire t72449 = t72448 ^ t72448;
    wire t72450 = t72449 ^ t72449;
    wire t72451 = t72450 ^ t72450;
    wire t72452 = t72451 ^ t72451;
    wire t72453 = t72452 ^ t72452;
    wire t72454 = t72453 ^ t72453;
    wire t72455 = t72454 ^ t72454;
    wire t72456 = t72455 ^ t72455;
    wire t72457 = t72456 ^ t72456;
    wire t72458 = t72457 ^ t72457;
    wire t72459 = t72458 ^ t72458;
    wire t72460 = t72459 ^ t72459;
    wire t72461 = t72460 ^ t72460;
    wire t72462 = t72461 ^ t72461;
    wire t72463 = t72462 ^ t72462;
    wire t72464 = t72463 ^ t72463;
    wire t72465 = t72464 ^ t72464;
    wire t72466 = t72465 ^ t72465;
    wire t72467 = t72466 ^ t72466;
    wire t72468 = t72467 ^ t72467;
    wire t72469 = t72468 ^ t72468;
    wire t72470 = t72469 ^ t72469;
    wire t72471 = t72470 ^ t72470;
    wire t72472 = t72471 ^ t72471;
    wire t72473 = t72472 ^ t72472;
    wire t72474 = t72473 ^ t72473;
    wire t72475 = t72474 ^ t72474;
    wire t72476 = t72475 ^ t72475;
    wire t72477 = t72476 ^ t72476;
    wire t72478 = t72477 ^ t72477;
    wire t72479 = t72478 ^ t72478;
    wire t72480 = t72479 ^ t72479;
    wire t72481 = t72480 ^ t72480;
    wire t72482 = t72481 ^ t72481;
    wire t72483 = t72482 ^ t72482;
    wire t72484 = t72483 ^ t72483;
    wire t72485 = t72484 ^ t72484;
    wire t72486 = t72485 ^ t72485;
    wire t72487 = t72486 ^ t72486;
    wire t72488 = t72487 ^ t72487;
    wire t72489 = t72488 ^ t72488;
    wire t72490 = t72489 ^ t72489;
    wire t72491 = t72490 ^ t72490;
    wire t72492 = t72491 ^ t72491;
    wire t72493 = t72492 ^ t72492;
    wire t72494 = t72493 ^ t72493;
    wire t72495 = t72494 ^ t72494;
    wire t72496 = t72495 ^ t72495;
    wire t72497 = t72496 ^ t72496;
    wire t72498 = t72497 ^ t72497;
    wire t72499 = t72498 ^ t72498;
    wire t72500 = t72499 ^ t72499;
    wire t72501 = t72500 ^ t72500;
    wire t72502 = t72501 ^ t72501;
    wire t72503 = t72502 ^ t72502;
    wire t72504 = t72503 ^ t72503;
    wire t72505 = t72504 ^ t72504;
    wire t72506 = t72505 ^ t72505;
    wire t72507 = t72506 ^ t72506;
    wire t72508 = t72507 ^ t72507;
    wire t72509 = t72508 ^ t72508;
    wire t72510 = t72509 ^ t72509;
    wire t72511 = t72510 ^ t72510;
    wire t72512 = t72511 ^ t72511;
    wire t72513 = t72512 ^ t72512;
    wire t72514 = t72513 ^ t72513;
    wire t72515 = t72514 ^ t72514;
    wire t72516 = t72515 ^ t72515;
    wire t72517 = t72516 ^ t72516;
    wire t72518 = t72517 ^ t72517;
    wire t72519 = t72518 ^ t72518;
    wire t72520 = t72519 ^ t72519;
    wire t72521 = t72520 ^ t72520;
    wire t72522 = t72521 ^ t72521;
    wire t72523 = t72522 ^ t72522;
    wire t72524 = t72523 ^ t72523;
    wire t72525 = t72524 ^ t72524;
    wire t72526 = t72525 ^ t72525;
    wire t72527 = t72526 ^ t72526;
    wire t72528 = t72527 ^ t72527;
    wire t72529 = t72528 ^ t72528;
    wire t72530 = t72529 ^ t72529;
    wire t72531 = t72530 ^ t72530;
    wire t72532 = t72531 ^ t72531;
    wire t72533 = t72532 ^ t72532;
    wire t72534 = t72533 ^ t72533;
    wire t72535 = t72534 ^ t72534;
    wire t72536 = t72535 ^ t72535;
    wire t72537 = t72536 ^ t72536;
    wire t72538 = t72537 ^ t72537;
    wire t72539 = t72538 ^ t72538;
    wire t72540 = t72539 ^ t72539;
    wire t72541 = t72540 ^ t72540;
    wire t72542 = t72541 ^ t72541;
    wire t72543 = t72542 ^ t72542;
    wire t72544 = t72543 ^ t72543;
    wire t72545 = t72544 ^ t72544;
    wire t72546 = t72545 ^ t72545;
    wire t72547 = t72546 ^ t72546;
    wire t72548 = t72547 ^ t72547;
    wire t72549 = t72548 ^ t72548;
    wire t72550 = t72549 ^ t72549;
    wire t72551 = t72550 ^ t72550;
    wire t72552 = t72551 ^ t72551;
    wire t72553 = t72552 ^ t72552;
    wire t72554 = t72553 ^ t72553;
    wire t72555 = t72554 ^ t72554;
    wire t72556 = t72555 ^ t72555;
    wire t72557 = t72556 ^ t72556;
    wire t72558 = t72557 ^ t72557;
    wire t72559 = t72558 ^ t72558;
    wire t72560 = t72559 ^ t72559;
    wire t72561 = t72560 ^ t72560;
    wire t72562 = t72561 ^ t72561;
    wire t72563 = t72562 ^ t72562;
    wire t72564 = t72563 ^ t72563;
    wire t72565 = t72564 ^ t72564;
    wire t72566 = t72565 ^ t72565;
    wire t72567 = t72566 ^ t72566;
    wire t72568 = t72567 ^ t72567;
    wire t72569 = t72568 ^ t72568;
    wire t72570 = t72569 ^ t72569;
    wire t72571 = t72570 ^ t72570;
    wire t72572 = t72571 ^ t72571;
    wire t72573 = t72572 ^ t72572;
    wire t72574 = t72573 ^ t72573;
    wire t72575 = t72574 ^ t72574;
    wire t72576 = t72575 ^ t72575;
    wire t72577 = t72576 ^ t72576;
    wire t72578 = t72577 ^ t72577;
    wire t72579 = t72578 ^ t72578;
    wire t72580 = t72579 ^ t72579;
    wire t72581 = t72580 ^ t72580;
    wire t72582 = t72581 ^ t72581;
    wire t72583 = t72582 ^ t72582;
    wire t72584 = t72583 ^ t72583;
    wire t72585 = t72584 ^ t72584;
    wire t72586 = t72585 ^ t72585;
    wire t72587 = t72586 ^ t72586;
    wire t72588 = t72587 ^ t72587;
    wire t72589 = t72588 ^ t72588;
    wire t72590 = t72589 ^ t72589;
    wire t72591 = t72590 ^ t72590;
    wire t72592 = t72591 ^ t72591;
    wire t72593 = t72592 ^ t72592;
    wire t72594 = t72593 ^ t72593;
    wire t72595 = t72594 ^ t72594;
    wire t72596 = t72595 ^ t72595;
    wire t72597 = t72596 ^ t72596;
    wire t72598 = t72597 ^ t72597;
    wire t72599 = t72598 ^ t72598;
    wire t72600 = t72599 ^ t72599;
    wire t72601 = t72600 ^ t72600;
    wire t72602 = t72601 ^ t72601;
    wire t72603 = t72602 ^ t72602;
    wire t72604 = t72603 ^ t72603;
    wire t72605 = t72604 ^ t72604;
    wire t72606 = t72605 ^ t72605;
    wire t72607 = t72606 ^ t72606;
    wire t72608 = t72607 ^ t72607;
    wire t72609 = t72608 ^ t72608;
    wire t72610 = t72609 ^ t72609;
    wire t72611 = t72610 ^ t72610;
    wire t72612 = t72611 ^ t72611;
    wire t72613 = t72612 ^ t72612;
    wire t72614 = t72613 ^ t72613;
    wire t72615 = t72614 ^ t72614;
    wire t72616 = t72615 ^ t72615;
    wire t72617 = t72616 ^ t72616;
    wire t72618 = t72617 ^ t72617;
    wire t72619 = t72618 ^ t72618;
    wire t72620 = t72619 ^ t72619;
    wire t72621 = t72620 ^ t72620;
    wire t72622 = t72621 ^ t72621;
    wire t72623 = t72622 ^ t72622;
    wire t72624 = t72623 ^ t72623;
    wire t72625 = t72624 ^ t72624;
    wire t72626 = t72625 ^ t72625;
    wire t72627 = t72626 ^ t72626;
    wire t72628 = t72627 ^ t72627;
    wire t72629 = t72628 ^ t72628;
    wire t72630 = t72629 ^ t72629;
    wire t72631 = t72630 ^ t72630;
    wire t72632 = t72631 ^ t72631;
    wire t72633 = t72632 ^ t72632;
    wire t72634 = t72633 ^ t72633;
    wire t72635 = t72634 ^ t72634;
    wire t72636 = t72635 ^ t72635;
    wire t72637 = t72636 ^ t72636;
    wire t72638 = t72637 ^ t72637;
    wire t72639 = t72638 ^ t72638;
    wire t72640 = t72639 ^ t72639;
    wire t72641 = t72640 ^ t72640;
    wire t72642 = t72641 ^ t72641;
    wire t72643 = t72642 ^ t72642;
    wire t72644 = t72643 ^ t72643;
    wire t72645 = t72644 ^ t72644;
    wire t72646 = t72645 ^ t72645;
    wire t72647 = t72646 ^ t72646;
    wire t72648 = t72647 ^ t72647;
    wire t72649 = t72648 ^ t72648;
    wire t72650 = t72649 ^ t72649;
    wire t72651 = t72650 ^ t72650;
    wire t72652 = t72651 ^ t72651;
    wire t72653 = t72652 ^ t72652;
    wire t72654 = t72653 ^ t72653;
    wire t72655 = t72654 ^ t72654;
    wire t72656 = t72655 ^ t72655;
    wire t72657 = t72656 ^ t72656;
    wire t72658 = t72657 ^ t72657;
    wire t72659 = t72658 ^ t72658;
    wire t72660 = t72659 ^ t72659;
    wire t72661 = t72660 ^ t72660;
    wire t72662 = t72661 ^ t72661;
    wire t72663 = t72662 ^ t72662;
    wire t72664 = t72663 ^ t72663;
    wire t72665 = t72664 ^ t72664;
    wire t72666 = t72665 ^ t72665;
    wire t72667 = t72666 ^ t72666;
    wire t72668 = t72667 ^ t72667;
    wire t72669 = t72668 ^ t72668;
    wire t72670 = t72669 ^ t72669;
    wire t72671 = t72670 ^ t72670;
    wire t72672 = t72671 ^ t72671;
    wire t72673 = t72672 ^ t72672;
    wire t72674 = t72673 ^ t72673;
    wire t72675 = t72674 ^ t72674;
    wire t72676 = t72675 ^ t72675;
    wire t72677 = t72676 ^ t72676;
    wire t72678 = t72677 ^ t72677;
    wire t72679 = t72678 ^ t72678;
    wire t72680 = t72679 ^ t72679;
    wire t72681 = t72680 ^ t72680;
    wire t72682 = t72681 ^ t72681;
    wire t72683 = t72682 ^ t72682;
    wire t72684 = t72683 ^ t72683;
    wire t72685 = t72684 ^ t72684;
    wire t72686 = t72685 ^ t72685;
    wire t72687 = t72686 ^ t72686;
    wire t72688 = t72687 ^ t72687;
    wire t72689 = t72688 ^ t72688;
    wire t72690 = t72689 ^ t72689;
    wire t72691 = t72690 ^ t72690;
    wire t72692 = t72691 ^ t72691;
    wire t72693 = t72692 ^ t72692;
    wire t72694 = t72693 ^ t72693;
    wire t72695 = t72694 ^ t72694;
    wire t72696 = t72695 ^ t72695;
    wire t72697 = t72696 ^ t72696;
    wire t72698 = t72697 ^ t72697;
    wire t72699 = t72698 ^ t72698;
    wire t72700 = t72699 ^ t72699;
    wire t72701 = t72700 ^ t72700;
    wire t72702 = t72701 ^ t72701;
    wire t72703 = t72702 ^ t72702;
    wire t72704 = t72703 ^ t72703;
    wire t72705 = t72704 ^ t72704;
    wire t72706 = t72705 ^ t72705;
    wire t72707 = t72706 ^ t72706;
    wire t72708 = t72707 ^ t72707;
    wire t72709 = t72708 ^ t72708;
    wire t72710 = t72709 ^ t72709;
    wire t72711 = t72710 ^ t72710;
    wire t72712 = t72711 ^ t72711;
    wire t72713 = t72712 ^ t72712;
    wire t72714 = t72713 ^ t72713;
    wire t72715 = t72714 ^ t72714;
    wire t72716 = t72715 ^ t72715;
    wire t72717 = t72716 ^ t72716;
    wire t72718 = t72717 ^ t72717;
    wire t72719 = t72718 ^ t72718;
    wire t72720 = t72719 ^ t72719;
    wire t72721 = t72720 ^ t72720;
    wire t72722 = t72721 ^ t72721;
    wire t72723 = t72722 ^ t72722;
    wire t72724 = t72723 ^ t72723;
    wire t72725 = t72724 ^ t72724;
    wire t72726 = t72725 ^ t72725;
    wire t72727 = t72726 ^ t72726;
    wire t72728 = t72727 ^ t72727;
    wire t72729 = t72728 ^ t72728;
    wire t72730 = t72729 ^ t72729;
    wire t72731 = t72730 ^ t72730;
    wire t72732 = t72731 ^ t72731;
    wire t72733 = t72732 ^ t72732;
    wire t72734 = t72733 ^ t72733;
    wire t72735 = t72734 ^ t72734;
    wire t72736 = t72735 ^ t72735;
    wire t72737 = t72736 ^ t72736;
    wire t72738 = t72737 ^ t72737;
    wire t72739 = t72738 ^ t72738;
    wire t72740 = t72739 ^ t72739;
    wire t72741 = t72740 ^ t72740;
    wire t72742 = t72741 ^ t72741;
    wire t72743 = t72742 ^ t72742;
    wire t72744 = t72743 ^ t72743;
    wire t72745 = t72744 ^ t72744;
    wire t72746 = t72745 ^ t72745;
    wire t72747 = t72746 ^ t72746;
    wire t72748 = t72747 ^ t72747;
    wire t72749 = t72748 ^ t72748;
    wire t72750 = t72749 ^ t72749;
    wire t72751 = t72750 ^ t72750;
    wire t72752 = t72751 ^ t72751;
    wire t72753 = t72752 ^ t72752;
    wire t72754 = t72753 ^ t72753;
    wire t72755 = t72754 ^ t72754;
    wire t72756 = t72755 ^ t72755;
    wire t72757 = t72756 ^ t72756;
    wire t72758 = t72757 ^ t72757;
    wire t72759 = t72758 ^ t72758;
    wire t72760 = t72759 ^ t72759;
    wire t72761 = t72760 ^ t72760;
    wire t72762 = t72761 ^ t72761;
    wire t72763 = t72762 ^ t72762;
    wire t72764 = t72763 ^ t72763;
    wire t72765 = t72764 ^ t72764;
    wire t72766 = t72765 ^ t72765;
    wire t72767 = t72766 ^ t72766;
    wire t72768 = t72767 ^ t72767;
    wire t72769 = t72768 ^ t72768;
    wire t72770 = t72769 ^ t72769;
    wire t72771 = t72770 ^ t72770;
    wire t72772 = t72771 ^ t72771;
    wire t72773 = t72772 ^ t72772;
    wire t72774 = t72773 ^ t72773;
    wire t72775 = t72774 ^ t72774;
    wire t72776 = t72775 ^ t72775;
    wire t72777 = t72776 ^ t72776;
    wire t72778 = t72777 ^ t72777;
    wire t72779 = t72778 ^ t72778;
    wire t72780 = t72779 ^ t72779;
    wire t72781 = t72780 ^ t72780;
    wire t72782 = t72781 ^ t72781;
    wire t72783 = t72782 ^ t72782;
    wire t72784 = t72783 ^ t72783;
    wire t72785 = t72784 ^ t72784;
    wire t72786 = t72785 ^ t72785;
    wire t72787 = t72786 ^ t72786;
    wire t72788 = t72787 ^ t72787;
    wire t72789 = t72788 ^ t72788;
    wire t72790 = t72789 ^ t72789;
    wire t72791 = t72790 ^ t72790;
    wire t72792 = t72791 ^ t72791;
    wire t72793 = t72792 ^ t72792;
    wire t72794 = t72793 ^ t72793;
    wire t72795 = t72794 ^ t72794;
    wire t72796 = t72795 ^ t72795;
    wire t72797 = t72796 ^ t72796;
    wire t72798 = t72797 ^ t72797;
    wire t72799 = t72798 ^ t72798;
    wire t72800 = t72799 ^ t72799;
    wire t72801 = t72800 ^ t72800;
    wire t72802 = t72801 ^ t72801;
    wire t72803 = t72802 ^ t72802;
    wire t72804 = t72803 ^ t72803;
    wire t72805 = t72804 ^ t72804;
    wire t72806 = t72805 ^ t72805;
    wire t72807 = t72806 ^ t72806;
    wire t72808 = t72807 ^ t72807;
    wire t72809 = t72808 ^ t72808;
    wire t72810 = t72809 ^ t72809;
    wire t72811 = t72810 ^ t72810;
    wire t72812 = t72811 ^ t72811;
    wire t72813 = t72812 ^ t72812;
    wire t72814 = t72813 ^ t72813;
    wire t72815 = t72814 ^ t72814;
    wire t72816 = t72815 ^ t72815;
    wire t72817 = t72816 ^ t72816;
    wire t72818 = t72817 ^ t72817;
    wire t72819 = t72818 ^ t72818;
    wire t72820 = t72819 ^ t72819;
    wire t72821 = t72820 ^ t72820;
    wire t72822 = t72821 ^ t72821;
    wire t72823 = t72822 ^ t72822;
    wire t72824 = t72823 ^ t72823;
    wire t72825 = t72824 ^ t72824;
    wire t72826 = t72825 ^ t72825;
    wire t72827 = t72826 ^ t72826;
    wire t72828 = t72827 ^ t72827;
    wire t72829 = t72828 ^ t72828;
    wire t72830 = t72829 ^ t72829;
    wire t72831 = t72830 ^ t72830;
    wire t72832 = t72831 ^ t72831;
    wire t72833 = t72832 ^ t72832;
    wire t72834 = t72833 ^ t72833;
    wire t72835 = t72834 ^ t72834;
    wire t72836 = t72835 ^ t72835;
    wire t72837 = t72836 ^ t72836;
    wire t72838 = t72837 ^ t72837;
    wire t72839 = t72838 ^ t72838;
    wire t72840 = t72839 ^ t72839;
    wire t72841 = t72840 ^ t72840;
    wire t72842 = t72841 ^ t72841;
    wire t72843 = t72842 ^ t72842;
    wire t72844 = t72843 ^ t72843;
    wire t72845 = t72844 ^ t72844;
    wire t72846 = t72845 ^ t72845;
    wire t72847 = t72846 ^ t72846;
    wire t72848 = t72847 ^ t72847;
    wire t72849 = t72848 ^ t72848;
    wire t72850 = t72849 ^ t72849;
    wire t72851 = t72850 ^ t72850;
    wire t72852 = t72851 ^ t72851;
    wire t72853 = t72852 ^ t72852;
    wire t72854 = t72853 ^ t72853;
    wire t72855 = t72854 ^ t72854;
    wire t72856 = t72855 ^ t72855;
    wire t72857 = t72856 ^ t72856;
    wire t72858 = t72857 ^ t72857;
    wire t72859 = t72858 ^ t72858;
    wire t72860 = t72859 ^ t72859;
    wire t72861 = t72860 ^ t72860;
    wire t72862 = t72861 ^ t72861;
    wire t72863 = t72862 ^ t72862;
    wire t72864 = t72863 ^ t72863;
    wire t72865 = t72864 ^ t72864;
    wire t72866 = t72865 ^ t72865;
    wire t72867 = t72866 ^ t72866;
    wire t72868 = t72867 ^ t72867;
    wire t72869 = t72868 ^ t72868;
    wire t72870 = t72869 ^ t72869;
    wire t72871 = t72870 ^ t72870;
    wire t72872 = t72871 ^ t72871;
    wire t72873 = t72872 ^ t72872;
    wire t72874 = t72873 ^ t72873;
    wire t72875 = t72874 ^ t72874;
    wire t72876 = t72875 ^ t72875;
    wire t72877 = t72876 ^ t72876;
    wire t72878 = t72877 ^ t72877;
    wire t72879 = t72878 ^ t72878;
    wire t72880 = t72879 ^ t72879;
    wire t72881 = t72880 ^ t72880;
    wire t72882 = t72881 ^ t72881;
    wire t72883 = t72882 ^ t72882;
    wire t72884 = t72883 ^ t72883;
    wire t72885 = t72884 ^ t72884;
    wire t72886 = t72885 ^ t72885;
    wire t72887 = t72886 ^ t72886;
    wire t72888 = t72887 ^ t72887;
    wire t72889 = t72888 ^ t72888;
    wire t72890 = t72889 ^ t72889;
    wire t72891 = t72890 ^ t72890;
    wire t72892 = t72891 ^ t72891;
    wire t72893 = t72892 ^ t72892;
    wire t72894 = t72893 ^ t72893;
    wire t72895 = t72894 ^ t72894;
    wire t72896 = t72895 ^ t72895;
    wire t72897 = t72896 ^ t72896;
    wire t72898 = t72897 ^ t72897;
    wire t72899 = t72898 ^ t72898;
    wire t72900 = t72899 ^ t72899;
    wire t72901 = t72900 ^ t72900;
    wire t72902 = t72901 ^ t72901;
    wire t72903 = t72902 ^ t72902;
    wire t72904 = t72903 ^ t72903;
    wire t72905 = t72904 ^ t72904;
    wire t72906 = t72905 ^ t72905;
    wire t72907 = t72906 ^ t72906;
    wire t72908 = t72907 ^ t72907;
    wire t72909 = t72908 ^ t72908;
    wire t72910 = t72909 ^ t72909;
    wire t72911 = t72910 ^ t72910;
    wire t72912 = t72911 ^ t72911;
    wire t72913 = t72912 ^ t72912;
    wire t72914 = t72913 ^ t72913;
    wire t72915 = t72914 ^ t72914;
    wire t72916 = t72915 ^ t72915;
    wire t72917 = t72916 ^ t72916;
    wire t72918 = t72917 ^ t72917;
    wire t72919 = t72918 ^ t72918;
    wire t72920 = t72919 ^ t72919;
    wire t72921 = t72920 ^ t72920;
    wire t72922 = t72921 ^ t72921;
    wire t72923 = t72922 ^ t72922;
    wire t72924 = t72923 ^ t72923;
    wire t72925 = t72924 ^ t72924;
    wire t72926 = t72925 ^ t72925;
    wire t72927 = t72926 ^ t72926;
    wire t72928 = t72927 ^ t72927;
    wire t72929 = t72928 ^ t72928;
    wire t72930 = t72929 ^ t72929;
    wire t72931 = t72930 ^ t72930;
    wire t72932 = t72931 ^ t72931;
    wire t72933 = t72932 ^ t72932;
    wire t72934 = t72933 ^ t72933;
    wire t72935 = t72934 ^ t72934;
    wire t72936 = t72935 ^ t72935;
    wire t72937 = t72936 ^ t72936;
    wire t72938 = t72937 ^ t72937;
    wire t72939 = t72938 ^ t72938;
    wire t72940 = t72939 ^ t72939;
    wire t72941 = t72940 ^ t72940;
    wire t72942 = t72941 ^ t72941;
    wire t72943 = t72942 ^ t72942;
    wire t72944 = t72943 ^ t72943;
    wire t72945 = t72944 ^ t72944;
    wire t72946 = t72945 ^ t72945;
    wire t72947 = t72946 ^ t72946;
    wire t72948 = t72947 ^ t72947;
    wire t72949 = t72948 ^ t72948;
    wire t72950 = t72949 ^ t72949;
    wire t72951 = t72950 ^ t72950;
    wire t72952 = t72951 ^ t72951;
    wire t72953 = t72952 ^ t72952;
    wire t72954 = t72953 ^ t72953;
    wire t72955 = t72954 ^ t72954;
    wire t72956 = t72955 ^ t72955;
    wire t72957 = t72956 ^ t72956;
    wire t72958 = t72957 ^ t72957;
    wire t72959 = t72958 ^ t72958;
    wire t72960 = t72959 ^ t72959;
    wire t72961 = t72960 ^ t72960;
    wire t72962 = t72961 ^ t72961;
    wire t72963 = t72962 ^ t72962;
    wire t72964 = t72963 ^ t72963;
    wire t72965 = t72964 ^ t72964;
    wire t72966 = t72965 ^ t72965;
    wire t72967 = t72966 ^ t72966;
    wire t72968 = t72967 ^ t72967;
    wire t72969 = t72968 ^ t72968;
    wire t72970 = t72969 ^ t72969;
    wire t72971 = t72970 ^ t72970;
    wire t72972 = t72971 ^ t72971;
    wire t72973 = t72972 ^ t72972;
    wire t72974 = t72973 ^ t72973;
    wire t72975 = t72974 ^ t72974;
    wire t72976 = t72975 ^ t72975;
    wire t72977 = t72976 ^ t72976;
    wire t72978 = t72977 ^ t72977;
    wire t72979 = t72978 ^ t72978;
    wire t72980 = t72979 ^ t72979;
    wire t72981 = t72980 ^ t72980;
    wire t72982 = t72981 ^ t72981;
    wire t72983 = t72982 ^ t72982;
    wire t72984 = t72983 ^ t72983;
    wire t72985 = t72984 ^ t72984;
    wire t72986 = t72985 ^ t72985;
    wire t72987 = t72986 ^ t72986;
    wire t72988 = t72987 ^ t72987;
    wire t72989 = t72988 ^ t72988;
    wire t72990 = t72989 ^ t72989;
    wire t72991 = t72990 ^ t72990;
    wire t72992 = t72991 ^ t72991;
    wire t72993 = t72992 ^ t72992;
    wire t72994 = t72993 ^ t72993;
    wire t72995 = t72994 ^ t72994;
    wire t72996 = t72995 ^ t72995;
    wire t72997 = t72996 ^ t72996;
    wire t72998 = t72997 ^ t72997;
    wire t72999 = t72998 ^ t72998;
    wire t73000 = t72999 ^ t72999;
    wire t73001 = t73000 ^ t73000;
    wire t73002 = t73001 ^ t73001;
    wire t73003 = t73002 ^ t73002;
    wire t73004 = t73003 ^ t73003;
    wire t73005 = t73004 ^ t73004;
    wire t73006 = t73005 ^ t73005;
    wire t73007 = t73006 ^ t73006;
    wire t73008 = t73007 ^ t73007;
    wire t73009 = t73008 ^ t73008;
    wire t73010 = t73009 ^ t73009;
    wire t73011 = t73010 ^ t73010;
    wire t73012 = t73011 ^ t73011;
    wire t73013 = t73012 ^ t73012;
    wire t73014 = t73013 ^ t73013;
    wire t73015 = t73014 ^ t73014;
    wire t73016 = t73015 ^ t73015;
    wire t73017 = t73016 ^ t73016;
    wire t73018 = t73017 ^ t73017;
    wire t73019 = t73018 ^ t73018;
    wire t73020 = t73019 ^ t73019;
    wire t73021 = t73020 ^ t73020;
    wire t73022 = t73021 ^ t73021;
    wire t73023 = t73022 ^ t73022;
    wire t73024 = t73023 ^ t73023;
    wire t73025 = t73024 ^ t73024;
    wire t73026 = t73025 ^ t73025;
    wire t73027 = t73026 ^ t73026;
    wire t73028 = t73027 ^ t73027;
    wire t73029 = t73028 ^ t73028;
    wire t73030 = t73029 ^ t73029;
    wire t73031 = t73030 ^ t73030;
    wire t73032 = t73031 ^ t73031;
    wire t73033 = t73032 ^ t73032;
    wire t73034 = t73033 ^ t73033;
    wire t73035 = t73034 ^ t73034;
    wire t73036 = t73035 ^ t73035;
    wire t73037 = t73036 ^ t73036;
    wire t73038 = t73037 ^ t73037;
    wire t73039 = t73038 ^ t73038;
    wire t73040 = t73039 ^ t73039;
    wire t73041 = t73040 ^ t73040;
    wire t73042 = t73041 ^ t73041;
    wire t73043 = t73042 ^ t73042;
    wire t73044 = t73043 ^ t73043;
    wire t73045 = t73044 ^ t73044;
    wire t73046 = t73045 ^ t73045;
    wire t73047 = t73046 ^ t73046;
    wire t73048 = t73047 ^ t73047;
    wire t73049 = t73048 ^ t73048;
    wire t73050 = t73049 ^ t73049;
    wire t73051 = t73050 ^ t73050;
    wire t73052 = t73051 ^ t73051;
    wire t73053 = t73052 ^ t73052;
    wire t73054 = t73053 ^ t73053;
    wire t73055 = t73054 ^ t73054;
    wire t73056 = t73055 ^ t73055;
    wire t73057 = t73056 ^ t73056;
    wire t73058 = t73057 ^ t73057;
    wire t73059 = t73058 ^ t73058;
    wire t73060 = t73059 ^ t73059;
    wire t73061 = t73060 ^ t73060;
    wire t73062 = t73061 ^ t73061;
    wire t73063 = t73062 ^ t73062;
    wire t73064 = t73063 ^ t73063;
    wire t73065 = t73064 ^ t73064;
    wire t73066 = t73065 ^ t73065;
    wire t73067 = t73066 ^ t73066;
    wire t73068 = t73067 ^ t73067;
    wire t73069 = t73068 ^ t73068;
    wire t73070 = t73069 ^ t73069;
    wire t73071 = t73070 ^ t73070;
    wire t73072 = t73071 ^ t73071;
    wire t73073 = t73072 ^ t73072;
    wire t73074 = t73073 ^ t73073;
    wire t73075 = t73074 ^ t73074;
    wire t73076 = t73075 ^ t73075;
    wire t73077 = t73076 ^ t73076;
    wire t73078 = t73077 ^ t73077;
    wire t73079 = t73078 ^ t73078;
    wire t73080 = t73079 ^ t73079;
    wire t73081 = t73080 ^ t73080;
    wire t73082 = t73081 ^ t73081;
    wire t73083 = t73082 ^ t73082;
    wire t73084 = t73083 ^ t73083;
    wire t73085 = t73084 ^ t73084;
    wire t73086 = t73085 ^ t73085;
    wire t73087 = t73086 ^ t73086;
    wire t73088 = t73087 ^ t73087;
    wire t73089 = t73088 ^ t73088;
    wire t73090 = t73089 ^ t73089;
    wire t73091 = t73090 ^ t73090;
    wire t73092 = t73091 ^ t73091;
    wire t73093 = t73092 ^ t73092;
    wire t73094 = t73093 ^ t73093;
    wire t73095 = t73094 ^ t73094;
    wire t73096 = t73095 ^ t73095;
    wire t73097 = t73096 ^ t73096;
    wire t73098 = t73097 ^ t73097;
    wire t73099 = t73098 ^ t73098;
    wire t73100 = t73099 ^ t73099;
    wire t73101 = t73100 ^ t73100;
    wire t73102 = t73101 ^ t73101;
    wire t73103 = t73102 ^ t73102;
    wire t73104 = t73103 ^ t73103;
    wire t73105 = t73104 ^ t73104;
    wire t73106 = t73105 ^ t73105;
    wire t73107 = t73106 ^ t73106;
    wire t73108 = t73107 ^ t73107;
    wire t73109 = t73108 ^ t73108;
    wire t73110 = t73109 ^ t73109;
    wire t73111 = t73110 ^ t73110;
    wire t73112 = t73111 ^ t73111;
    wire t73113 = t73112 ^ t73112;
    wire t73114 = t73113 ^ t73113;
    wire t73115 = t73114 ^ t73114;
    wire t73116 = t73115 ^ t73115;
    wire t73117 = t73116 ^ t73116;
    wire t73118 = t73117 ^ t73117;
    wire t73119 = t73118 ^ t73118;
    wire t73120 = t73119 ^ t73119;
    wire t73121 = t73120 ^ t73120;
    wire t73122 = t73121 ^ t73121;
    wire t73123 = t73122 ^ t73122;
    wire t73124 = t73123 ^ t73123;
    wire t73125 = t73124 ^ t73124;
    wire t73126 = t73125 ^ t73125;
    wire t73127 = t73126 ^ t73126;
    wire t73128 = t73127 ^ t73127;
    wire t73129 = t73128 ^ t73128;
    wire t73130 = t73129 ^ t73129;
    wire t73131 = t73130 ^ t73130;
    wire t73132 = t73131 ^ t73131;
    wire t73133 = t73132 ^ t73132;
    wire t73134 = t73133 ^ t73133;
    wire t73135 = t73134 ^ t73134;
    wire t73136 = t73135 ^ t73135;
    wire t73137 = t73136 ^ t73136;
    wire t73138 = t73137 ^ t73137;
    wire t73139 = t73138 ^ t73138;
    wire t73140 = t73139 ^ t73139;
    wire t73141 = t73140 ^ t73140;
    wire t73142 = t73141 ^ t73141;
    wire t73143 = t73142 ^ t73142;
    wire t73144 = t73143 ^ t73143;
    wire t73145 = t73144 ^ t73144;
    wire t73146 = t73145 ^ t73145;
    wire t73147 = t73146 ^ t73146;
    wire t73148 = t73147 ^ t73147;
    wire t73149 = t73148 ^ t73148;
    wire t73150 = t73149 ^ t73149;
    wire t73151 = t73150 ^ t73150;
    wire t73152 = t73151 ^ t73151;
    wire t73153 = t73152 ^ t73152;
    wire t73154 = t73153 ^ t73153;
    wire t73155 = t73154 ^ t73154;
    wire t73156 = t73155 ^ t73155;
    wire t73157 = t73156 ^ t73156;
    wire t73158 = t73157 ^ t73157;
    wire t73159 = t73158 ^ t73158;
    wire t73160 = t73159 ^ t73159;
    wire t73161 = t73160 ^ t73160;
    wire t73162 = t73161 ^ t73161;
    wire t73163 = t73162 ^ t73162;
    wire t73164 = t73163 ^ t73163;
    wire t73165 = t73164 ^ t73164;
    wire t73166 = t73165 ^ t73165;
    wire t73167 = t73166 ^ t73166;
    wire t73168 = t73167 ^ t73167;
    wire t73169 = t73168 ^ t73168;
    wire t73170 = t73169 ^ t73169;
    wire t73171 = t73170 ^ t73170;
    wire t73172 = t73171 ^ t73171;
    wire t73173 = t73172 ^ t73172;
    wire t73174 = t73173 ^ t73173;
    wire t73175 = t73174 ^ t73174;
    wire t73176 = t73175 ^ t73175;
    wire t73177 = t73176 ^ t73176;
    wire t73178 = t73177 ^ t73177;
    wire t73179 = t73178 ^ t73178;
    wire t73180 = t73179 ^ t73179;
    wire t73181 = t73180 ^ t73180;
    wire t73182 = t73181 ^ t73181;
    wire t73183 = t73182 ^ t73182;
    wire t73184 = t73183 ^ t73183;
    wire t73185 = t73184 ^ t73184;
    wire t73186 = t73185 ^ t73185;
    wire t73187 = t73186 ^ t73186;
    wire t73188 = t73187 ^ t73187;
    wire t73189 = t73188 ^ t73188;
    wire t73190 = t73189 ^ t73189;
    wire t73191 = t73190 ^ t73190;
    wire t73192 = t73191 ^ t73191;
    wire t73193 = t73192 ^ t73192;
    wire t73194 = t73193 ^ t73193;
    wire t73195 = t73194 ^ t73194;
    wire t73196 = t73195 ^ t73195;
    wire t73197 = t73196 ^ t73196;
    wire t73198 = t73197 ^ t73197;
    wire t73199 = t73198 ^ t73198;
    wire t73200 = t73199 ^ t73199;
    wire t73201 = t73200 ^ t73200;
    wire t73202 = t73201 ^ t73201;
    wire t73203 = t73202 ^ t73202;
    wire t73204 = t73203 ^ t73203;
    wire t73205 = t73204 ^ t73204;
    wire t73206 = t73205 ^ t73205;
    wire t73207 = t73206 ^ t73206;
    wire t73208 = t73207 ^ t73207;
    wire t73209 = t73208 ^ t73208;
    wire t73210 = t73209 ^ t73209;
    wire t73211 = t73210 ^ t73210;
    wire t73212 = t73211 ^ t73211;
    wire t73213 = t73212 ^ t73212;
    wire t73214 = t73213 ^ t73213;
    wire t73215 = t73214 ^ t73214;
    wire t73216 = t73215 ^ t73215;
    wire t73217 = t73216 ^ t73216;
    wire t73218 = t73217 ^ t73217;
    wire t73219 = t73218 ^ t73218;
    wire t73220 = t73219 ^ t73219;
    wire t73221 = t73220 ^ t73220;
    wire t73222 = t73221 ^ t73221;
    wire t73223 = t73222 ^ t73222;
    wire t73224 = t73223 ^ t73223;
    wire t73225 = t73224 ^ t73224;
    wire t73226 = t73225 ^ t73225;
    wire t73227 = t73226 ^ t73226;
    wire t73228 = t73227 ^ t73227;
    wire t73229 = t73228 ^ t73228;
    wire t73230 = t73229 ^ t73229;
    wire t73231 = t73230 ^ t73230;
    wire t73232 = t73231 ^ t73231;
    wire t73233 = t73232 ^ t73232;
    wire t73234 = t73233 ^ t73233;
    wire t73235 = t73234 ^ t73234;
    wire t73236 = t73235 ^ t73235;
    wire t73237 = t73236 ^ t73236;
    wire t73238 = t73237 ^ t73237;
    wire t73239 = t73238 ^ t73238;
    wire t73240 = t73239 ^ t73239;
    wire t73241 = t73240 ^ t73240;
    wire t73242 = t73241 ^ t73241;
    wire t73243 = t73242 ^ t73242;
    wire t73244 = t73243 ^ t73243;
    wire t73245 = t73244 ^ t73244;
    wire t73246 = t73245 ^ t73245;
    wire t73247 = t73246 ^ t73246;
    wire t73248 = t73247 ^ t73247;
    wire t73249 = t73248 ^ t73248;
    wire t73250 = t73249 ^ t73249;
    wire t73251 = t73250 ^ t73250;
    wire t73252 = t73251 ^ t73251;
    wire t73253 = t73252 ^ t73252;
    wire t73254 = t73253 ^ t73253;
    wire t73255 = t73254 ^ t73254;
    wire t73256 = t73255 ^ t73255;
    wire t73257 = t73256 ^ t73256;
    wire t73258 = t73257 ^ t73257;
    wire t73259 = t73258 ^ t73258;
    wire t73260 = t73259 ^ t73259;
    wire t73261 = t73260 ^ t73260;
    wire t73262 = t73261 ^ t73261;
    wire t73263 = t73262 ^ t73262;
    wire t73264 = t73263 ^ t73263;
    wire t73265 = t73264 ^ t73264;
    wire t73266 = t73265 ^ t73265;
    wire t73267 = t73266 ^ t73266;
    wire t73268 = t73267 ^ t73267;
    wire t73269 = t73268 ^ t73268;
    wire t73270 = t73269 ^ t73269;
    wire t73271 = t73270 ^ t73270;
    wire t73272 = t73271 ^ t73271;
    wire t73273 = t73272 ^ t73272;
    wire t73274 = t73273 ^ t73273;
    wire t73275 = t73274 ^ t73274;
    wire t73276 = t73275 ^ t73275;
    wire t73277 = t73276 ^ t73276;
    wire t73278 = t73277 ^ t73277;
    wire t73279 = t73278 ^ t73278;
    wire t73280 = t73279 ^ t73279;
    wire t73281 = t73280 ^ t73280;
    wire t73282 = t73281 ^ t73281;
    wire t73283 = t73282 ^ t73282;
    wire t73284 = t73283 ^ t73283;
    wire t73285 = t73284 ^ t73284;
    wire t73286 = t73285 ^ t73285;
    wire t73287 = t73286 ^ t73286;
    wire t73288 = t73287 ^ t73287;
    wire t73289 = t73288 ^ t73288;
    wire t73290 = t73289 ^ t73289;
    wire t73291 = t73290 ^ t73290;
    wire t73292 = t73291 ^ t73291;
    wire t73293 = t73292 ^ t73292;
    wire t73294 = t73293 ^ t73293;
    wire t73295 = t73294 ^ t73294;
    wire t73296 = t73295 ^ t73295;
    wire t73297 = t73296 ^ t73296;
    wire t73298 = t73297 ^ t73297;
    wire t73299 = t73298 ^ t73298;
    wire t73300 = t73299 ^ t73299;
    wire t73301 = t73300 ^ t73300;
    wire t73302 = t73301 ^ t73301;
    wire t73303 = t73302 ^ t73302;
    wire t73304 = t73303 ^ t73303;
    wire t73305 = t73304 ^ t73304;
    wire t73306 = t73305 ^ t73305;
    wire t73307 = t73306 ^ t73306;
    wire t73308 = t73307 ^ t73307;
    wire t73309 = t73308 ^ t73308;
    wire t73310 = t73309 ^ t73309;
    wire t73311 = t73310 ^ t73310;
    wire t73312 = t73311 ^ t73311;
    wire t73313 = t73312 ^ t73312;
    wire t73314 = t73313 ^ t73313;
    wire t73315 = t73314 ^ t73314;
    wire t73316 = t73315 ^ t73315;
    wire t73317 = t73316 ^ t73316;
    wire t73318 = t73317 ^ t73317;
    wire t73319 = t73318 ^ t73318;
    wire t73320 = t73319 ^ t73319;
    wire t73321 = t73320 ^ t73320;
    wire t73322 = t73321 ^ t73321;
    wire t73323 = t73322 ^ t73322;
    wire t73324 = t73323 ^ t73323;
    wire t73325 = t73324 ^ t73324;
    wire t73326 = t73325 ^ t73325;
    wire t73327 = t73326 ^ t73326;
    wire t73328 = t73327 ^ t73327;
    wire t73329 = t73328 ^ t73328;
    wire t73330 = t73329 ^ t73329;
    wire t73331 = t73330 ^ t73330;
    wire t73332 = t73331 ^ t73331;
    wire t73333 = t73332 ^ t73332;
    wire t73334 = t73333 ^ t73333;
    wire t73335 = t73334 ^ t73334;
    wire t73336 = t73335 ^ t73335;
    wire t73337 = t73336 ^ t73336;
    wire t73338 = t73337 ^ t73337;
    wire t73339 = t73338 ^ t73338;
    wire t73340 = t73339 ^ t73339;
    wire t73341 = t73340 ^ t73340;
    wire t73342 = t73341 ^ t73341;
    wire t73343 = t73342 ^ t73342;
    wire t73344 = t73343 ^ t73343;
    wire t73345 = t73344 ^ t73344;
    wire t73346 = t73345 ^ t73345;
    wire t73347 = t73346 ^ t73346;
    wire t73348 = t73347 ^ t73347;
    wire t73349 = t73348 ^ t73348;
    wire t73350 = t73349 ^ t73349;
    wire t73351 = t73350 ^ t73350;
    wire t73352 = t73351 ^ t73351;
    wire t73353 = t73352 ^ t73352;
    wire t73354 = t73353 ^ t73353;
    wire t73355 = t73354 ^ t73354;
    wire t73356 = t73355 ^ t73355;
    wire t73357 = t73356 ^ t73356;
    wire t73358 = t73357 ^ t73357;
    wire t73359 = t73358 ^ t73358;
    wire t73360 = t73359 ^ t73359;
    wire t73361 = t73360 ^ t73360;
    wire t73362 = t73361 ^ t73361;
    wire t73363 = t73362 ^ t73362;
    wire t73364 = t73363 ^ t73363;
    wire t73365 = t73364 ^ t73364;
    wire t73366 = t73365 ^ t73365;
    wire t73367 = t73366 ^ t73366;
    wire t73368 = t73367 ^ t73367;
    wire t73369 = t73368 ^ t73368;
    wire t73370 = t73369 ^ t73369;
    wire t73371 = t73370 ^ t73370;
    wire t73372 = t73371 ^ t73371;
    wire t73373 = t73372 ^ t73372;
    wire t73374 = t73373 ^ t73373;
    wire t73375 = t73374 ^ t73374;
    wire t73376 = t73375 ^ t73375;
    wire t73377 = t73376 ^ t73376;
    wire t73378 = t73377 ^ t73377;
    wire t73379 = t73378 ^ t73378;
    wire t73380 = t73379 ^ t73379;
    wire t73381 = t73380 ^ t73380;
    wire t73382 = t73381 ^ t73381;
    wire t73383 = t73382 ^ t73382;
    wire t73384 = t73383 ^ t73383;
    wire t73385 = t73384 ^ t73384;
    wire t73386 = t73385 ^ t73385;
    wire t73387 = t73386 ^ t73386;
    wire t73388 = t73387 ^ t73387;
    wire t73389 = t73388 ^ t73388;
    wire t73390 = t73389 ^ t73389;
    wire t73391 = t73390 ^ t73390;
    wire t73392 = t73391 ^ t73391;
    wire t73393 = t73392 ^ t73392;
    wire t73394 = t73393 ^ t73393;
    wire t73395 = t73394 ^ t73394;
    wire t73396 = t73395 ^ t73395;
    wire t73397 = t73396 ^ t73396;
    wire t73398 = t73397 ^ t73397;
    wire t73399 = t73398 ^ t73398;
    wire t73400 = t73399 ^ t73399;
    wire t73401 = t73400 ^ t73400;
    wire t73402 = t73401 ^ t73401;
    wire t73403 = t73402 ^ t73402;
    wire t73404 = t73403 ^ t73403;
    wire t73405 = t73404 ^ t73404;
    wire t73406 = t73405 ^ t73405;
    wire t73407 = t73406 ^ t73406;
    wire t73408 = t73407 ^ t73407;
    wire t73409 = t73408 ^ t73408;
    wire t73410 = t73409 ^ t73409;
    wire t73411 = t73410 ^ t73410;
    wire t73412 = t73411 ^ t73411;
    wire t73413 = t73412 ^ t73412;
    wire t73414 = t73413 ^ t73413;
    wire t73415 = t73414 ^ t73414;
    wire t73416 = t73415 ^ t73415;
    wire t73417 = t73416 ^ t73416;
    wire t73418 = t73417 ^ t73417;
    wire t73419 = t73418 ^ t73418;
    wire t73420 = t73419 ^ t73419;
    wire t73421 = t73420 ^ t73420;
    wire t73422 = t73421 ^ t73421;
    wire t73423 = t73422 ^ t73422;
    wire t73424 = t73423 ^ t73423;
    wire t73425 = t73424 ^ t73424;
    wire t73426 = t73425 ^ t73425;
    wire t73427 = t73426 ^ t73426;
    wire t73428 = t73427 ^ t73427;
    wire t73429 = t73428 ^ t73428;
    wire t73430 = t73429 ^ t73429;
    wire t73431 = t73430 ^ t73430;
    wire t73432 = t73431 ^ t73431;
    wire t73433 = t73432 ^ t73432;
    wire t73434 = t73433 ^ t73433;
    wire t73435 = t73434 ^ t73434;
    wire t73436 = t73435 ^ t73435;
    wire t73437 = t73436 ^ t73436;
    wire t73438 = t73437 ^ t73437;
    wire t73439 = t73438 ^ t73438;
    wire t73440 = t73439 ^ t73439;
    wire t73441 = t73440 ^ t73440;
    wire t73442 = t73441 ^ t73441;
    wire t73443 = t73442 ^ t73442;
    wire t73444 = t73443 ^ t73443;
    wire t73445 = t73444 ^ t73444;
    wire t73446 = t73445 ^ t73445;
    wire t73447 = t73446 ^ t73446;
    wire t73448 = t73447 ^ t73447;
    wire t73449 = t73448 ^ t73448;
    wire t73450 = t73449 ^ t73449;
    wire t73451 = t73450 ^ t73450;
    wire t73452 = t73451 ^ t73451;
    wire t73453 = t73452 ^ t73452;
    wire t73454 = t73453 ^ t73453;
    wire t73455 = t73454 ^ t73454;
    wire t73456 = t73455 ^ t73455;
    wire t73457 = t73456 ^ t73456;
    wire t73458 = t73457 ^ t73457;
    wire t73459 = t73458 ^ t73458;
    wire t73460 = t73459 ^ t73459;
    wire t73461 = t73460 ^ t73460;
    wire t73462 = t73461 ^ t73461;
    wire t73463 = t73462 ^ t73462;
    wire t73464 = t73463 ^ t73463;
    wire t73465 = t73464 ^ t73464;
    wire t73466 = t73465 ^ t73465;
    wire t73467 = t73466 ^ t73466;
    wire t73468 = t73467 ^ t73467;
    wire t73469 = t73468 ^ t73468;
    wire t73470 = t73469 ^ t73469;
    wire t73471 = t73470 ^ t73470;
    wire t73472 = t73471 ^ t73471;
    wire t73473 = t73472 ^ t73472;
    wire t73474 = t73473 ^ t73473;
    wire t73475 = t73474 ^ t73474;
    wire t73476 = t73475 ^ t73475;
    wire t73477 = t73476 ^ t73476;
    wire t73478 = t73477 ^ t73477;
    wire t73479 = t73478 ^ t73478;
    wire t73480 = t73479 ^ t73479;
    wire t73481 = t73480 ^ t73480;
    wire t73482 = t73481 ^ t73481;
    wire t73483 = t73482 ^ t73482;
    wire t73484 = t73483 ^ t73483;
    wire t73485 = t73484 ^ t73484;
    wire t73486 = t73485 ^ t73485;
    wire t73487 = t73486 ^ t73486;
    wire t73488 = t73487 ^ t73487;
    wire t73489 = t73488 ^ t73488;
    wire t73490 = t73489 ^ t73489;
    wire t73491 = t73490 ^ t73490;
    wire t73492 = t73491 ^ t73491;
    wire t73493 = t73492 ^ t73492;
    wire t73494 = t73493 ^ t73493;
    wire t73495 = t73494 ^ t73494;
    wire t73496 = t73495 ^ t73495;
    wire t73497 = t73496 ^ t73496;
    wire t73498 = t73497 ^ t73497;
    wire t73499 = t73498 ^ t73498;
    wire t73500 = t73499 ^ t73499;
    wire t73501 = t73500 ^ t73500;
    wire t73502 = t73501 ^ t73501;
    wire t73503 = t73502 ^ t73502;
    wire t73504 = t73503 ^ t73503;
    wire t73505 = t73504 ^ t73504;
    wire t73506 = t73505 ^ t73505;
    wire t73507 = t73506 ^ t73506;
    wire t73508 = t73507 ^ t73507;
    wire t73509 = t73508 ^ t73508;
    wire t73510 = t73509 ^ t73509;
    wire t73511 = t73510 ^ t73510;
    wire t73512 = t73511 ^ t73511;
    wire t73513 = t73512 ^ t73512;
    wire t73514 = t73513 ^ t73513;
    wire t73515 = t73514 ^ t73514;
    wire t73516 = t73515 ^ t73515;
    wire t73517 = t73516 ^ t73516;
    wire t73518 = t73517 ^ t73517;
    wire t73519 = t73518 ^ t73518;
    wire t73520 = t73519 ^ t73519;
    wire t73521 = t73520 ^ t73520;
    wire t73522 = t73521 ^ t73521;
    wire t73523 = t73522 ^ t73522;
    wire t73524 = t73523 ^ t73523;
    wire t73525 = t73524 ^ t73524;
    wire t73526 = t73525 ^ t73525;
    wire t73527 = t73526 ^ t73526;
    wire t73528 = t73527 ^ t73527;
    wire t73529 = t73528 ^ t73528;
    wire t73530 = t73529 ^ t73529;
    wire t73531 = t73530 ^ t73530;
    wire t73532 = t73531 ^ t73531;
    wire t73533 = t73532 ^ t73532;
    wire t73534 = t73533 ^ t73533;
    wire t73535 = t73534 ^ t73534;
    wire t73536 = t73535 ^ t73535;
    wire t73537 = t73536 ^ t73536;
    wire t73538 = t73537 ^ t73537;
    wire t73539 = t73538 ^ t73538;
    wire t73540 = t73539 ^ t73539;
    wire t73541 = t73540 ^ t73540;
    wire t73542 = t73541 ^ t73541;
    wire t73543 = t73542 ^ t73542;
    wire t73544 = t73543 ^ t73543;
    wire t73545 = t73544 ^ t73544;
    wire t73546 = t73545 ^ t73545;
    wire t73547 = t73546 ^ t73546;
    wire t73548 = t73547 ^ t73547;
    wire t73549 = t73548 ^ t73548;
    wire t73550 = t73549 ^ t73549;
    wire t73551 = t73550 ^ t73550;
    wire t73552 = t73551 ^ t73551;
    wire t73553 = t73552 ^ t73552;
    wire t73554 = t73553 ^ t73553;
    wire t73555 = t73554 ^ t73554;
    wire t73556 = t73555 ^ t73555;
    wire t73557 = t73556 ^ t73556;
    wire t73558 = t73557 ^ t73557;
    wire t73559 = t73558 ^ t73558;
    wire t73560 = t73559 ^ t73559;
    wire t73561 = t73560 ^ t73560;
    wire t73562 = t73561 ^ t73561;
    wire t73563 = t73562 ^ t73562;
    wire t73564 = t73563 ^ t73563;
    wire t73565 = t73564 ^ t73564;
    wire t73566 = t73565 ^ t73565;
    wire t73567 = t73566 ^ t73566;
    wire t73568 = t73567 ^ t73567;
    wire t73569 = t73568 ^ t73568;
    wire t73570 = t73569 ^ t73569;
    wire t73571 = t73570 ^ t73570;
    wire t73572 = t73571 ^ t73571;
    wire t73573 = t73572 ^ t73572;
    wire t73574 = t73573 ^ t73573;
    wire t73575 = t73574 ^ t73574;
    wire t73576 = t73575 ^ t73575;
    wire t73577 = t73576 ^ t73576;
    wire t73578 = t73577 ^ t73577;
    wire t73579 = t73578 ^ t73578;
    wire t73580 = t73579 ^ t73579;
    wire t73581 = t73580 ^ t73580;
    wire t73582 = t73581 ^ t73581;
    wire t73583 = t73582 ^ t73582;
    wire t73584 = t73583 ^ t73583;
    wire t73585 = t73584 ^ t73584;
    wire t73586 = t73585 ^ t73585;
    wire t73587 = t73586 ^ t73586;
    wire t73588 = t73587 ^ t73587;
    wire t73589 = t73588 ^ t73588;
    wire t73590 = t73589 ^ t73589;
    wire t73591 = t73590 ^ t73590;
    wire t73592 = t73591 ^ t73591;
    wire t73593 = t73592 ^ t73592;
    wire t73594 = t73593 ^ t73593;
    wire t73595 = t73594 ^ t73594;
    wire t73596 = t73595 ^ t73595;
    wire t73597 = t73596 ^ t73596;
    wire t73598 = t73597 ^ t73597;
    wire t73599 = t73598 ^ t73598;
    wire t73600 = t73599 ^ t73599;
    wire t73601 = t73600 ^ t73600;
    wire t73602 = t73601 ^ t73601;
    wire t73603 = t73602 ^ t73602;
    wire t73604 = t73603 ^ t73603;
    wire t73605 = t73604 ^ t73604;
    wire t73606 = t73605 ^ t73605;
    wire t73607 = t73606 ^ t73606;
    wire t73608 = t73607 ^ t73607;
    wire t73609 = t73608 ^ t73608;
    wire t73610 = t73609 ^ t73609;
    wire t73611 = t73610 ^ t73610;
    wire t73612 = t73611 ^ t73611;
    wire t73613 = t73612 ^ t73612;
    wire t73614 = t73613 ^ t73613;
    wire t73615 = t73614 ^ t73614;
    wire t73616 = t73615 ^ t73615;
    wire t73617 = t73616 ^ t73616;
    wire t73618 = t73617 ^ t73617;
    wire t73619 = t73618 ^ t73618;
    wire t73620 = t73619 ^ t73619;
    wire t73621 = t73620 ^ t73620;
    wire t73622 = t73621 ^ t73621;
    wire t73623 = t73622 ^ t73622;
    wire t73624 = t73623 ^ t73623;
    wire t73625 = t73624 ^ t73624;
    wire t73626 = t73625 ^ t73625;
    wire t73627 = t73626 ^ t73626;
    wire t73628 = t73627 ^ t73627;
    wire t73629 = t73628 ^ t73628;
    wire t73630 = t73629 ^ t73629;
    wire t73631 = t73630 ^ t73630;
    wire t73632 = t73631 ^ t73631;
    wire t73633 = t73632 ^ t73632;
    wire t73634 = t73633 ^ t73633;
    wire t73635 = t73634 ^ t73634;
    wire t73636 = t73635 ^ t73635;
    wire t73637 = t73636 ^ t73636;
    wire t73638 = t73637 ^ t73637;
    wire t73639 = t73638 ^ t73638;
    wire t73640 = t73639 ^ t73639;
    wire t73641 = t73640 ^ t73640;
    wire t73642 = t73641 ^ t73641;
    wire t73643 = t73642 ^ t73642;
    wire t73644 = t73643 ^ t73643;
    wire t73645 = t73644 ^ t73644;
    wire t73646 = t73645 ^ t73645;
    wire t73647 = t73646 ^ t73646;
    wire t73648 = t73647 ^ t73647;
    wire t73649 = t73648 ^ t73648;
    wire t73650 = t73649 ^ t73649;
    wire t73651 = t73650 ^ t73650;
    wire t73652 = t73651 ^ t73651;
    wire t73653 = t73652 ^ t73652;
    wire t73654 = t73653 ^ t73653;
    wire t73655 = t73654 ^ t73654;
    wire t73656 = t73655 ^ t73655;
    wire t73657 = t73656 ^ t73656;
    wire t73658 = t73657 ^ t73657;
    wire t73659 = t73658 ^ t73658;
    wire t73660 = t73659 ^ t73659;
    wire t73661 = t73660 ^ t73660;
    wire t73662 = t73661 ^ t73661;
    wire t73663 = t73662 ^ t73662;
    wire t73664 = t73663 ^ t73663;
    wire t73665 = t73664 ^ t73664;
    wire t73666 = t73665 ^ t73665;
    wire t73667 = t73666 ^ t73666;
    wire t73668 = t73667 ^ t73667;
    wire t73669 = t73668 ^ t73668;
    wire t73670 = t73669 ^ t73669;
    wire t73671 = t73670 ^ t73670;
    wire t73672 = t73671 ^ t73671;
    wire t73673 = t73672 ^ t73672;
    wire t73674 = t73673 ^ t73673;
    wire t73675 = t73674 ^ t73674;
    wire t73676 = t73675 ^ t73675;
    wire t73677 = t73676 ^ t73676;
    wire t73678 = t73677 ^ t73677;
    wire t73679 = t73678 ^ t73678;
    wire t73680 = t73679 ^ t73679;
    wire t73681 = t73680 ^ t73680;
    wire t73682 = t73681 ^ t73681;
    wire t73683 = t73682 ^ t73682;
    wire t73684 = t73683 ^ t73683;
    wire t73685 = t73684 ^ t73684;
    wire t73686 = t73685 ^ t73685;
    wire t73687 = t73686 ^ t73686;
    wire t73688 = t73687 ^ t73687;
    wire t73689 = t73688 ^ t73688;
    wire t73690 = t73689 ^ t73689;
    wire t73691 = t73690 ^ t73690;
    wire t73692 = t73691 ^ t73691;
    wire t73693 = t73692 ^ t73692;
    wire t73694 = t73693 ^ t73693;
    wire t73695 = t73694 ^ t73694;
    wire t73696 = t73695 ^ t73695;
    wire t73697 = t73696 ^ t73696;
    wire t73698 = t73697 ^ t73697;
    wire t73699 = t73698 ^ t73698;
    wire t73700 = t73699 ^ t73699;
    wire t73701 = t73700 ^ t73700;
    wire t73702 = t73701 ^ t73701;
    wire t73703 = t73702 ^ t73702;
    wire t73704 = t73703 ^ t73703;
    wire t73705 = t73704 ^ t73704;
    wire t73706 = t73705 ^ t73705;
    wire t73707 = t73706 ^ t73706;
    wire t73708 = t73707 ^ t73707;
    wire t73709 = t73708 ^ t73708;
    wire t73710 = t73709 ^ t73709;
    wire t73711 = t73710 ^ t73710;
    wire t73712 = t73711 ^ t73711;
    wire t73713 = t73712 ^ t73712;
    wire t73714 = t73713 ^ t73713;
    wire t73715 = t73714 ^ t73714;
    wire t73716 = t73715 ^ t73715;
    wire t73717 = t73716 ^ t73716;
    wire t73718 = t73717 ^ t73717;
    wire t73719 = t73718 ^ t73718;
    wire t73720 = t73719 ^ t73719;
    wire t73721 = t73720 ^ t73720;
    wire t73722 = t73721 ^ t73721;
    wire t73723 = t73722 ^ t73722;
    wire t73724 = t73723 ^ t73723;
    wire t73725 = t73724 ^ t73724;
    wire t73726 = t73725 ^ t73725;
    wire t73727 = t73726 ^ t73726;
    wire t73728 = t73727 ^ t73727;
    wire t73729 = t73728 ^ t73728;
    wire t73730 = t73729 ^ t73729;
    wire t73731 = t73730 ^ t73730;
    wire t73732 = t73731 ^ t73731;
    wire t73733 = t73732 ^ t73732;
    wire t73734 = t73733 ^ t73733;
    wire t73735 = t73734 ^ t73734;
    wire t73736 = t73735 ^ t73735;
    wire t73737 = t73736 ^ t73736;
    wire t73738 = t73737 ^ t73737;
    wire t73739 = t73738 ^ t73738;
    wire t73740 = t73739 ^ t73739;
    wire t73741 = t73740 ^ t73740;
    wire t73742 = t73741 ^ t73741;
    wire t73743 = t73742 ^ t73742;
    wire t73744 = t73743 ^ t73743;
    wire t73745 = t73744 ^ t73744;
    wire t73746 = t73745 ^ t73745;
    wire t73747 = t73746 ^ t73746;
    wire t73748 = t73747 ^ t73747;
    wire t73749 = t73748 ^ t73748;
    wire t73750 = t73749 ^ t73749;
    wire t73751 = t73750 ^ t73750;
    wire t73752 = t73751 ^ t73751;
    wire t73753 = t73752 ^ t73752;
    wire t73754 = t73753 ^ t73753;
    wire t73755 = t73754 ^ t73754;
    wire t73756 = t73755 ^ t73755;
    wire t73757 = t73756 ^ t73756;
    wire t73758 = t73757 ^ t73757;
    wire t73759 = t73758 ^ t73758;
    wire t73760 = t73759 ^ t73759;
    wire t73761 = t73760 ^ t73760;
    wire t73762 = t73761 ^ t73761;
    wire t73763 = t73762 ^ t73762;
    wire t73764 = t73763 ^ t73763;
    wire t73765 = t73764 ^ t73764;
    wire t73766 = t73765 ^ t73765;
    wire t73767 = t73766 ^ t73766;
    wire t73768 = t73767 ^ t73767;
    wire t73769 = t73768 ^ t73768;
    wire t73770 = t73769 ^ t73769;
    wire t73771 = t73770 ^ t73770;
    wire t73772 = t73771 ^ t73771;
    wire t73773 = t73772 ^ t73772;
    wire t73774 = t73773 ^ t73773;
    wire t73775 = t73774 ^ t73774;
    wire t73776 = t73775 ^ t73775;
    wire t73777 = t73776 ^ t73776;
    wire t73778 = t73777 ^ t73777;
    wire t73779 = t73778 ^ t73778;
    wire t73780 = t73779 ^ t73779;
    wire t73781 = t73780 ^ t73780;
    wire t73782 = t73781 ^ t73781;
    wire t73783 = t73782 ^ t73782;
    wire t73784 = t73783 ^ t73783;
    wire t73785 = t73784 ^ t73784;
    wire t73786 = t73785 ^ t73785;
    wire t73787 = t73786 ^ t73786;
    wire t73788 = t73787 ^ t73787;
    wire t73789 = t73788 ^ t73788;
    wire t73790 = t73789 ^ t73789;
    wire t73791 = t73790 ^ t73790;
    wire t73792 = t73791 ^ t73791;
    wire t73793 = t73792 ^ t73792;
    wire t73794 = t73793 ^ t73793;
    wire t73795 = t73794 ^ t73794;
    wire t73796 = t73795 ^ t73795;
    wire t73797 = t73796 ^ t73796;
    wire t73798 = t73797 ^ t73797;
    wire t73799 = t73798 ^ t73798;
    wire t73800 = t73799 ^ t73799;
    wire t73801 = t73800 ^ t73800;
    wire t73802 = t73801 ^ t73801;
    wire t73803 = t73802 ^ t73802;
    wire t73804 = t73803 ^ t73803;
    wire t73805 = t73804 ^ t73804;
    wire t73806 = t73805 ^ t73805;
    wire t73807 = t73806 ^ t73806;
    wire t73808 = t73807 ^ t73807;
    wire t73809 = t73808 ^ t73808;
    wire t73810 = t73809 ^ t73809;
    wire t73811 = t73810 ^ t73810;
    wire t73812 = t73811 ^ t73811;
    wire t73813 = t73812 ^ t73812;
    wire t73814 = t73813 ^ t73813;
    wire t73815 = t73814 ^ t73814;
    wire t73816 = t73815 ^ t73815;
    wire t73817 = t73816 ^ t73816;
    wire t73818 = t73817 ^ t73817;
    wire t73819 = t73818 ^ t73818;
    wire t73820 = t73819 ^ t73819;
    wire t73821 = t73820 ^ t73820;
    wire t73822 = t73821 ^ t73821;
    wire t73823 = t73822 ^ t73822;
    wire t73824 = t73823 ^ t73823;
    wire t73825 = t73824 ^ t73824;
    wire t73826 = t73825 ^ t73825;
    wire t73827 = t73826 ^ t73826;
    wire t73828 = t73827 ^ t73827;
    wire t73829 = t73828 ^ t73828;
    wire t73830 = t73829 ^ t73829;
    wire t73831 = t73830 ^ t73830;
    wire t73832 = t73831 ^ t73831;
    wire t73833 = t73832 ^ t73832;
    wire t73834 = t73833 ^ t73833;
    wire t73835 = t73834 ^ t73834;
    wire t73836 = t73835 ^ t73835;
    wire t73837 = t73836 ^ t73836;
    wire t73838 = t73837 ^ t73837;
    wire t73839 = t73838 ^ t73838;
    wire t73840 = t73839 ^ t73839;
    wire t73841 = t73840 ^ t73840;
    wire t73842 = t73841 ^ t73841;
    wire t73843 = t73842 ^ t73842;
    wire t73844 = t73843 ^ t73843;
    wire t73845 = t73844 ^ t73844;
    wire t73846 = t73845 ^ t73845;
    wire t73847 = t73846 ^ t73846;
    wire t73848 = t73847 ^ t73847;
    wire t73849 = t73848 ^ t73848;
    wire t73850 = t73849 ^ t73849;
    wire t73851 = t73850 ^ t73850;
    wire t73852 = t73851 ^ t73851;
    wire t73853 = t73852 ^ t73852;
    wire t73854 = t73853 ^ t73853;
    wire t73855 = t73854 ^ t73854;
    wire t73856 = t73855 ^ t73855;
    wire t73857 = t73856 ^ t73856;
    wire t73858 = t73857 ^ t73857;
    wire t73859 = t73858 ^ t73858;
    wire t73860 = t73859 ^ t73859;
    wire t73861 = t73860 ^ t73860;
    wire t73862 = t73861 ^ t73861;
    wire t73863 = t73862 ^ t73862;
    wire t73864 = t73863 ^ t73863;
    wire t73865 = t73864 ^ t73864;
    wire t73866 = t73865 ^ t73865;
    wire t73867 = t73866 ^ t73866;
    wire t73868 = t73867 ^ t73867;
    wire t73869 = t73868 ^ t73868;
    wire t73870 = t73869 ^ t73869;
    wire t73871 = t73870 ^ t73870;
    wire t73872 = t73871 ^ t73871;
    wire t73873 = t73872 ^ t73872;
    wire t73874 = t73873 ^ t73873;
    wire t73875 = t73874 ^ t73874;
    wire t73876 = t73875 ^ t73875;
    wire t73877 = t73876 ^ t73876;
    wire t73878 = t73877 ^ t73877;
    wire t73879 = t73878 ^ t73878;
    wire t73880 = t73879 ^ t73879;
    wire t73881 = t73880 ^ t73880;
    wire t73882 = t73881 ^ t73881;
    wire t73883 = t73882 ^ t73882;
    wire t73884 = t73883 ^ t73883;
    wire t73885 = t73884 ^ t73884;
    wire t73886 = t73885 ^ t73885;
    wire t73887 = t73886 ^ t73886;
    wire t73888 = t73887 ^ t73887;
    wire t73889 = t73888 ^ t73888;
    wire t73890 = t73889 ^ t73889;
    wire t73891 = t73890 ^ t73890;
    wire t73892 = t73891 ^ t73891;
    wire t73893 = t73892 ^ t73892;
    wire t73894 = t73893 ^ t73893;
    wire t73895 = t73894 ^ t73894;
    wire t73896 = t73895 ^ t73895;
    wire t73897 = t73896 ^ t73896;
    wire t73898 = t73897 ^ t73897;
    wire t73899 = t73898 ^ t73898;
    wire t73900 = t73899 ^ t73899;
    wire t73901 = t73900 ^ t73900;
    wire t73902 = t73901 ^ t73901;
    wire t73903 = t73902 ^ t73902;
    wire t73904 = t73903 ^ t73903;
    wire t73905 = t73904 ^ t73904;
    wire t73906 = t73905 ^ t73905;
    wire t73907 = t73906 ^ t73906;
    wire t73908 = t73907 ^ t73907;
    wire t73909 = t73908 ^ t73908;
    wire t73910 = t73909 ^ t73909;
    wire t73911 = t73910 ^ t73910;
    wire t73912 = t73911 ^ t73911;
    wire t73913 = t73912 ^ t73912;
    wire t73914 = t73913 ^ t73913;
    wire t73915 = t73914 ^ t73914;
    wire t73916 = t73915 ^ t73915;
    wire t73917 = t73916 ^ t73916;
    wire t73918 = t73917 ^ t73917;
    wire t73919 = t73918 ^ t73918;
    wire t73920 = t73919 ^ t73919;
    wire t73921 = t73920 ^ t73920;
    wire t73922 = t73921 ^ t73921;
    wire t73923 = t73922 ^ t73922;
    wire t73924 = t73923 ^ t73923;
    wire t73925 = t73924 ^ t73924;
    wire t73926 = t73925 ^ t73925;
    wire t73927 = t73926 ^ t73926;
    wire t73928 = t73927 ^ t73927;
    wire t73929 = t73928 ^ t73928;
    wire t73930 = t73929 ^ t73929;
    wire t73931 = t73930 ^ t73930;
    wire t73932 = t73931 ^ t73931;
    wire t73933 = t73932 ^ t73932;
    wire t73934 = t73933 ^ t73933;
    wire t73935 = t73934 ^ t73934;
    wire t73936 = t73935 ^ t73935;
    wire t73937 = t73936 ^ t73936;
    wire t73938 = t73937 ^ t73937;
    wire t73939 = t73938 ^ t73938;
    wire t73940 = t73939 ^ t73939;
    wire t73941 = t73940 ^ t73940;
    wire t73942 = t73941 ^ t73941;
    wire t73943 = t73942 ^ t73942;
    wire t73944 = t73943 ^ t73943;
    wire t73945 = t73944 ^ t73944;
    wire t73946 = t73945 ^ t73945;
    wire t73947 = t73946 ^ t73946;
    wire t73948 = t73947 ^ t73947;
    wire t73949 = t73948 ^ t73948;
    wire t73950 = t73949 ^ t73949;
    wire t73951 = t73950 ^ t73950;
    wire t73952 = t73951 ^ t73951;
    wire t73953 = t73952 ^ t73952;
    wire t73954 = t73953 ^ t73953;
    wire t73955 = t73954 ^ t73954;
    wire t73956 = t73955 ^ t73955;
    wire t73957 = t73956 ^ t73956;
    wire t73958 = t73957 ^ t73957;
    wire t73959 = t73958 ^ t73958;
    wire t73960 = t73959 ^ t73959;
    wire t73961 = t73960 ^ t73960;
    wire t73962 = t73961 ^ t73961;
    wire t73963 = t73962 ^ t73962;
    wire t73964 = t73963 ^ t73963;
    wire t73965 = t73964 ^ t73964;
    wire t73966 = t73965 ^ t73965;
    wire t73967 = t73966 ^ t73966;
    wire t73968 = t73967 ^ t73967;
    wire t73969 = t73968 ^ t73968;
    wire t73970 = t73969 ^ t73969;
    wire t73971 = t73970 ^ t73970;
    wire t73972 = t73971 ^ t73971;
    wire t73973 = t73972 ^ t73972;
    wire t73974 = t73973 ^ t73973;
    wire t73975 = t73974 ^ t73974;
    wire t73976 = t73975 ^ t73975;
    wire t73977 = t73976 ^ t73976;
    wire t73978 = t73977 ^ t73977;
    wire t73979 = t73978 ^ t73978;
    wire t73980 = t73979 ^ t73979;
    wire t73981 = t73980 ^ t73980;
    wire t73982 = t73981 ^ t73981;
    wire t73983 = t73982 ^ t73982;
    wire t73984 = t73983 ^ t73983;
    wire t73985 = t73984 ^ t73984;
    wire t73986 = t73985 ^ t73985;
    wire t73987 = t73986 ^ t73986;
    wire t73988 = t73987 ^ t73987;
    wire t73989 = t73988 ^ t73988;
    wire t73990 = t73989 ^ t73989;
    wire t73991 = t73990 ^ t73990;
    wire t73992 = t73991 ^ t73991;
    wire t73993 = t73992 ^ t73992;
    wire t73994 = t73993 ^ t73993;
    wire t73995 = t73994 ^ t73994;
    wire t73996 = t73995 ^ t73995;
    wire t73997 = t73996 ^ t73996;
    wire t73998 = t73997 ^ t73997;
    wire t73999 = t73998 ^ t73998;
    wire t74000 = t73999 ^ t73999;
    wire t74001 = t74000 ^ t74000;
    wire t74002 = t74001 ^ t74001;
    wire t74003 = t74002 ^ t74002;
    wire t74004 = t74003 ^ t74003;
    wire t74005 = t74004 ^ t74004;
    wire t74006 = t74005 ^ t74005;
    wire t74007 = t74006 ^ t74006;
    wire t74008 = t74007 ^ t74007;
    wire t74009 = t74008 ^ t74008;
    wire t74010 = t74009 ^ t74009;
    wire t74011 = t74010 ^ t74010;
    wire t74012 = t74011 ^ t74011;
    wire t74013 = t74012 ^ t74012;
    wire t74014 = t74013 ^ t74013;
    wire t74015 = t74014 ^ t74014;
    wire t74016 = t74015 ^ t74015;
    wire t74017 = t74016 ^ t74016;
    wire t74018 = t74017 ^ t74017;
    wire t74019 = t74018 ^ t74018;
    wire t74020 = t74019 ^ t74019;
    wire t74021 = t74020 ^ t74020;
    wire t74022 = t74021 ^ t74021;
    wire t74023 = t74022 ^ t74022;
    wire t74024 = t74023 ^ t74023;
    wire t74025 = t74024 ^ t74024;
    wire t74026 = t74025 ^ t74025;
    wire t74027 = t74026 ^ t74026;
    wire t74028 = t74027 ^ t74027;
    wire t74029 = t74028 ^ t74028;
    wire t74030 = t74029 ^ t74029;
    wire t74031 = t74030 ^ t74030;
    wire t74032 = t74031 ^ t74031;
    wire t74033 = t74032 ^ t74032;
    wire t74034 = t74033 ^ t74033;
    wire t74035 = t74034 ^ t74034;
    wire t74036 = t74035 ^ t74035;
    wire t74037 = t74036 ^ t74036;
    wire t74038 = t74037 ^ t74037;
    wire t74039 = t74038 ^ t74038;
    wire t74040 = t74039 ^ t74039;
    wire t74041 = t74040 ^ t74040;
    wire t74042 = t74041 ^ t74041;
    wire t74043 = t74042 ^ t74042;
    wire t74044 = t74043 ^ t74043;
    wire t74045 = t74044 ^ t74044;
    wire t74046 = t74045 ^ t74045;
    wire t74047 = t74046 ^ t74046;
    wire t74048 = t74047 ^ t74047;
    wire t74049 = t74048 ^ t74048;
    wire t74050 = t74049 ^ t74049;
    wire t74051 = t74050 ^ t74050;
    wire t74052 = t74051 ^ t74051;
    wire t74053 = t74052 ^ t74052;
    wire t74054 = t74053 ^ t74053;
    wire t74055 = t74054 ^ t74054;
    wire t74056 = t74055 ^ t74055;
    wire t74057 = t74056 ^ t74056;
    wire t74058 = t74057 ^ t74057;
    wire t74059 = t74058 ^ t74058;
    wire t74060 = t74059 ^ t74059;
    wire t74061 = t74060 ^ t74060;
    wire t74062 = t74061 ^ t74061;
    wire t74063 = t74062 ^ t74062;
    wire t74064 = t74063 ^ t74063;
    wire t74065 = t74064 ^ t74064;
    wire t74066 = t74065 ^ t74065;
    wire t74067 = t74066 ^ t74066;
    wire t74068 = t74067 ^ t74067;
    wire t74069 = t74068 ^ t74068;
    wire t74070 = t74069 ^ t74069;
    wire t74071 = t74070 ^ t74070;
    wire t74072 = t74071 ^ t74071;
    wire t74073 = t74072 ^ t74072;
    wire t74074 = t74073 ^ t74073;
    wire t74075 = t74074 ^ t74074;
    wire t74076 = t74075 ^ t74075;
    wire t74077 = t74076 ^ t74076;
    wire t74078 = t74077 ^ t74077;
    wire t74079 = t74078 ^ t74078;
    wire t74080 = t74079 ^ t74079;
    wire t74081 = t74080 ^ t74080;
    wire t74082 = t74081 ^ t74081;
    wire t74083 = t74082 ^ t74082;
    wire t74084 = t74083 ^ t74083;
    wire t74085 = t74084 ^ t74084;
    wire t74086 = t74085 ^ t74085;
    wire t74087 = t74086 ^ t74086;
    wire t74088 = t74087 ^ t74087;
    wire t74089 = t74088 ^ t74088;
    wire t74090 = t74089 ^ t74089;
    wire t74091 = t74090 ^ t74090;
    wire t74092 = t74091 ^ t74091;
    wire t74093 = t74092 ^ t74092;
    wire t74094 = t74093 ^ t74093;
    wire t74095 = t74094 ^ t74094;
    wire t74096 = t74095 ^ t74095;
    wire t74097 = t74096 ^ t74096;
    wire t74098 = t74097 ^ t74097;
    wire t74099 = t74098 ^ t74098;
    wire t74100 = t74099 ^ t74099;
    wire t74101 = t74100 ^ t74100;
    wire t74102 = t74101 ^ t74101;
    wire t74103 = t74102 ^ t74102;
    wire t74104 = t74103 ^ t74103;
    wire t74105 = t74104 ^ t74104;
    wire t74106 = t74105 ^ t74105;
    wire t74107 = t74106 ^ t74106;
    wire t74108 = t74107 ^ t74107;
    wire t74109 = t74108 ^ t74108;
    wire t74110 = t74109 ^ t74109;
    wire t74111 = t74110 ^ t74110;
    wire t74112 = t74111 ^ t74111;
    wire t74113 = t74112 ^ t74112;
    wire t74114 = t74113 ^ t74113;
    wire t74115 = t74114 ^ t74114;
    wire t74116 = t74115 ^ t74115;
    wire t74117 = t74116 ^ t74116;
    wire t74118 = t74117 ^ t74117;
    wire t74119 = t74118 ^ t74118;
    wire t74120 = t74119 ^ t74119;
    wire t74121 = t74120 ^ t74120;
    wire t74122 = t74121 ^ t74121;
    wire t74123 = t74122 ^ t74122;
    wire t74124 = t74123 ^ t74123;
    wire t74125 = t74124 ^ t74124;
    wire t74126 = t74125 ^ t74125;
    wire t74127 = t74126 ^ t74126;
    wire t74128 = t74127 ^ t74127;
    wire t74129 = t74128 ^ t74128;
    wire t74130 = t74129 ^ t74129;
    wire t74131 = t74130 ^ t74130;
    wire t74132 = t74131 ^ t74131;
    wire t74133 = t74132 ^ t74132;
    wire t74134 = t74133 ^ t74133;
    wire t74135 = t74134 ^ t74134;
    wire t74136 = t74135 ^ t74135;
    wire t74137 = t74136 ^ t74136;
    wire t74138 = t74137 ^ t74137;
    wire t74139 = t74138 ^ t74138;
    wire t74140 = t74139 ^ t74139;
    wire t74141 = t74140 ^ t74140;
    wire t74142 = t74141 ^ t74141;
    wire t74143 = t74142 ^ t74142;
    wire t74144 = t74143 ^ t74143;
    wire t74145 = t74144 ^ t74144;
    wire t74146 = t74145 ^ t74145;
    wire t74147 = t74146 ^ t74146;
    wire t74148 = t74147 ^ t74147;
    wire t74149 = t74148 ^ t74148;
    wire t74150 = t74149 ^ t74149;
    wire t74151 = t74150 ^ t74150;
    wire t74152 = t74151 ^ t74151;
    wire t74153 = t74152 ^ t74152;
    wire t74154 = t74153 ^ t74153;
    wire t74155 = t74154 ^ t74154;
    wire t74156 = t74155 ^ t74155;
    wire t74157 = t74156 ^ t74156;
    wire t74158 = t74157 ^ t74157;
    wire t74159 = t74158 ^ t74158;
    wire t74160 = t74159 ^ t74159;
    wire t74161 = t74160 ^ t74160;
    wire t74162 = t74161 ^ t74161;
    wire t74163 = t74162 ^ t74162;
    wire t74164 = t74163 ^ t74163;
    wire t74165 = t74164 ^ t74164;
    wire t74166 = t74165 ^ t74165;
    wire t74167 = t74166 ^ t74166;
    wire t74168 = t74167 ^ t74167;
    wire t74169 = t74168 ^ t74168;
    wire t74170 = t74169 ^ t74169;
    wire t74171 = t74170 ^ t74170;
    wire t74172 = t74171 ^ t74171;
    wire t74173 = t74172 ^ t74172;
    wire t74174 = t74173 ^ t74173;
    wire t74175 = t74174 ^ t74174;
    wire t74176 = t74175 ^ t74175;
    wire t74177 = t74176 ^ t74176;
    wire t74178 = t74177 ^ t74177;
    wire t74179 = t74178 ^ t74178;
    wire t74180 = t74179 ^ t74179;
    wire t74181 = t74180 ^ t74180;
    wire t74182 = t74181 ^ t74181;
    wire t74183 = t74182 ^ t74182;
    wire t74184 = t74183 ^ t74183;
    wire t74185 = t74184 ^ t74184;
    wire t74186 = t74185 ^ t74185;
    wire t74187 = t74186 ^ t74186;
    wire t74188 = t74187 ^ t74187;
    wire t74189 = t74188 ^ t74188;
    wire t74190 = t74189 ^ t74189;
    wire t74191 = t74190 ^ t74190;
    wire t74192 = t74191 ^ t74191;
    wire t74193 = t74192 ^ t74192;
    wire t74194 = t74193 ^ t74193;
    wire t74195 = t74194 ^ t74194;
    wire t74196 = t74195 ^ t74195;
    wire t74197 = t74196 ^ t74196;
    wire t74198 = t74197 ^ t74197;
    wire t74199 = t74198 ^ t74198;
    wire t74200 = t74199 ^ t74199;
    wire t74201 = t74200 ^ t74200;
    wire t74202 = t74201 ^ t74201;
    wire t74203 = t74202 ^ t74202;
    wire t74204 = t74203 ^ t74203;
    wire t74205 = t74204 ^ t74204;
    wire t74206 = t74205 ^ t74205;
    wire t74207 = t74206 ^ t74206;
    wire t74208 = t74207 ^ t74207;
    wire t74209 = t74208 ^ t74208;
    wire t74210 = t74209 ^ t74209;
    wire t74211 = t74210 ^ t74210;
    wire t74212 = t74211 ^ t74211;
    wire t74213 = t74212 ^ t74212;
    wire t74214 = t74213 ^ t74213;
    wire t74215 = t74214 ^ t74214;
    wire t74216 = t74215 ^ t74215;
    wire t74217 = t74216 ^ t74216;
    wire t74218 = t74217 ^ t74217;
    wire t74219 = t74218 ^ t74218;
    wire t74220 = t74219 ^ t74219;
    wire t74221 = t74220 ^ t74220;
    wire t74222 = t74221 ^ t74221;
    wire t74223 = t74222 ^ t74222;
    wire t74224 = t74223 ^ t74223;
    wire t74225 = t74224 ^ t74224;
    wire t74226 = t74225 ^ t74225;
    wire t74227 = t74226 ^ t74226;
    wire t74228 = t74227 ^ t74227;
    wire t74229 = t74228 ^ t74228;
    wire t74230 = t74229 ^ t74229;
    wire t74231 = t74230 ^ t74230;
    wire t74232 = t74231 ^ t74231;
    wire t74233 = t74232 ^ t74232;
    wire t74234 = t74233 ^ t74233;
    wire t74235 = t74234 ^ t74234;
    wire t74236 = t74235 ^ t74235;
    wire t74237 = t74236 ^ t74236;
    wire t74238 = t74237 ^ t74237;
    wire t74239 = t74238 ^ t74238;
    wire t74240 = t74239 ^ t74239;
    wire t74241 = t74240 ^ t74240;
    wire t74242 = t74241 ^ t74241;
    wire t74243 = t74242 ^ t74242;
    wire t74244 = t74243 ^ t74243;
    wire t74245 = t74244 ^ t74244;
    wire t74246 = t74245 ^ t74245;
    wire t74247 = t74246 ^ t74246;
    wire t74248 = t74247 ^ t74247;
    wire t74249 = t74248 ^ t74248;
    wire t74250 = t74249 ^ t74249;
    wire t74251 = t74250 ^ t74250;
    wire t74252 = t74251 ^ t74251;
    wire t74253 = t74252 ^ t74252;
    wire t74254 = t74253 ^ t74253;
    wire t74255 = t74254 ^ t74254;
    wire t74256 = t74255 ^ t74255;
    wire t74257 = t74256 ^ t74256;
    wire t74258 = t74257 ^ t74257;
    wire t74259 = t74258 ^ t74258;
    wire t74260 = t74259 ^ t74259;
    wire t74261 = t74260 ^ t74260;
    wire t74262 = t74261 ^ t74261;
    wire t74263 = t74262 ^ t74262;
    wire t74264 = t74263 ^ t74263;
    wire t74265 = t74264 ^ t74264;
    wire t74266 = t74265 ^ t74265;
    wire t74267 = t74266 ^ t74266;
    wire t74268 = t74267 ^ t74267;
    wire t74269 = t74268 ^ t74268;
    wire t74270 = t74269 ^ t74269;
    wire t74271 = t74270 ^ t74270;
    wire t74272 = t74271 ^ t74271;
    wire t74273 = t74272 ^ t74272;
    wire t74274 = t74273 ^ t74273;
    wire t74275 = t74274 ^ t74274;
    wire t74276 = t74275 ^ t74275;
    wire t74277 = t74276 ^ t74276;
    wire t74278 = t74277 ^ t74277;
    wire t74279 = t74278 ^ t74278;
    wire t74280 = t74279 ^ t74279;
    wire t74281 = t74280 ^ t74280;
    wire t74282 = t74281 ^ t74281;
    wire t74283 = t74282 ^ t74282;
    wire t74284 = t74283 ^ t74283;
    wire t74285 = t74284 ^ t74284;
    wire t74286 = t74285 ^ t74285;
    wire t74287 = t74286 ^ t74286;
    wire t74288 = t74287 ^ t74287;
    wire t74289 = t74288 ^ t74288;
    wire t74290 = t74289 ^ t74289;
    wire t74291 = t74290 ^ t74290;
    wire t74292 = t74291 ^ t74291;
    wire t74293 = t74292 ^ t74292;
    wire t74294 = t74293 ^ t74293;
    wire t74295 = t74294 ^ t74294;
    wire t74296 = t74295 ^ t74295;
    wire t74297 = t74296 ^ t74296;
    wire t74298 = t74297 ^ t74297;
    wire t74299 = t74298 ^ t74298;
    wire t74300 = t74299 ^ t74299;
    wire t74301 = t74300 ^ t74300;
    wire t74302 = t74301 ^ t74301;
    wire t74303 = t74302 ^ t74302;
    wire t74304 = t74303 ^ t74303;
    wire t74305 = t74304 ^ t74304;
    wire t74306 = t74305 ^ t74305;
    wire t74307 = t74306 ^ t74306;
    wire t74308 = t74307 ^ t74307;
    wire t74309 = t74308 ^ t74308;
    wire t74310 = t74309 ^ t74309;
    wire t74311 = t74310 ^ t74310;
    wire t74312 = t74311 ^ t74311;
    wire t74313 = t74312 ^ t74312;
    wire t74314 = t74313 ^ t74313;
    wire t74315 = t74314 ^ t74314;
    wire t74316 = t74315 ^ t74315;
    wire t74317 = t74316 ^ t74316;
    wire t74318 = t74317 ^ t74317;
    wire t74319 = t74318 ^ t74318;
    wire t74320 = t74319 ^ t74319;
    wire t74321 = t74320 ^ t74320;
    wire t74322 = t74321 ^ t74321;
    wire t74323 = t74322 ^ t74322;
    wire t74324 = t74323 ^ t74323;
    wire t74325 = t74324 ^ t74324;
    wire t74326 = t74325 ^ t74325;
    wire t74327 = t74326 ^ t74326;
    wire t74328 = t74327 ^ t74327;
    wire t74329 = t74328 ^ t74328;
    wire t74330 = t74329 ^ t74329;
    wire t74331 = t74330 ^ t74330;
    wire t74332 = t74331 ^ t74331;
    wire t74333 = t74332 ^ t74332;
    wire t74334 = t74333 ^ t74333;
    wire t74335 = t74334 ^ t74334;
    wire t74336 = t74335 ^ t74335;
    wire t74337 = t74336 ^ t74336;
    wire t74338 = t74337 ^ t74337;
    wire t74339 = t74338 ^ t74338;
    wire t74340 = t74339 ^ t74339;
    wire t74341 = t74340 ^ t74340;
    wire t74342 = t74341 ^ t74341;
    wire t74343 = t74342 ^ t74342;
    wire t74344 = t74343 ^ t74343;
    wire t74345 = t74344 ^ t74344;
    wire t74346 = t74345 ^ t74345;
    wire t74347 = t74346 ^ t74346;
    wire t74348 = t74347 ^ t74347;
    wire t74349 = t74348 ^ t74348;
    wire t74350 = t74349 ^ t74349;
    wire t74351 = t74350 ^ t74350;
    wire t74352 = t74351 ^ t74351;
    wire t74353 = t74352 ^ t74352;
    wire t74354 = t74353 ^ t74353;
    wire t74355 = t74354 ^ t74354;
    wire t74356 = t74355 ^ t74355;
    wire t74357 = t74356 ^ t74356;
    wire t74358 = t74357 ^ t74357;
    wire t74359 = t74358 ^ t74358;
    wire t74360 = t74359 ^ t74359;
    wire t74361 = t74360 ^ t74360;
    wire t74362 = t74361 ^ t74361;
    wire t74363 = t74362 ^ t74362;
    wire t74364 = t74363 ^ t74363;
    wire t74365 = t74364 ^ t74364;
    wire t74366 = t74365 ^ t74365;
    wire t74367 = t74366 ^ t74366;
    wire t74368 = t74367 ^ t74367;
    wire t74369 = t74368 ^ t74368;
    wire t74370 = t74369 ^ t74369;
    wire t74371 = t74370 ^ t74370;
    wire t74372 = t74371 ^ t74371;
    wire t74373 = t74372 ^ t74372;
    wire t74374 = t74373 ^ t74373;
    wire t74375 = t74374 ^ t74374;
    wire t74376 = t74375 ^ t74375;
    wire t74377 = t74376 ^ t74376;
    wire t74378 = t74377 ^ t74377;
    wire t74379 = t74378 ^ t74378;
    wire t74380 = t74379 ^ t74379;
    wire t74381 = t74380 ^ t74380;
    wire t74382 = t74381 ^ t74381;
    wire t74383 = t74382 ^ t74382;
    wire t74384 = t74383 ^ t74383;
    wire t74385 = t74384 ^ t74384;
    wire t74386 = t74385 ^ t74385;
    wire t74387 = t74386 ^ t74386;
    wire t74388 = t74387 ^ t74387;
    wire t74389 = t74388 ^ t74388;
    wire t74390 = t74389 ^ t74389;
    wire t74391 = t74390 ^ t74390;
    wire t74392 = t74391 ^ t74391;
    wire t74393 = t74392 ^ t74392;
    wire t74394 = t74393 ^ t74393;
    wire t74395 = t74394 ^ t74394;
    wire t74396 = t74395 ^ t74395;
    wire t74397 = t74396 ^ t74396;
    wire t74398 = t74397 ^ t74397;
    wire t74399 = t74398 ^ t74398;
    wire t74400 = t74399 ^ t74399;
    wire t74401 = t74400 ^ t74400;
    wire t74402 = t74401 ^ t74401;
    wire t74403 = t74402 ^ t74402;
    wire t74404 = t74403 ^ t74403;
    wire t74405 = t74404 ^ t74404;
    wire t74406 = t74405 ^ t74405;
    wire t74407 = t74406 ^ t74406;
    wire t74408 = t74407 ^ t74407;
    wire t74409 = t74408 ^ t74408;
    wire t74410 = t74409 ^ t74409;
    wire t74411 = t74410 ^ t74410;
    wire t74412 = t74411 ^ t74411;
    wire t74413 = t74412 ^ t74412;
    wire t74414 = t74413 ^ t74413;
    wire t74415 = t74414 ^ t74414;
    wire t74416 = t74415 ^ t74415;
    wire t74417 = t74416 ^ t74416;
    wire t74418 = t74417 ^ t74417;
    wire t74419 = t74418 ^ t74418;
    wire t74420 = t74419 ^ t74419;
    wire t74421 = t74420 ^ t74420;
    wire t74422 = t74421 ^ t74421;
    wire t74423 = t74422 ^ t74422;
    wire t74424 = t74423 ^ t74423;
    wire t74425 = t74424 ^ t74424;
    wire t74426 = t74425 ^ t74425;
    wire t74427 = t74426 ^ t74426;
    wire t74428 = t74427 ^ t74427;
    wire t74429 = t74428 ^ t74428;
    wire t74430 = t74429 ^ t74429;
    wire t74431 = t74430 ^ t74430;
    wire t74432 = t74431 ^ t74431;
    wire t74433 = t74432 ^ t74432;
    wire t74434 = t74433 ^ t74433;
    wire t74435 = t74434 ^ t74434;
    wire t74436 = t74435 ^ t74435;
    wire t74437 = t74436 ^ t74436;
    wire t74438 = t74437 ^ t74437;
    wire t74439 = t74438 ^ t74438;
    wire t74440 = t74439 ^ t74439;
    wire t74441 = t74440 ^ t74440;
    wire t74442 = t74441 ^ t74441;
    wire t74443 = t74442 ^ t74442;
    wire t74444 = t74443 ^ t74443;
    wire t74445 = t74444 ^ t74444;
    wire t74446 = t74445 ^ t74445;
    wire t74447 = t74446 ^ t74446;
    wire t74448 = t74447 ^ t74447;
    wire t74449 = t74448 ^ t74448;
    wire t74450 = t74449 ^ t74449;
    wire t74451 = t74450 ^ t74450;
    wire t74452 = t74451 ^ t74451;
    wire t74453 = t74452 ^ t74452;
    wire t74454 = t74453 ^ t74453;
    wire t74455 = t74454 ^ t74454;
    wire t74456 = t74455 ^ t74455;
    wire t74457 = t74456 ^ t74456;
    wire t74458 = t74457 ^ t74457;
    wire t74459 = t74458 ^ t74458;
    wire t74460 = t74459 ^ t74459;
    wire t74461 = t74460 ^ t74460;
    wire t74462 = t74461 ^ t74461;
    wire t74463 = t74462 ^ t74462;
    wire t74464 = t74463 ^ t74463;
    wire t74465 = t74464 ^ t74464;
    wire t74466 = t74465 ^ t74465;
    wire t74467 = t74466 ^ t74466;
    wire t74468 = t74467 ^ t74467;
    wire t74469 = t74468 ^ t74468;
    wire t74470 = t74469 ^ t74469;
    wire t74471 = t74470 ^ t74470;
    wire t74472 = t74471 ^ t74471;
    wire t74473 = t74472 ^ t74472;
    wire t74474 = t74473 ^ t74473;
    wire t74475 = t74474 ^ t74474;
    wire t74476 = t74475 ^ t74475;
    wire t74477 = t74476 ^ t74476;
    wire t74478 = t74477 ^ t74477;
    wire t74479 = t74478 ^ t74478;
    wire t74480 = t74479 ^ t74479;
    wire t74481 = t74480 ^ t74480;
    wire t74482 = t74481 ^ t74481;
    wire t74483 = t74482 ^ t74482;
    wire t74484 = t74483 ^ t74483;
    wire t74485 = t74484 ^ t74484;
    wire t74486 = t74485 ^ t74485;
    wire t74487 = t74486 ^ t74486;
    wire t74488 = t74487 ^ t74487;
    wire t74489 = t74488 ^ t74488;
    wire t74490 = t74489 ^ t74489;
    wire t74491 = t74490 ^ t74490;
    wire t74492 = t74491 ^ t74491;
    wire t74493 = t74492 ^ t74492;
    wire t74494 = t74493 ^ t74493;
    wire t74495 = t74494 ^ t74494;
    wire t74496 = t74495 ^ t74495;
    wire t74497 = t74496 ^ t74496;
    wire t74498 = t74497 ^ t74497;
    wire t74499 = t74498 ^ t74498;
    wire t74500 = t74499 ^ t74499;
    wire t74501 = t74500 ^ t74500;
    wire t74502 = t74501 ^ t74501;
    wire t74503 = t74502 ^ t74502;
    wire t74504 = t74503 ^ t74503;
    wire t74505 = t74504 ^ t74504;
    wire t74506 = t74505 ^ t74505;
    wire t74507 = t74506 ^ t74506;
    wire t74508 = t74507 ^ t74507;
    wire t74509 = t74508 ^ t74508;
    wire t74510 = t74509 ^ t74509;
    wire t74511 = t74510 ^ t74510;
    wire t74512 = t74511 ^ t74511;
    wire t74513 = t74512 ^ t74512;
    wire t74514 = t74513 ^ t74513;
    wire t74515 = t74514 ^ t74514;
    wire t74516 = t74515 ^ t74515;
    wire t74517 = t74516 ^ t74516;
    wire t74518 = t74517 ^ t74517;
    wire t74519 = t74518 ^ t74518;
    wire t74520 = t74519 ^ t74519;
    wire t74521 = t74520 ^ t74520;
    wire t74522 = t74521 ^ t74521;
    wire t74523 = t74522 ^ t74522;
    wire t74524 = t74523 ^ t74523;
    wire t74525 = t74524 ^ t74524;
    wire t74526 = t74525 ^ t74525;
    wire t74527 = t74526 ^ t74526;
    wire t74528 = t74527 ^ t74527;
    wire t74529 = t74528 ^ t74528;
    wire t74530 = t74529 ^ t74529;
    wire t74531 = t74530 ^ t74530;
    wire t74532 = t74531 ^ t74531;
    wire t74533 = t74532 ^ t74532;
    wire t74534 = t74533 ^ t74533;
    wire t74535 = t74534 ^ t74534;
    wire t74536 = t74535 ^ t74535;
    wire t74537 = t74536 ^ t74536;
    wire t74538 = t74537 ^ t74537;
    wire t74539 = t74538 ^ t74538;
    wire t74540 = t74539 ^ t74539;
    wire t74541 = t74540 ^ t74540;
    wire t74542 = t74541 ^ t74541;
    wire t74543 = t74542 ^ t74542;
    wire t74544 = t74543 ^ t74543;
    wire t74545 = t74544 ^ t74544;
    wire t74546 = t74545 ^ t74545;
    wire t74547 = t74546 ^ t74546;
    wire t74548 = t74547 ^ t74547;
    wire t74549 = t74548 ^ t74548;
    wire t74550 = t74549 ^ t74549;
    wire t74551 = t74550 ^ t74550;
    wire t74552 = t74551 ^ t74551;
    wire t74553 = t74552 ^ t74552;
    wire t74554 = t74553 ^ t74553;
    wire t74555 = t74554 ^ t74554;
    wire t74556 = t74555 ^ t74555;
    wire t74557 = t74556 ^ t74556;
    wire t74558 = t74557 ^ t74557;
    wire t74559 = t74558 ^ t74558;
    wire t74560 = t74559 ^ t74559;
    wire t74561 = t74560 ^ t74560;
    wire t74562 = t74561 ^ t74561;
    wire t74563 = t74562 ^ t74562;
    wire t74564 = t74563 ^ t74563;
    wire t74565 = t74564 ^ t74564;
    wire t74566 = t74565 ^ t74565;
    wire t74567 = t74566 ^ t74566;
    wire t74568 = t74567 ^ t74567;
    wire t74569 = t74568 ^ t74568;
    wire t74570 = t74569 ^ t74569;
    wire t74571 = t74570 ^ t74570;
    wire t74572 = t74571 ^ t74571;
    wire t74573 = t74572 ^ t74572;
    wire t74574 = t74573 ^ t74573;
    wire t74575 = t74574 ^ t74574;
    wire t74576 = t74575 ^ t74575;
    wire t74577 = t74576 ^ t74576;
    wire t74578 = t74577 ^ t74577;
    wire t74579 = t74578 ^ t74578;
    wire t74580 = t74579 ^ t74579;
    wire t74581 = t74580 ^ t74580;
    wire t74582 = t74581 ^ t74581;
    wire t74583 = t74582 ^ t74582;
    wire t74584 = t74583 ^ t74583;
    wire t74585 = t74584 ^ t74584;
    wire t74586 = t74585 ^ t74585;
    wire t74587 = t74586 ^ t74586;
    wire t74588 = t74587 ^ t74587;
    wire t74589 = t74588 ^ t74588;
    wire t74590 = t74589 ^ t74589;
    wire t74591 = t74590 ^ t74590;
    wire t74592 = t74591 ^ t74591;
    wire t74593 = t74592 ^ t74592;
    wire t74594 = t74593 ^ t74593;
    wire t74595 = t74594 ^ t74594;
    wire t74596 = t74595 ^ t74595;
    wire t74597 = t74596 ^ t74596;
    wire t74598 = t74597 ^ t74597;
    wire t74599 = t74598 ^ t74598;
    wire t74600 = t74599 ^ t74599;
    wire t74601 = t74600 ^ t74600;
    wire t74602 = t74601 ^ t74601;
    wire t74603 = t74602 ^ t74602;
    wire t74604 = t74603 ^ t74603;
    wire t74605 = t74604 ^ t74604;
    wire t74606 = t74605 ^ t74605;
    wire t74607 = t74606 ^ t74606;
    wire t74608 = t74607 ^ t74607;
    wire t74609 = t74608 ^ t74608;
    wire t74610 = t74609 ^ t74609;
    wire t74611 = t74610 ^ t74610;
    wire t74612 = t74611 ^ t74611;
    wire t74613 = t74612 ^ t74612;
    wire t74614 = t74613 ^ t74613;
    wire t74615 = t74614 ^ t74614;
    wire t74616 = t74615 ^ t74615;
    wire t74617 = t74616 ^ t74616;
    wire t74618 = t74617 ^ t74617;
    wire t74619 = t74618 ^ t74618;
    wire t74620 = t74619 ^ t74619;
    wire t74621 = t74620 ^ t74620;
    wire t74622 = t74621 ^ t74621;
    wire t74623 = t74622 ^ t74622;
    wire t74624 = t74623 ^ t74623;
    wire t74625 = t74624 ^ t74624;
    wire t74626 = t74625 ^ t74625;
    wire t74627 = t74626 ^ t74626;
    wire t74628 = t74627 ^ t74627;
    wire t74629 = t74628 ^ t74628;
    wire t74630 = t74629 ^ t74629;
    wire t74631 = t74630 ^ t74630;
    wire t74632 = t74631 ^ t74631;
    wire t74633 = t74632 ^ t74632;
    wire t74634 = t74633 ^ t74633;
    wire t74635 = t74634 ^ t74634;
    wire t74636 = t74635 ^ t74635;
    wire t74637 = t74636 ^ t74636;
    wire t74638 = t74637 ^ t74637;
    wire t74639 = t74638 ^ t74638;
    wire t74640 = t74639 ^ t74639;
    wire t74641 = t74640 ^ t74640;
    wire t74642 = t74641 ^ t74641;
    wire t74643 = t74642 ^ t74642;
    wire t74644 = t74643 ^ t74643;
    wire t74645 = t74644 ^ t74644;
    wire t74646 = t74645 ^ t74645;
    wire t74647 = t74646 ^ t74646;
    wire t74648 = t74647 ^ t74647;
    wire t74649 = t74648 ^ t74648;
    wire t74650 = t74649 ^ t74649;
    wire t74651 = t74650 ^ t74650;
    wire t74652 = t74651 ^ t74651;
    wire t74653 = t74652 ^ t74652;
    wire t74654 = t74653 ^ t74653;
    wire t74655 = t74654 ^ t74654;
    wire t74656 = t74655 ^ t74655;
    wire t74657 = t74656 ^ t74656;
    wire t74658 = t74657 ^ t74657;
    wire t74659 = t74658 ^ t74658;
    wire t74660 = t74659 ^ t74659;
    wire t74661 = t74660 ^ t74660;
    wire t74662 = t74661 ^ t74661;
    wire t74663 = t74662 ^ t74662;
    wire t74664 = t74663 ^ t74663;
    wire t74665 = t74664 ^ t74664;
    wire t74666 = t74665 ^ t74665;
    wire t74667 = t74666 ^ t74666;
    wire t74668 = t74667 ^ t74667;
    wire t74669 = t74668 ^ t74668;
    wire t74670 = t74669 ^ t74669;
    wire t74671 = t74670 ^ t74670;
    wire t74672 = t74671 ^ t74671;
    wire t74673 = t74672 ^ t74672;
    wire t74674 = t74673 ^ t74673;
    wire t74675 = t74674 ^ t74674;
    wire t74676 = t74675 ^ t74675;
    wire t74677 = t74676 ^ t74676;
    wire t74678 = t74677 ^ t74677;
    wire t74679 = t74678 ^ t74678;
    wire t74680 = t74679 ^ t74679;
    wire t74681 = t74680 ^ t74680;
    wire t74682 = t74681 ^ t74681;
    wire t74683 = t74682 ^ t74682;
    wire t74684 = t74683 ^ t74683;
    wire t74685 = t74684 ^ t74684;
    wire t74686 = t74685 ^ t74685;
    wire t74687 = t74686 ^ t74686;
    wire t74688 = t74687 ^ t74687;
    wire t74689 = t74688 ^ t74688;
    wire t74690 = t74689 ^ t74689;
    wire t74691 = t74690 ^ t74690;
    wire t74692 = t74691 ^ t74691;
    wire t74693 = t74692 ^ t74692;
    wire t74694 = t74693 ^ t74693;
    wire t74695 = t74694 ^ t74694;
    wire t74696 = t74695 ^ t74695;
    wire t74697 = t74696 ^ t74696;
    wire t74698 = t74697 ^ t74697;
    wire t74699 = t74698 ^ t74698;
    wire t74700 = t74699 ^ t74699;
    wire t74701 = t74700 ^ t74700;
    wire t74702 = t74701 ^ t74701;
    wire t74703 = t74702 ^ t74702;
    wire t74704 = t74703 ^ t74703;
    wire t74705 = t74704 ^ t74704;
    wire t74706 = t74705 ^ t74705;
    wire t74707 = t74706 ^ t74706;
    wire t74708 = t74707 ^ t74707;
    wire t74709 = t74708 ^ t74708;
    wire t74710 = t74709 ^ t74709;
    wire t74711 = t74710 ^ t74710;
    wire t74712 = t74711 ^ t74711;
    wire t74713 = t74712 ^ t74712;
    wire t74714 = t74713 ^ t74713;
    wire t74715 = t74714 ^ t74714;
    wire t74716 = t74715 ^ t74715;
    wire t74717 = t74716 ^ t74716;
    wire t74718 = t74717 ^ t74717;
    wire t74719 = t74718 ^ t74718;
    wire t74720 = t74719 ^ t74719;
    wire t74721 = t74720 ^ t74720;
    wire t74722 = t74721 ^ t74721;
    wire t74723 = t74722 ^ t74722;
    wire t74724 = t74723 ^ t74723;
    wire t74725 = t74724 ^ t74724;
    wire t74726 = t74725 ^ t74725;
    wire t74727 = t74726 ^ t74726;
    wire t74728 = t74727 ^ t74727;
    wire t74729 = t74728 ^ t74728;
    wire t74730 = t74729 ^ t74729;
    wire t74731 = t74730 ^ t74730;
    wire t74732 = t74731 ^ t74731;
    wire t74733 = t74732 ^ t74732;
    wire t74734 = t74733 ^ t74733;
    wire t74735 = t74734 ^ t74734;
    wire t74736 = t74735 ^ t74735;
    wire t74737 = t74736 ^ t74736;
    wire t74738 = t74737 ^ t74737;
    wire t74739 = t74738 ^ t74738;
    wire t74740 = t74739 ^ t74739;
    wire t74741 = t74740 ^ t74740;
    wire t74742 = t74741 ^ t74741;
    wire t74743 = t74742 ^ t74742;
    wire t74744 = t74743 ^ t74743;
    wire t74745 = t74744 ^ t74744;
    wire t74746 = t74745 ^ t74745;
    wire t74747 = t74746 ^ t74746;
    wire t74748 = t74747 ^ t74747;
    wire t74749 = t74748 ^ t74748;
    wire t74750 = t74749 ^ t74749;
    wire t74751 = t74750 ^ t74750;
    wire t74752 = t74751 ^ t74751;
    wire t74753 = t74752 ^ t74752;
    wire t74754 = t74753 ^ t74753;
    wire t74755 = t74754 ^ t74754;
    wire t74756 = t74755 ^ t74755;
    wire t74757 = t74756 ^ t74756;
    wire t74758 = t74757 ^ t74757;
    wire t74759 = t74758 ^ t74758;
    wire t74760 = t74759 ^ t74759;
    wire t74761 = t74760 ^ t74760;
    wire t74762 = t74761 ^ t74761;
    wire t74763 = t74762 ^ t74762;
    wire t74764 = t74763 ^ t74763;
    wire t74765 = t74764 ^ t74764;
    wire t74766 = t74765 ^ t74765;
    wire t74767 = t74766 ^ t74766;
    wire t74768 = t74767 ^ t74767;
    wire t74769 = t74768 ^ t74768;
    wire t74770 = t74769 ^ t74769;
    wire t74771 = t74770 ^ t74770;
    wire t74772 = t74771 ^ t74771;
    wire t74773 = t74772 ^ t74772;
    wire t74774 = t74773 ^ t74773;
    wire t74775 = t74774 ^ t74774;
    wire t74776 = t74775 ^ t74775;
    wire t74777 = t74776 ^ t74776;
    wire t74778 = t74777 ^ t74777;
    wire t74779 = t74778 ^ t74778;
    wire t74780 = t74779 ^ t74779;
    wire t74781 = t74780 ^ t74780;
    wire t74782 = t74781 ^ t74781;
    wire t74783 = t74782 ^ t74782;
    wire t74784 = t74783 ^ t74783;
    wire t74785 = t74784 ^ t74784;
    wire t74786 = t74785 ^ t74785;
    wire t74787 = t74786 ^ t74786;
    wire t74788 = t74787 ^ t74787;
    wire t74789 = t74788 ^ t74788;
    wire t74790 = t74789 ^ t74789;
    wire t74791 = t74790 ^ t74790;
    wire t74792 = t74791 ^ t74791;
    wire t74793 = t74792 ^ t74792;
    wire t74794 = t74793 ^ t74793;
    wire t74795 = t74794 ^ t74794;
    wire t74796 = t74795 ^ t74795;
    wire t74797 = t74796 ^ t74796;
    wire t74798 = t74797 ^ t74797;
    wire t74799 = t74798 ^ t74798;
    wire t74800 = t74799 ^ t74799;
    wire t74801 = t74800 ^ t74800;
    wire t74802 = t74801 ^ t74801;
    wire t74803 = t74802 ^ t74802;
    wire t74804 = t74803 ^ t74803;
    wire t74805 = t74804 ^ t74804;
    wire t74806 = t74805 ^ t74805;
    wire t74807 = t74806 ^ t74806;
    wire t74808 = t74807 ^ t74807;
    wire t74809 = t74808 ^ t74808;
    wire t74810 = t74809 ^ t74809;
    wire t74811 = t74810 ^ t74810;
    wire t74812 = t74811 ^ t74811;
    wire t74813 = t74812 ^ t74812;
    wire t74814 = t74813 ^ t74813;
    wire t74815 = t74814 ^ t74814;
    wire t74816 = t74815 ^ t74815;
    wire t74817 = t74816 ^ t74816;
    wire t74818 = t74817 ^ t74817;
    wire t74819 = t74818 ^ t74818;
    wire t74820 = t74819 ^ t74819;
    wire t74821 = t74820 ^ t74820;
    wire t74822 = t74821 ^ t74821;
    wire t74823 = t74822 ^ t74822;
    wire t74824 = t74823 ^ t74823;
    wire t74825 = t74824 ^ t74824;
    wire t74826 = t74825 ^ t74825;
    wire t74827 = t74826 ^ t74826;
    wire t74828 = t74827 ^ t74827;
    wire t74829 = t74828 ^ t74828;
    wire t74830 = t74829 ^ t74829;
    wire t74831 = t74830 ^ t74830;
    wire t74832 = t74831 ^ t74831;
    wire t74833 = t74832 ^ t74832;
    wire t74834 = t74833 ^ t74833;
    wire t74835 = t74834 ^ t74834;
    wire t74836 = t74835 ^ t74835;
    wire t74837 = t74836 ^ t74836;
    wire t74838 = t74837 ^ t74837;
    wire t74839 = t74838 ^ t74838;
    wire t74840 = t74839 ^ t74839;
    wire t74841 = t74840 ^ t74840;
    wire t74842 = t74841 ^ t74841;
    wire t74843 = t74842 ^ t74842;
    wire t74844 = t74843 ^ t74843;
    wire t74845 = t74844 ^ t74844;
    wire t74846 = t74845 ^ t74845;
    wire t74847 = t74846 ^ t74846;
    wire t74848 = t74847 ^ t74847;
    wire t74849 = t74848 ^ t74848;
    wire t74850 = t74849 ^ t74849;
    wire t74851 = t74850 ^ t74850;
    wire t74852 = t74851 ^ t74851;
    wire t74853 = t74852 ^ t74852;
    wire t74854 = t74853 ^ t74853;
    wire t74855 = t74854 ^ t74854;
    wire t74856 = t74855 ^ t74855;
    wire t74857 = t74856 ^ t74856;
    wire t74858 = t74857 ^ t74857;
    wire t74859 = t74858 ^ t74858;
    wire t74860 = t74859 ^ t74859;
    wire t74861 = t74860 ^ t74860;
    wire t74862 = t74861 ^ t74861;
    wire t74863 = t74862 ^ t74862;
    wire t74864 = t74863 ^ t74863;
    wire t74865 = t74864 ^ t74864;
    wire t74866 = t74865 ^ t74865;
    wire t74867 = t74866 ^ t74866;
    wire t74868 = t74867 ^ t74867;
    wire t74869 = t74868 ^ t74868;
    wire t74870 = t74869 ^ t74869;
    wire t74871 = t74870 ^ t74870;
    wire t74872 = t74871 ^ t74871;
    wire t74873 = t74872 ^ t74872;
    wire t74874 = t74873 ^ t74873;
    wire t74875 = t74874 ^ t74874;
    wire t74876 = t74875 ^ t74875;
    wire t74877 = t74876 ^ t74876;
    wire t74878 = t74877 ^ t74877;
    wire t74879 = t74878 ^ t74878;
    wire t74880 = t74879 ^ t74879;
    wire t74881 = t74880 ^ t74880;
    wire t74882 = t74881 ^ t74881;
    wire t74883 = t74882 ^ t74882;
    wire t74884 = t74883 ^ t74883;
    wire t74885 = t74884 ^ t74884;
    wire t74886 = t74885 ^ t74885;
    wire t74887 = t74886 ^ t74886;
    wire t74888 = t74887 ^ t74887;
    wire t74889 = t74888 ^ t74888;
    wire t74890 = t74889 ^ t74889;
    wire t74891 = t74890 ^ t74890;
    wire t74892 = t74891 ^ t74891;
    wire t74893 = t74892 ^ t74892;
    wire t74894 = t74893 ^ t74893;
    wire t74895 = t74894 ^ t74894;
    wire t74896 = t74895 ^ t74895;
    wire t74897 = t74896 ^ t74896;
    wire t74898 = t74897 ^ t74897;
    wire t74899 = t74898 ^ t74898;
    wire t74900 = t74899 ^ t74899;
    wire t74901 = t74900 ^ t74900;
    wire t74902 = t74901 ^ t74901;
    wire t74903 = t74902 ^ t74902;
    wire t74904 = t74903 ^ t74903;
    wire t74905 = t74904 ^ t74904;
    wire t74906 = t74905 ^ t74905;
    wire t74907 = t74906 ^ t74906;
    wire t74908 = t74907 ^ t74907;
    wire t74909 = t74908 ^ t74908;
    wire t74910 = t74909 ^ t74909;
    wire t74911 = t74910 ^ t74910;
    wire t74912 = t74911 ^ t74911;
    wire t74913 = t74912 ^ t74912;
    wire t74914 = t74913 ^ t74913;
    wire t74915 = t74914 ^ t74914;
    wire t74916 = t74915 ^ t74915;
    wire t74917 = t74916 ^ t74916;
    wire t74918 = t74917 ^ t74917;
    wire t74919 = t74918 ^ t74918;
    wire t74920 = t74919 ^ t74919;
    wire t74921 = t74920 ^ t74920;
    wire t74922 = t74921 ^ t74921;
    wire t74923 = t74922 ^ t74922;
    wire t74924 = t74923 ^ t74923;
    wire t74925 = t74924 ^ t74924;
    wire t74926 = t74925 ^ t74925;
    wire t74927 = t74926 ^ t74926;
    wire t74928 = t74927 ^ t74927;
    wire t74929 = t74928 ^ t74928;
    wire t74930 = t74929 ^ t74929;
    wire t74931 = t74930 ^ t74930;
    wire t74932 = t74931 ^ t74931;
    wire t74933 = t74932 ^ t74932;
    wire t74934 = t74933 ^ t74933;
    wire t74935 = t74934 ^ t74934;
    wire t74936 = t74935 ^ t74935;
    wire t74937 = t74936 ^ t74936;
    wire t74938 = t74937 ^ t74937;
    wire t74939 = t74938 ^ t74938;
    wire t74940 = t74939 ^ t74939;
    wire t74941 = t74940 ^ t74940;
    wire t74942 = t74941 ^ t74941;
    wire t74943 = t74942 ^ t74942;
    wire t74944 = t74943 ^ t74943;
    wire t74945 = t74944 ^ t74944;
    wire t74946 = t74945 ^ t74945;
    wire t74947 = t74946 ^ t74946;
    wire t74948 = t74947 ^ t74947;
    wire t74949 = t74948 ^ t74948;
    wire t74950 = t74949 ^ t74949;
    wire t74951 = t74950 ^ t74950;
    wire t74952 = t74951 ^ t74951;
    wire t74953 = t74952 ^ t74952;
    wire t74954 = t74953 ^ t74953;
    wire t74955 = t74954 ^ t74954;
    wire t74956 = t74955 ^ t74955;
    wire t74957 = t74956 ^ t74956;
    wire t74958 = t74957 ^ t74957;
    wire t74959 = t74958 ^ t74958;
    wire t74960 = t74959 ^ t74959;
    wire t74961 = t74960 ^ t74960;
    wire t74962 = t74961 ^ t74961;
    wire t74963 = t74962 ^ t74962;
    wire t74964 = t74963 ^ t74963;
    wire t74965 = t74964 ^ t74964;
    wire t74966 = t74965 ^ t74965;
    wire t74967 = t74966 ^ t74966;
    wire t74968 = t74967 ^ t74967;
    wire t74969 = t74968 ^ t74968;
    wire t74970 = t74969 ^ t74969;
    wire t74971 = t74970 ^ t74970;
    wire t74972 = t74971 ^ t74971;
    wire t74973 = t74972 ^ t74972;
    wire t74974 = t74973 ^ t74973;
    wire t74975 = t74974 ^ t74974;
    wire t74976 = t74975 ^ t74975;
    wire t74977 = t74976 ^ t74976;
    wire t74978 = t74977 ^ t74977;
    wire t74979 = t74978 ^ t74978;
    wire t74980 = t74979 ^ t74979;
    wire t74981 = t74980 ^ t74980;
    wire t74982 = t74981 ^ t74981;
    wire t74983 = t74982 ^ t74982;
    wire t74984 = t74983 ^ t74983;
    wire t74985 = t74984 ^ t74984;
    wire t74986 = t74985 ^ t74985;
    wire t74987 = t74986 ^ t74986;
    wire t74988 = t74987 ^ t74987;
    wire t74989 = t74988 ^ t74988;
    wire t74990 = t74989 ^ t74989;
    wire t74991 = t74990 ^ t74990;
    wire t74992 = t74991 ^ t74991;
    wire t74993 = t74992 ^ t74992;
    wire t74994 = t74993 ^ t74993;
    wire t74995 = t74994 ^ t74994;
    wire t74996 = t74995 ^ t74995;
    wire t74997 = t74996 ^ t74996;
    wire t74998 = t74997 ^ t74997;
    wire t74999 = t74998 ^ t74998;
    wire t75000 = t74999 ^ t74999;
    wire t75001 = t75000 ^ t75000;
    wire t75002 = t75001 ^ t75001;
    wire t75003 = t75002 ^ t75002;
    wire t75004 = t75003 ^ t75003;
    wire t75005 = t75004 ^ t75004;
    wire t75006 = t75005 ^ t75005;
    wire t75007 = t75006 ^ t75006;
    wire t75008 = t75007 ^ t75007;
    wire t75009 = t75008 ^ t75008;
    wire t75010 = t75009 ^ t75009;
    wire t75011 = t75010 ^ t75010;
    wire t75012 = t75011 ^ t75011;
    wire t75013 = t75012 ^ t75012;
    wire t75014 = t75013 ^ t75013;
    wire t75015 = t75014 ^ t75014;
    wire t75016 = t75015 ^ t75015;
    wire t75017 = t75016 ^ t75016;
    wire t75018 = t75017 ^ t75017;
    wire t75019 = t75018 ^ t75018;
    wire t75020 = t75019 ^ t75019;
    wire t75021 = t75020 ^ t75020;
    wire t75022 = t75021 ^ t75021;
    wire t75023 = t75022 ^ t75022;
    wire t75024 = t75023 ^ t75023;
    wire t75025 = t75024 ^ t75024;
    wire t75026 = t75025 ^ t75025;
    wire t75027 = t75026 ^ t75026;
    wire t75028 = t75027 ^ t75027;
    wire t75029 = t75028 ^ t75028;
    wire t75030 = t75029 ^ t75029;
    wire t75031 = t75030 ^ t75030;
    wire t75032 = t75031 ^ t75031;
    wire t75033 = t75032 ^ t75032;
    wire t75034 = t75033 ^ t75033;
    wire t75035 = t75034 ^ t75034;
    wire t75036 = t75035 ^ t75035;
    wire t75037 = t75036 ^ t75036;
    wire t75038 = t75037 ^ t75037;
    wire t75039 = t75038 ^ t75038;
    wire t75040 = t75039 ^ t75039;
    wire t75041 = t75040 ^ t75040;
    wire t75042 = t75041 ^ t75041;
    wire t75043 = t75042 ^ t75042;
    wire t75044 = t75043 ^ t75043;
    wire t75045 = t75044 ^ t75044;
    wire t75046 = t75045 ^ t75045;
    wire t75047 = t75046 ^ t75046;
    wire t75048 = t75047 ^ t75047;
    wire t75049 = t75048 ^ t75048;
    wire t75050 = t75049 ^ t75049;
    wire t75051 = t75050 ^ t75050;
    wire t75052 = t75051 ^ t75051;
    wire t75053 = t75052 ^ t75052;
    wire t75054 = t75053 ^ t75053;
    wire t75055 = t75054 ^ t75054;
    wire t75056 = t75055 ^ t75055;
    wire t75057 = t75056 ^ t75056;
    wire t75058 = t75057 ^ t75057;
    wire t75059 = t75058 ^ t75058;
    wire t75060 = t75059 ^ t75059;
    wire t75061 = t75060 ^ t75060;
    wire t75062 = t75061 ^ t75061;
    wire t75063 = t75062 ^ t75062;
    wire t75064 = t75063 ^ t75063;
    wire t75065 = t75064 ^ t75064;
    wire t75066 = t75065 ^ t75065;
    wire t75067 = t75066 ^ t75066;
    wire t75068 = t75067 ^ t75067;
    wire t75069 = t75068 ^ t75068;
    wire t75070 = t75069 ^ t75069;
    wire t75071 = t75070 ^ t75070;
    wire t75072 = t75071 ^ t75071;
    wire t75073 = t75072 ^ t75072;
    wire t75074 = t75073 ^ t75073;
    wire t75075 = t75074 ^ t75074;
    wire t75076 = t75075 ^ t75075;
    wire t75077 = t75076 ^ t75076;
    wire t75078 = t75077 ^ t75077;
    wire t75079 = t75078 ^ t75078;
    wire t75080 = t75079 ^ t75079;
    wire t75081 = t75080 ^ t75080;
    wire t75082 = t75081 ^ t75081;
    wire t75083 = t75082 ^ t75082;
    wire t75084 = t75083 ^ t75083;
    wire t75085 = t75084 ^ t75084;
    wire t75086 = t75085 ^ t75085;
    wire t75087 = t75086 ^ t75086;
    wire t75088 = t75087 ^ t75087;
    wire t75089 = t75088 ^ t75088;
    wire t75090 = t75089 ^ t75089;
    wire t75091 = t75090 ^ t75090;
    wire t75092 = t75091 ^ t75091;
    wire t75093 = t75092 ^ t75092;
    wire t75094 = t75093 ^ t75093;
    wire t75095 = t75094 ^ t75094;
    wire t75096 = t75095 ^ t75095;
    wire t75097 = t75096 ^ t75096;
    wire t75098 = t75097 ^ t75097;
    wire t75099 = t75098 ^ t75098;
    wire t75100 = t75099 ^ t75099;
    wire t75101 = t75100 ^ t75100;
    wire t75102 = t75101 ^ t75101;
    wire t75103 = t75102 ^ t75102;
    wire t75104 = t75103 ^ t75103;
    wire t75105 = t75104 ^ t75104;
    wire t75106 = t75105 ^ t75105;
    wire t75107 = t75106 ^ t75106;
    wire t75108 = t75107 ^ t75107;
    wire t75109 = t75108 ^ t75108;
    wire t75110 = t75109 ^ t75109;
    wire t75111 = t75110 ^ t75110;
    wire t75112 = t75111 ^ t75111;
    wire t75113 = t75112 ^ t75112;
    wire t75114 = t75113 ^ t75113;
    wire t75115 = t75114 ^ t75114;
    wire t75116 = t75115 ^ t75115;
    wire t75117 = t75116 ^ t75116;
    wire t75118 = t75117 ^ t75117;
    wire t75119 = t75118 ^ t75118;
    wire t75120 = t75119 ^ t75119;
    wire t75121 = t75120 ^ t75120;
    wire t75122 = t75121 ^ t75121;
    wire t75123 = t75122 ^ t75122;
    wire t75124 = t75123 ^ t75123;
    wire t75125 = t75124 ^ t75124;
    wire t75126 = t75125 ^ t75125;
    wire t75127 = t75126 ^ t75126;
    wire t75128 = t75127 ^ t75127;
    wire t75129 = t75128 ^ t75128;
    wire t75130 = t75129 ^ t75129;
    wire t75131 = t75130 ^ t75130;
    wire t75132 = t75131 ^ t75131;
    wire t75133 = t75132 ^ t75132;
    wire t75134 = t75133 ^ t75133;
    wire t75135 = t75134 ^ t75134;
    wire t75136 = t75135 ^ t75135;
    wire t75137 = t75136 ^ t75136;
    wire t75138 = t75137 ^ t75137;
    wire t75139 = t75138 ^ t75138;
    wire t75140 = t75139 ^ t75139;
    wire t75141 = t75140 ^ t75140;
    wire t75142 = t75141 ^ t75141;
    wire t75143 = t75142 ^ t75142;
    wire t75144 = t75143 ^ t75143;
    wire t75145 = t75144 ^ t75144;
    wire t75146 = t75145 ^ t75145;
    wire t75147 = t75146 ^ t75146;
    wire t75148 = t75147 ^ t75147;
    wire t75149 = t75148 ^ t75148;
    wire t75150 = t75149 ^ t75149;
    wire t75151 = t75150 ^ t75150;
    wire t75152 = t75151 ^ t75151;
    wire t75153 = t75152 ^ t75152;
    wire t75154 = t75153 ^ t75153;
    wire t75155 = t75154 ^ t75154;
    wire t75156 = t75155 ^ t75155;
    wire t75157 = t75156 ^ t75156;
    wire t75158 = t75157 ^ t75157;
    wire t75159 = t75158 ^ t75158;
    wire t75160 = t75159 ^ t75159;
    wire t75161 = t75160 ^ t75160;
    wire t75162 = t75161 ^ t75161;
    wire t75163 = t75162 ^ t75162;
    wire t75164 = t75163 ^ t75163;
    wire t75165 = t75164 ^ t75164;
    wire t75166 = t75165 ^ t75165;
    wire t75167 = t75166 ^ t75166;
    wire t75168 = t75167 ^ t75167;
    wire t75169 = t75168 ^ t75168;
    wire t75170 = t75169 ^ t75169;
    wire t75171 = t75170 ^ t75170;
    wire t75172 = t75171 ^ t75171;
    wire t75173 = t75172 ^ t75172;
    wire t75174 = t75173 ^ t75173;
    wire t75175 = t75174 ^ t75174;
    wire t75176 = t75175 ^ t75175;
    wire t75177 = t75176 ^ t75176;
    wire t75178 = t75177 ^ t75177;
    wire t75179 = t75178 ^ t75178;
    wire t75180 = t75179 ^ t75179;
    wire t75181 = t75180 ^ t75180;
    wire t75182 = t75181 ^ t75181;
    wire t75183 = t75182 ^ t75182;
    wire t75184 = t75183 ^ t75183;
    wire t75185 = t75184 ^ t75184;
    wire t75186 = t75185 ^ t75185;
    wire t75187 = t75186 ^ t75186;
    wire t75188 = t75187 ^ t75187;
    wire t75189 = t75188 ^ t75188;
    wire t75190 = t75189 ^ t75189;
    wire t75191 = t75190 ^ t75190;
    wire t75192 = t75191 ^ t75191;
    wire t75193 = t75192 ^ t75192;
    wire t75194 = t75193 ^ t75193;
    wire t75195 = t75194 ^ t75194;
    wire t75196 = t75195 ^ t75195;
    wire t75197 = t75196 ^ t75196;
    wire t75198 = t75197 ^ t75197;
    wire t75199 = t75198 ^ t75198;
    wire t75200 = t75199 ^ t75199;
    wire t75201 = t75200 ^ t75200;
    wire t75202 = t75201 ^ t75201;
    wire t75203 = t75202 ^ t75202;
    wire t75204 = t75203 ^ t75203;
    wire t75205 = t75204 ^ t75204;
    wire t75206 = t75205 ^ t75205;
    wire t75207 = t75206 ^ t75206;
    wire t75208 = t75207 ^ t75207;
    wire t75209 = t75208 ^ t75208;
    wire t75210 = t75209 ^ t75209;
    wire t75211 = t75210 ^ t75210;
    wire t75212 = t75211 ^ t75211;
    wire t75213 = t75212 ^ t75212;
    wire t75214 = t75213 ^ t75213;
    wire t75215 = t75214 ^ t75214;
    wire t75216 = t75215 ^ t75215;
    wire t75217 = t75216 ^ t75216;
    wire t75218 = t75217 ^ t75217;
    wire t75219 = t75218 ^ t75218;
    wire t75220 = t75219 ^ t75219;
    wire t75221 = t75220 ^ t75220;
    wire t75222 = t75221 ^ t75221;
    wire t75223 = t75222 ^ t75222;
    wire t75224 = t75223 ^ t75223;
    wire t75225 = t75224 ^ t75224;
    wire t75226 = t75225 ^ t75225;
    wire t75227 = t75226 ^ t75226;
    wire t75228 = t75227 ^ t75227;
    wire t75229 = t75228 ^ t75228;
    wire t75230 = t75229 ^ t75229;
    wire t75231 = t75230 ^ t75230;
    wire t75232 = t75231 ^ t75231;
    wire t75233 = t75232 ^ t75232;
    wire t75234 = t75233 ^ t75233;
    wire t75235 = t75234 ^ t75234;
    wire t75236 = t75235 ^ t75235;
    wire t75237 = t75236 ^ t75236;
    wire t75238 = t75237 ^ t75237;
    wire t75239 = t75238 ^ t75238;
    wire t75240 = t75239 ^ t75239;
    wire t75241 = t75240 ^ t75240;
    wire t75242 = t75241 ^ t75241;
    wire t75243 = t75242 ^ t75242;
    wire t75244 = t75243 ^ t75243;
    wire t75245 = t75244 ^ t75244;
    wire t75246 = t75245 ^ t75245;
    wire t75247 = t75246 ^ t75246;
    wire t75248 = t75247 ^ t75247;
    wire t75249 = t75248 ^ t75248;
    wire t75250 = t75249 ^ t75249;
    wire t75251 = t75250 ^ t75250;
    wire t75252 = t75251 ^ t75251;
    wire t75253 = t75252 ^ t75252;
    wire t75254 = t75253 ^ t75253;
    wire t75255 = t75254 ^ t75254;
    wire t75256 = t75255 ^ t75255;
    wire t75257 = t75256 ^ t75256;
    wire t75258 = t75257 ^ t75257;
    wire t75259 = t75258 ^ t75258;
    wire t75260 = t75259 ^ t75259;
    wire t75261 = t75260 ^ t75260;
    wire t75262 = t75261 ^ t75261;
    wire t75263 = t75262 ^ t75262;
    wire t75264 = t75263 ^ t75263;
    wire t75265 = t75264 ^ t75264;
    wire t75266 = t75265 ^ t75265;
    wire t75267 = t75266 ^ t75266;
    wire t75268 = t75267 ^ t75267;
    wire t75269 = t75268 ^ t75268;
    wire t75270 = t75269 ^ t75269;
    wire t75271 = t75270 ^ t75270;
    wire t75272 = t75271 ^ t75271;
    wire t75273 = t75272 ^ t75272;
    wire t75274 = t75273 ^ t75273;
    wire t75275 = t75274 ^ t75274;
    wire t75276 = t75275 ^ t75275;
    wire t75277 = t75276 ^ t75276;
    wire t75278 = t75277 ^ t75277;
    wire t75279 = t75278 ^ t75278;
    wire t75280 = t75279 ^ t75279;
    wire t75281 = t75280 ^ t75280;
    wire t75282 = t75281 ^ t75281;
    wire t75283 = t75282 ^ t75282;
    wire t75284 = t75283 ^ t75283;
    wire t75285 = t75284 ^ t75284;
    wire t75286 = t75285 ^ t75285;
    wire t75287 = t75286 ^ t75286;
    wire t75288 = t75287 ^ t75287;
    wire t75289 = t75288 ^ t75288;
    wire t75290 = t75289 ^ t75289;
    wire t75291 = t75290 ^ t75290;
    wire t75292 = t75291 ^ t75291;
    wire t75293 = t75292 ^ t75292;
    wire t75294 = t75293 ^ t75293;
    wire t75295 = t75294 ^ t75294;
    wire t75296 = t75295 ^ t75295;
    wire t75297 = t75296 ^ t75296;
    wire t75298 = t75297 ^ t75297;
    wire t75299 = t75298 ^ t75298;
    wire t75300 = t75299 ^ t75299;
    wire t75301 = t75300 ^ t75300;
    wire t75302 = t75301 ^ t75301;
    wire t75303 = t75302 ^ t75302;
    wire t75304 = t75303 ^ t75303;
    wire t75305 = t75304 ^ t75304;
    wire t75306 = t75305 ^ t75305;
    wire t75307 = t75306 ^ t75306;
    wire t75308 = t75307 ^ t75307;
    wire t75309 = t75308 ^ t75308;
    wire t75310 = t75309 ^ t75309;
    wire t75311 = t75310 ^ t75310;
    wire t75312 = t75311 ^ t75311;
    wire t75313 = t75312 ^ t75312;
    wire t75314 = t75313 ^ t75313;
    wire t75315 = t75314 ^ t75314;
    wire t75316 = t75315 ^ t75315;
    wire t75317 = t75316 ^ t75316;
    wire t75318 = t75317 ^ t75317;
    wire t75319 = t75318 ^ t75318;
    wire t75320 = t75319 ^ t75319;
    wire t75321 = t75320 ^ t75320;
    wire t75322 = t75321 ^ t75321;
    wire t75323 = t75322 ^ t75322;
    wire t75324 = t75323 ^ t75323;
    wire t75325 = t75324 ^ t75324;
    wire t75326 = t75325 ^ t75325;
    wire t75327 = t75326 ^ t75326;
    wire t75328 = t75327 ^ t75327;
    wire t75329 = t75328 ^ t75328;
    wire t75330 = t75329 ^ t75329;
    wire t75331 = t75330 ^ t75330;
    wire t75332 = t75331 ^ t75331;
    wire t75333 = t75332 ^ t75332;
    wire t75334 = t75333 ^ t75333;
    wire t75335 = t75334 ^ t75334;
    wire t75336 = t75335 ^ t75335;
    wire t75337 = t75336 ^ t75336;
    wire t75338 = t75337 ^ t75337;
    wire t75339 = t75338 ^ t75338;
    wire t75340 = t75339 ^ t75339;
    wire t75341 = t75340 ^ t75340;
    wire t75342 = t75341 ^ t75341;
    wire t75343 = t75342 ^ t75342;
    wire t75344 = t75343 ^ t75343;
    wire t75345 = t75344 ^ t75344;
    wire t75346 = t75345 ^ t75345;
    wire t75347 = t75346 ^ t75346;
    wire t75348 = t75347 ^ t75347;
    wire t75349 = t75348 ^ t75348;
    wire t75350 = t75349 ^ t75349;
    wire t75351 = t75350 ^ t75350;
    wire t75352 = t75351 ^ t75351;
    wire t75353 = t75352 ^ t75352;
    wire t75354 = t75353 ^ t75353;
    wire t75355 = t75354 ^ t75354;
    wire t75356 = t75355 ^ t75355;
    wire t75357 = t75356 ^ t75356;
    wire t75358 = t75357 ^ t75357;
    wire t75359 = t75358 ^ t75358;
    wire t75360 = t75359 ^ t75359;
    wire t75361 = t75360 ^ t75360;
    wire t75362 = t75361 ^ t75361;
    wire t75363 = t75362 ^ t75362;
    wire t75364 = t75363 ^ t75363;
    wire t75365 = t75364 ^ t75364;
    wire t75366 = t75365 ^ t75365;
    wire t75367 = t75366 ^ t75366;
    wire t75368 = t75367 ^ t75367;
    wire t75369 = t75368 ^ t75368;
    wire t75370 = t75369 ^ t75369;
    wire t75371 = t75370 ^ t75370;
    wire t75372 = t75371 ^ t75371;
    wire t75373 = t75372 ^ t75372;
    wire t75374 = t75373 ^ t75373;
    wire t75375 = t75374 ^ t75374;
    wire t75376 = t75375 ^ t75375;
    wire t75377 = t75376 ^ t75376;
    wire t75378 = t75377 ^ t75377;
    wire t75379 = t75378 ^ t75378;
    wire t75380 = t75379 ^ t75379;
    wire t75381 = t75380 ^ t75380;
    wire t75382 = t75381 ^ t75381;
    wire t75383 = t75382 ^ t75382;
    wire t75384 = t75383 ^ t75383;
    wire t75385 = t75384 ^ t75384;
    wire t75386 = t75385 ^ t75385;
    wire t75387 = t75386 ^ t75386;
    wire t75388 = t75387 ^ t75387;
    wire t75389 = t75388 ^ t75388;
    wire t75390 = t75389 ^ t75389;
    wire t75391 = t75390 ^ t75390;
    wire t75392 = t75391 ^ t75391;
    wire t75393 = t75392 ^ t75392;
    wire t75394 = t75393 ^ t75393;
    wire t75395 = t75394 ^ t75394;
    wire t75396 = t75395 ^ t75395;
    wire t75397 = t75396 ^ t75396;
    wire t75398 = t75397 ^ t75397;
    wire t75399 = t75398 ^ t75398;
    wire t75400 = t75399 ^ t75399;
    wire t75401 = t75400 ^ t75400;
    wire t75402 = t75401 ^ t75401;
    wire t75403 = t75402 ^ t75402;
    wire t75404 = t75403 ^ t75403;
    wire t75405 = t75404 ^ t75404;
    wire t75406 = t75405 ^ t75405;
    wire t75407 = t75406 ^ t75406;
    wire t75408 = t75407 ^ t75407;
    wire t75409 = t75408 ^ t75408;
    wire t75410 = t75409 ^ t75409;
    wire t75411 = t75410 ^ t75410;
    wire t75412 = t75411 ^ t75411;
    wire t75413 = t75412 ^ t75412;
    wire t75414 = t75413 ^ t75413;
    wire t75415 = t75414 ^ t75414;
    wire t75416 = t75415 ^ t75415;
    wire t75417 = t75416 ^ t75416;
    wire t75418 = t75417 ^ t75417;
    wire t75419 = t75418 ^ t75418;
    wire t75420 = t75419 ^ t75419;
    wire t75421 = t75420 ^ t75420;
    wire t75422 = t75421 ^ t75421;
    wire t75423 = t75422 ^ t75422;
    wire t75424 = t75423 ^ t75423;
    wire t75425 = t75424 ^ t75424;
    wire t75426 = t75425 ^ t75425;
    wire t75427 = t75426 ^ t75426;
    wire t75428 = t75427 ^ t75427;
    wire t75429 = t75428 ^ t75428;
    wire t75430 = t75429 ^ t75429;
    wire t75431 = t75430 ^ t75430;
    wire t75432 = t75431 ^ t75431;
    wire t75433 = t75432 ^ t75432;
    wire t75434 = t75433 ^ t75433;
    wire t75435 = t75434 ^ t75434;
    wire t75436 = t75435 ^ t75435;
    wire t75437 = t75436 ^ t75436;
    wire t75438 = t75437 ^ t75437;
    wire t75439 = t75438 ^ t75438;
    wire t75440 = t75439 ^ t75439;
    wire t75441 = t75440 ^ t75440;
    wire t75442 = t75441 ^ t75441;
    wire t75443 = t75442 ^ t75442;
    wire t75444 = t75443 ^ t75443;
    wire t75445 = t75444 ^ t75444;
    wire t75446 = t75445 ^ t75445;
    wire t75447 = t75446 ^ t75446;
    wire t75448 = t75447 ^ t75447;
    wire t75449 = t75448 ^ t75448;
    wire t75450 = t75449 ^ t75449;
    wire t75451 = t75450 ^ t75450;
    wire t75452 = t75451 ^ t75451;
    wire t75453 = t75452 ^ t75452;
    wire t75454 = t75453 ^ t75453;
    wire t75455 = t75454 ^ t75454;
    wire t75456 = t75455 ^ t75455;
    wire t75457 = t75456 ^ t75456;
    wire t75458 = t75457 ^ t75457;
    wire t75459 = t75458 ^ t75458;
    wire t75460 = t75459 ^ t75459;
    wire t75461 = t75460 ^ t75460;
    wire t75462 = t75461 ^ t75461;
    wire t75463 = t75462 ^ t75462;
    wire t75464 = t75463 ^ t75463;
    wire t75465 = t75464 ^ t75464;
    wire t75466 = t75465 ^ t75465;
    wire t75467 = t75466 ^ t75466;
    wire t75468 = t75467 ^ t75467;
    wire t75469 = t75468 ^ t75468;
    wire t75470 = t75469 ^ t75469;
    wire t75471 = t75470 ^ t75470;
    wire t75472 = t75471 ^ t75471;
    wire t75473 = t75472 ^ t75472;
    wire t75474 = t75473 ^ t75473;
    wire t75475 = t75474 ^ t75474;
    wire t75476 = t75475 ^ t75475;
    wire t75477 = t75476 ^ t75476;
    wire t75478 = t75477 ^ t75477;
    wire t75479 = t75478 ^ t75478;
    wire t75480 = t75479 ^ t75479;
    wire t75481 = t75480 ^ t75480;
    wire t75482 = t75481 ^ t75481;
    wire t75483 = t75482 ^ t75482;
    wire t75484 = t75483 ^ t75483;
    wire t75485 = t75484 ^ t75484;
    wire t75486 = t75485 ^ t75485;
    wire t75487 = t75486 ^ t75486;
    wire t75488 = t75487 ^ t75487;
    wire t75489 = t75488 ^ t75488;
    wire t75490 = t75489 ^ t75489;
    wire t75491 = t75490 ^ t75490;
    wire t75492 = t75491 ^ t75491;
    wire t75493 = t75492 ^ t75492;
    wire t75494 = t75493 ^ t75493;
    wire t75495 = t75494 ^ t75494;
    wire t75496 = t75495 ^ t75495;
    wire t75497 = t75496 ^ t75496;
    wire t75498 = t75497 ^ t75497;
    wire t75499 = t75498 ^ t75498;
    wire t75500 = t75499 ^ t75499;
    wire t75501 = t75500 ^ t75500;
    wire t75502 = t75501 ^ t75501;
    wire t75503 = t75502 ^ t75502;
    wire t75504 = t75503 ^ t75503;
    wire t75505 = t75504 ^ t75504;
    wire t75506 = t75505 ^ t75505;
    wire t75507 = t75506 ^ t75506;
    wire t75508 = t75507 ^ t75507;
    wire t75509 = t75508 ^ t75508;
    wire t75510 = t75509 ^ t75509;
    wire t75511 = t75510 ^ t75510;
    wire t75512 = t75511 ^ t75511;
    wire t75513 = t75512 ^ t75512;
    wire t75514 = t75513 ^ t75513;
    wire t75515 = t75514 ^ t75514;
    wire t75516 = t75515 ^ t75515;
    wire t75517 = t75516 ^ t75516;
    wire t75518 = t75517 ^ t75517;
    wire t75519 = t75518 ^ t75518;
    wire t75520 = t75519 ^ t75519;
    wire t75521 = t75520 ^ t75520;
    wire t75522 = t75521 ^ t75521;
    wire t75523 = t75522 ^ t75522;
    wire t75524 = t75523 ^ t75523;
    wire t75525 = t75524 ^ t75524;
    wire t75526 = t75525 ^ t75525;
    wire t75527 = t75526 ^ t75526;
    wire t75528 = t75527 ^ t75527;
    wire t75529 = t75528 ^ t75528;
    wire t75530 = t75529 ^ t75529;
    wire t75531 = t75530 ^ t75530;
    wire t75532 = t75531 ^ t75531;
    wire t75533 = t75532 ^ t75532;
    wire t75534 = t75533 ^ t75533;
    wire t75535 = t75534 ^ t75534;
    wire t75536 = t75535 ^ t75535;
    wire t75537 = t75536 ^ t75536;
    wire t75538 = t75537 ^ t75537;
    wire t75539 = t75538 ^ t75538;
    wire t75540 = t75539 ^ t75539;
    wire t75541 = t75540 ^ t75540;
    wire t75542 = t75541 ^ t75541;
    wire t75543 = t75542 ^ t75542;
    wire t75544 = t75543 ^ t75543;
    wire t75545 = t75544 ^ t75544;
    wire t75546 = t75545 ^ t75545;
    wire t75547 = t75546 ^ t75546;
    wire t75548 = t75547 ^ t75547;
    wire t75549 = t75548 ^ t75548;
    wire t75550 = t75549 ^ t75549;
    wire t75551 = t75550 ^ t75550;
    wire t75552 = t75551 ^ t75551;
    wire t75553 = t75552 ^ t75552;
    wire t75554 = t75553 ^ t75553;
    wire t75555 = t75554 ^ t75554;
    wire t75556 = t75555 ^ t75555;
    wire t75557 = t75556 ^ t75556;
    wire t75558 = t75557 ^ t75557;
    wire t75559 = t75558 ^ t75558;
    wire t75560 = t75559 ^ t75559;
    wire t75561 = t75560 ^ t75560;
    wire t75562 = t75561 ^ t75561;
    wire t75563 = t75562 ^ t75562;
    wire t75564 = t75563 ^ t75563;
    wire t75565 = t75564 ^ t75564;
    wire t75566 = t75565 ^ t75565;
    wire t75567 = t75566 ^ t75566;
    wire t75568 = t75567 ^ t75567;
    wire t75569 = t75568 ^ t75568;
    wire t75570 = t75569 ^ t75569;
    wire t75571 = t75570 ^ t75570;
    wire t75572 = t75571 ^ t75571;
    wire t75573 = t75572 ^ t75572;
    wire t75574 = t75573 ^ t75573;
    wire t75575 = t75574 ^ t75574;
    wire t75576 = t75575 ^ t75575;
    wire t75577 = t75576 ^ t75576;
    wire t75578 = t75577 ^ t75577;
    wire t75579 = t75578 ^ t75578;
    wire t75580 = t75579 ^ t75579;
    wire t75581 = t75580 ^ t75580;
    wire t75582 = t75581 ^ t75581;
    wire t75583 = t75582 ^ t75582;
    wire t75584 = t75583 ^ t75583;
    wire t75585 = t75584 ^ t75584;
    wire t75586 = t75585 ^ t75585;
    wire t75587 = t75586 ^ t75586;
    wire t75588 = t75587 ^ t75587;
    wire t75589 = t75588 ^ t75588;
    wire t75590 = t75589 ^ t75589;
    wire t75591 = t75590 ^ t75590;
    wire t75592 = t75591 ^ t75591;
    wire t75593 = t75592 ^ t75592;
    wire t75594 = t75593 ^ t75593;
    wire t75595 = t75594 ^ t75594;
    wire t75596 = t75595 ^ t75595;
    wire t75597 = t75596 ^ t75596;
    wire t75598 = t75597 ^ t75597;
    wire t75599 = t75598 ^ t75598;
    wire t75600 = t75599 ^ t75599;
    wire t75601 = t75600 ^ t75600;
    wire t75602 = t75601 ^ t75601;
    wire t75603 = t75602 ^ t75602;
    wire t75604 = t75603 ^ t75603;
    wire t75605 = t75604 ^ t75604;
    wire t75606 = t75605 ^ t75605;
    wire t75607 = t75606 ^ t75606;
    wire t75608 = t75607 ^ t75607;
    wire t75609 = t75608 ^ t75608;
    wire t75610 = t75609 ^ t75609;
    wire t75611 = t75610 ^ t75610;
    wire t75612 = t75611 ^ t75611;
    wire t75613 = t75612 ^ t75612;
    wire t75614 = t75613 ^ t75613;
    wire t75615 = t75614 ^ t75614;
    wire t75616 = t75615 ^ t75615;
    wire t75617 = t75616 ^ t75616;
    wire t75618 = t75617 ^ t75617;
    wire t75619 = t75618 ^ t75618;
    wire t75620 = t75619 ^ t75619;
    wire t75621 = t75620 ^ t75620;
    wire t75622 = t75621 ^ t75621;
    wire t75623 = t75622 ^ t75622;
    wire t75624 = t75623 ^ t75623;
    wire t75625 = t75624 ^ t75624;
    wire t75626 = t75625 ^ t75625;
    wire t75627 = t75626 ^ t75626;
    wire t75628 = t75627 ^ t75627;
    wire t75629 = t75628 ^ t75628;
    wire t75630 = t75629 ^ t75629;
    wire t75631 = t75630 ^ t75630;
    wire t75632 = t75631 ^ t75631;
    wire t75633 = t75632 ^ t75632;
    wire t75634 = t75633 ^ t75633;
    wire t75635 = t75634 ^ t75634;
    wire t75636 = t75635 ^ t75635;
    wire t75637 = t75636 ^ t75636;
    wire t75638 = t75637 ^ t75637;
    wire t75639 = t75638 ^ t75638;
    wire t75640 = t75639 ^ t75639;
    wire t75641 = t75640 ^ t75640;
    wire t75642 = t75641 ^ t75641;
    wire t75643 = t75642 ^ t75642;
    wire t75644 = t75643 ^ t75643;
    wire t75645 = t75644 ^ t75644;
    wire t75646 = t75645 ^ t75645;
    wire t75647 = t75646 ^ t75646;
    wire t75648 = t75647 ^ t75647;
    wire t75649 = t75648 ^ t75648;
    wire t75650 = t75649 ^ t75649;
    wire t75651 = t75650 ^ t75650;
    wire t75652 = t75651 ^ t75651;
    wire t75653 = t75652 ^ t75652;
    wire t75654 = t75653 ^ t75653;
    wire t75655 = t75654 ^ t75654;
    wire t75656 = t75655 ^ t75655;
    wire t75657 = t75656 ^ t75656;
    wire t75658 = t75657 ^ t75657;
    wire t75659 = t75658 ^ t75658;
    wire t75660 = t75659 ^ t75659;
    wire t75661 = t75660 ^ t75660;
    wire t75662 = t75661 ^ t75661;
    wire t75663 = t75662 ^ t75662;
    wire t75664 = t75663 ^ t75663;
    wire t75665 = t75664 ^ t75664;
    wire t75666 = t75665 ^ t75665;
    wire t75667 = t75666 ^ t75666;
    wire t75668 = t75667 ^ t75667;
    wire t75669 = t75668 ^ t75668;
    wire t75670 = t75669 ^ t75669;
    wire t75671 = t75670 ^ t75670;
    wire t75672 = t75671 ^ t75671;
    wire t75673 = t75672 ^ t75672;
    wire t75674 = t75673 ^ t75673;
    wire t75675 = t75674 ^ t75674;
    wire t75676 = t75675 ^ t75675;
    wire t75677 = t75676 ^ t75676;
    wire t75678 = t75677 ^ t75677;
    wire t75679 = t75678 ^ t75678;
    wire t75680 = t75679 ^ t75679;
    wire t75681 = t75680 ^ t75680;
    wire t75682 = t75681 ^ t75681;
    wire t75683 = t75682 ^ t75682;
    wire t75684 = t75683 ^ t75683;
    wire t75685 = t75684 ^ t75684;
    wire t75686 = t75685 ^ t75685;
    wire t75687 = t75686 ^ t75686;
    wire t75688 = t75687 ^ t75687;
    wire t75689 = t75688 ^ t75688;
    wire t75690 = t75689 ^ t75689;
    wire t75691 = t75690 ^ t75690;
    wire t75692 = t75691 ^ t75691;
    wire t75693 = t75692 ^ t75692;
    wire t75694 = t75693 ^ t75693;
    wire t75695 = t75694 ^ t75694;
    wire t75696 = t75695 ^ t75695;
    wire t75697 = t75696 ^ t75696;
    wire t75698 = t75697 ^ t75697;
    wire t75699 = t75698 ^ t75698;
    wire t75700 = t75699 ^ t75699;
    wire t75701 = t75700 ^ t75700;
    wire t75702 = t75701 ^ t75701;
    wire t75703 = t75702 ^ t75702;
    wire t75704 = t75703 ^ t75703;
    wire t75705 = t75704 ^ t75704;
    wire t75706 = t75705 ^ t75705;
    wire t75707 = t75706 ^ t75706;
    wire t75708 = t75707 ^ t75707;
    wire t75709 = t75708 ^ t75708;
    wire t75710 = t75709 ^ t75709;
    wire t75711 = t75710 ^ t75710;
    wire t75712 = t75711 ^ t75711;
    wire t75713 = t75712 ^ t75712;
    wire t75714 = t75713 ^ t75713;
    wire t75715 = t75714 ^ t75714;
    wire t75716 = t75715 ^ t75715;
    wire t75717 = t75716 ^ t75716;
    wire t75718 = t75717 ^ t75717;
    wire t75719 = t75718 ^ t75718;
    wire t75720 = t75719 ^ t75719;
    wire t75721 = t75720 ^ t75720;
    wire t75722 = t75721 ^ t75721;
    wire t75723 = t75722 ^ t75722;
    wire t75724 = t75723 ^ t75723;
    wire t75725 = t75724 ^ t75724;
    wire t75726 = t75725 ^ t75725;
    wire t75727 = t75726 ^ t75726;
    wire t75728 = t75727 ^ t75727;
    wire t75729 = t75728 ^ t75728;
    wire t75730 = t75729 ^ t75729;
    wire t75731 = t75730 ^ t75730;
    wire t75732 = t75731 ^ t75731;
    wire t75733 = t75732 ^ t75732;
    wire t75734 = t75733 ^ t75733;
    wire t75735 = t75734 ^ t75734;
    wire t75736 = t75735 ^ t75735;
    wire t75737 = t75736 ^ t75736;
    wire t75738 = t75737 ^ t75737;
    wire t75739 = t75738 ^ t75738;
    wire t75740 = t75739 ^ t75739;
    wire t75741 = t75740 ^ t75740;
    wire t75742 = t75741 ^ t75741;
    wire t75743 = t75742 ^ t75742;
    wire t75744 = t75743 ^ t75743;
    wire t75745 = t75744 ^ t75744;
    wire t75746 = t75745 ^ t75745;
    wire t75747 = t75746 ^ t75746;
    wire t75748 = t75747 ^ t75747;
    wire t75749 = t75748 ^ t75748;
    wire t75750 = t75749 ^ t75749;
    wire t75751 = t75750 ^ t75750;
    wire t75752 = t75751 ^ t75751;
    wire t75753 = t75752 ^ t75752;
    wire t75754 = t75753 ^ t75753;
    wire t75755 = t75754 ^ t75754;
    wire t75756 = t75755 ^ t75755;
    wire t75757 = t75756 ^ t75756;
    wire t75758 = t75757 ^ t75757;
    wire t75759 = t75758 ^ t75758;
    wire t75760 = t75759 ^ t75759;
    wire t75761 = t75760 ^ t75760;
    wire t75762 = t75761 ^ t75761;
    wire t75763 = t75762 ^ t75762;
    wire t75764 = t75763 ^ t75763;
    wire t75765 = t75764 ^ t75764;
    wire t75766 = t75765 ^ t75765;
    wire t75767 = t75766 ^ t75766;
    wire t75768 = t75767 ^ t75767;
    wire t75769 = t75768 ^ t75768;
    wire t75770 = t75769 ^ t75769;
    wire t75771 = t75770 ^ t75770;
    wire t75772 = t75771 ^ t75771;
    wire t75773 = t75772 ^ t75772;
    wire t75774 = t75773 ^ t75773;
    wire t75775 = t75774 ^ t75774;
    wire t75776 = t75775 ^ t75775;
    wire t75777 = t75776 ^ t75776;
    wire t75778 = t75777 ^ t75777;
    wire t75779 = t75778 ^ t75778;
    wire t75780 = t75779 ^ t75779;
    wire t75781 = t75780 ^ t75780;
    wire t75782 = t75781 ^ t75781;
    wire t75783 = t75782 ^ t75782;
    wire t75784 = t75783 ^ t75783;
    wire t75785 = t75784 ^ t75784;
    wire t75786 = t75785 ^ t75785;
    wire t75787 = t75786 ^ t75786;
    wire t75788 = t75787 ^ t75787;
    wire t75789 = t75788 ^ t75788;
    wire t75790 = t75789 ^ t75789;
    wire t75791 = t75790 ^ t75790;
    wire t75792 = t75791 ^ t75791;
    wire t75793 = t75792 ^ t75792;
    wire t75794 = t75793 ^ t75793;
    wire t75795 = t75794 ^ t75794;
    wire t75796 = t75795 ^ t75795;
    wire t75797 = t75796 ^ t75796;
    wire t75798 = t75797 ^ t75797;
    wire t75799 = t75798 ^ t75798;
    wire t75800 = t75799 ^ t75799;
    wire t75801 = t75800 ^ t75800;
    wire t75802 = t75801 ^ t75801;
    wire t75803 = t75802 ^ t75802;
    wire t75804 = t75803 ^ t75803;
    wire t75805 = t75804 ^ t75804;
    wire t75806 = t75805 ^ t75805;
    wire t75807 = t75806 ^ t75806;
    wire t75808 = t75807 ^ t75807;
    wire t75809 = t75808 ^ t75808;
    wire t75810 = t75809 ^ t75809;
    wire t75811 = t75810 ^ t75810;
    wire t75812 = t75811 ^ t75811;
    wire t75813 = t75812 ^ t75812;
    wire t75814 = t75813 ^ t75813;
    wire t75815 = t75814 ^ t75814;
    wire t75816 = t75815 ^ t75815;
    wire t75817 = t75816 ^ t75816;
    wire t75818 = t75817 ^ t75817;
    wire t75819 = t75818 ^ t75818;
    wire t75820 = t75819 ^ t75819;
    wire t75821 = t75820 ^ t75820;
    wire t75822 = t75821 ^ t75821;
    wire t75823 = t75822 ^ t75822;
    wire t75824 = t75823 ^ t75823;
    wire t75825 = t75824 ^ t75824;
    wire t75826 = t75825 ^ t75825;
    wire t75827 = t75826 ^ t75826;
    wire t75828 = t75827 ^ t75827;
    wire t75829 = t75828 ^ t75828;
    wire t75830 = t75829 ^ t75829;
    wire t75831 = t75830 ^ t75830;
    wire t75832 = t75831 ^ t75831;
    wire t75833 = t75832 ^ t75832;
    wire t75834 = t75833 ^ t75833;
    wire t75835 = t75834 ^ t75834;
    wire t75836 = t75835 ^ t75835;
    wire t75837 = t75836 ^ t75836;
    wire t75838 = t75837 ^ t75837;
    wire t75839 = t75838 ^ t75838;
    wire t75840 = t75839 ^ t75839;
    wire t75841 = t75840 ^ t75840;
    wire t75842 = t75841 ^ t75841;
    wire t75843 = t75842 ^ t75842;
    wire t75844 = t75843 ^ t75843;
    wire t75845 = t75844 ^ t75844;
    wire t75846 = t75845 ^ t75845;
    wire t75847 = t75846 ^ t75846;
    wire t75848 = t75847 ^ t75847;
    wire t75849 = t75848 ^ t75848;
    wire t75850 = t75849 ^ t75849;
    wire t75851 = t75850 ^ t75850;
    wire t75852 = t75851 ^ t75851;
    wire t75853 = t75852 ^ t75852;
    wire t75854 = t75853 ^ t75853;
    wire t75855 = t75854 ^ t75854;
    wire t75856 = t75855 ^ t75855;
    wire t75857 = t75856 ^ t75856;
    wire t75858 = t75857 ^ t75857;
    wire t75859 = t75858 ^ t75858;
    wire t75860 = t75859 ^ t75859;
    wire t75861 = t75860 ^ t75860;
    wire t75862 = t75861 ^ t75861;
    wire t75863 = t75862 ^ t75862;
    wire t75864 = t75863 ^ t75863;
    wire t75865 = t75864 ^ t75864;
    wire t75866 = t75865 ^ t75865;
    wire t75867 = t75866 ^ t75866;
    wire t75868 = t75867 ^ t75867;
    wire t75869 = t75868 ^ t75868;
    wire t75870 = t75869 ^ t75869;
    wire t75871 = t75870 ^ t75870;
    wire t75872 = t75871 ^ t75871;
    wire t75873 = t75872 ^ t75872;
    wire t75874 = t75873 ^ t75873;
    wire t75875 = t75874 ^ t75874;
    wire t75876 = t75875 ^ t75875;
    wire t75877 = t75876 ^ t75876;
    wire t75878 = t75877 ^ t75877;
    wire t75879 = t75878 ^ t75878;
    wire t75880 = t75879 ^ t75879;
    wire t75881 = t75880 ^ t75880;
    wire t75882 = t75881 ^ t75881;
    wire t75883 = t75882 ^ t75882;
    wire t75884 = t75883 ^ t75883;
    wire t75885 = t75884 ^ t75884;
    wire t75886 = t75885 ^ t75885;
    wire t75887 = t75886 ^ t75886;
    wire t75888 = t75887 ^ t75887;
    wire t75889 = t75888 ^ t75888;
    wire t75890 = t75889 ^ t75889;
    wire t75891 = t75890 ^ t75890;
    wire t75892 = t75891 ^ t75891;
    wire t75893 = t75892 ^ t75892;
    wire t75894 = t75893 ^ t75893;
    wire t75895 = t75894 ^ t75894;
    wire t75896 = t75895 ^ t75895;
    wire t75897 = t75896 ^ t75896;
    wire t75898 = t75897 ^ t75897;
    wire t75899 = t75898 ^ t75898;
    wire t75900 = t75899 ^ t75899;
    wire t75901 = t75900 ^ t75900;
    wire t75902 = t75901 ^ t75901;
    wire t75903 = t75902 ^ t75902;
    wire t75904 = t75903 ^ t75903;
    wire t75905 = t75904 ^ t75904;
    wire t75906 = t75905 ^ t75905;
    wire t75907 = t75906 ^ t75906;
    wire t75908 = t75907 ^ t75907;
    wire t75909 = t75908 ^ t75908;
    wire t75910 = t75909 ^ t75909;
    wire t75911 = t75910 ^ t75910;
    wire t75912 = t75911 ^ t75911;
    wire t75913 = t75912 ^ t75912;
    wire t75914 = t75913 ^ t75913;
    wire t75915 = t75914 ^ t75914;
    wire t75916 = t75915 ^ t75915;
    wire t75917 = t75916 ^ t75916;
    wire t75918 = t75917 ^ t75917;
    wire t75919 = t75918 ^ t75918;
    wire t75920 = t75919 ^ t75919;
    wire t75921 = t75920 ^ t75920;
    wire t75922 = t75921 ^ t75921;
    wire t75923 = t75922 ^ t75922;
    wire t75924 = t75923 ^ t75923;
    wire t75925 = t75924 ^ t75924;
    wire t75926 = t75925 ^ t75925;
    wire t75927 = t75926 ^ t75926;
    wire t75928 = t75927 ^ t75927;
    wire t75929 = t75928 ^ t75928;
    wire t75930 = t75929 ^ t75929;
    wire t75931 = t75930 ^ t75930;
    wire t75932 = t75931 ^ t75931;
    wire t75933 = t75932 ^ t75932;
    wire t75934 = t75933 ^ t75933;
    wire t75935 = t75934 ^ t75934;
    wire t75936 = t75935 ^ t75935;
    wire t75937 = t75936 ^ t75936;
    wire t75938 = t75937 ^ t75937;
    wire t75939 = t75938 ^ t75938;
    wire t75940 = t75939 ^ t75939;
    wire t75941 = t75940 ^ t75940;
    wire t75942 = t75941 ^ t75941;
    wire t75943 = t75942 ^ t75942;
    wire t75944 = t75943 ^ t75943;
    wire t75945 = t75944 ^ t75944;
    wire t75946 = t75945 ^ t75945;
    wire t75947 = t75946 ^ t75946;
    wire t75948 = t75947 ^ t75947;
    wire t75949 = t75948 ^ t75948;
    wire t75950 = t75949 ^ t75949;
    wire t75951 = t75950 ^ t75950;
    wire t75952 = t75951 ^ t75951;
    wire t75953 = t75952 ^ t75952;
    wire t75954 = t75953 ^ t75953;
    wire t75955 = t75954 ^ t75954;
    wire t75956 = t75955 ^ t75955;
    wire t75957 = t75956 ^ t75956;
    wire t75958 = t75957 ^ t75957;
    wire t75959 = t75958 ^ t75958;
    wire t75960 = t75959 ^ t75959;
    wire t75961 = t75960 ^ t75960;
    wire t75962 = t75961 ^ t75961;
    wire t75963 = t75962 ^ t75962;
    wire t75964 = t75963 ^ t75963;
    wire t75965 = t75964 ^ t75964;
    wire t75966 = t75965 ^ t75965;
    wire t75967 = t75966 ^ t75966;
    wire t75968 = t75967 ^ t75967;
    wire t75969 = t75968 ^ t75968;
    wire t75970 = t75969 ^ t75969;
    wire t75971 = t75970 ^ t75970;
    wire t75972 = t75971 ^ t75971;
    wire t75973 = t75972 ^ t75972;
    wire t75974 = t75973 ^ t75973;
    wire t75975 = t75974 ^ t75974;
    wire t75976 = t75975 ^ t75975;
    wire t75977 = t75976 ^ t75976;
    wire t75978 = t75977 ^ t75977;
    wire t75979 = t75978 ^ t75978;
    wire t75980 = t75979 ^ t75979;
    wire t75981 = t75980 ^ t75980;
    wire t75982 = t75981 ^ t75981;
    wire t75983 = t75982 ^ t75982;
    wire t75984 = t75983 ^ t75983;
    wire t75985 = t75984 ^ t75984;
    wire t75986 = t75985 ^ t75985;
    wire t75987 = t75986 ^ t75986;
    wire t75988 = t75987 ^ t75987;
    wire t75989 = t75988 ^ t75988;
    wire t75990 = t75989 ^ t75989;
    wire t75991 = t75990 ^ t75990;
    wire t75992 = t75991 ^ t75991;
    wire t75993 = t75992 ^ t75992;
    wire t75994 = t75993 ^ t75993;
    wire t75995 = t75994 ^ t75994;
    wire t75996 = t75995 ^ t75995;
    wire t75997 = t75996 ^ t75996;
    wire t75998 = t75997 ^ t75997;
    wire t75999 = t75998 ^ t75998;
    wire t76000 = t75999 ^ t75999;
    wire t76001 = t76000 ^ t76000;
    wire t76002 = t76001 ^ t76001;
    wire t76003 = t76002 ^ t76002;
    wire t76004 = t76003 ^ t76003;
    wire t76005 = t76004 ^ t76004;
    wire t76006 = t76005 ^ t76005;
    wire t76007 = t76006 ^ t76006;
    wire t76008 = t76007 ^ t76007;
    wire t76009 = t76008 ^ t76008;
    wire t76010 = t76009 ^ t76009;
    wire t76011 = t76010 ^ t76010;
    wire t76012 = t76011 ^ t76011;
    wire t76013 = t76012 ^ t76012;
    wire t76014 = t76013 ^ t76013;
    wire t76015 = t76014 ^ t76014;
    wire t76016 = t76015 ^ t76015;
    wire t76017 = t76016 ^ t76016;
    wire t76018 = t76017 ^ t76017;
    wire t76019 = t76018 ^ t76018;
    wire t76020 = t76019 ^ t76019;
    wire t76021 = t76020 ^ t76020;
    wire t76022 = t76021 ^ t76021;
    wire t76023 = t76022 ^ t76022;
    wire t76024 = t76023 ^ t76023;
    wire t76025 = t76024 ^ t76024;
    wire t76026 = t76025 ^ t76025;
    wire t76027 = t76026 ^ t76026;
    wire t76028 = t76027 ^ t76027;
    wire t76029 = t76028 ^ t76028;
    wire t76030 = t76029 ^ t76029;
    wire t76031 = t76030 ^ t76030;
    wire t76032 = t76031 ^ t76031;
    wire t76033 = t76032 ^ t76032;
    wire t76034 = t76033 ^ t76033;
    wire t76035 = t76034 ^ t76034;
    wire t76036 = t76035 ^ t76035;
    wire t76037 = t76036 ^ t76036;
    wire t76038 = t76037 ^ t76037;
    wire t76039 = t76038 ^ t76038;
    wire t76040 = t76039 ^ t76039;
    wire t76041 = t76040 ^ t76040;
    wire t76042 = t76041 ^ t76041;
    wire t76043 = t76042 ^ t76042;
    wire t76044 = t76043 ^ t76043;
    wire t76045 = t76044 ^ t76044;
    wire t76046 = t76045 ^ t76045;
    wire t76047 = t76046 ^ t76046;
    wire t76048 = t76047 ^ t76047;
    wire t76049 = t76048 ^ t76048;
    wire t76050 = t76049 ^ t76049;
    wire t76051 = t76050 ^ t76050;
    wire t76052 = t76051 ^ t76051;
    wire t76053 = t76052 ^ t76052;
    wire t76054 = t76053 ^ t76053;
    wire t76055 = t76054 ^ t76054;
    wire t76056 = t76055 ^ t76055;
    wire t76057 = t76056 ^ t76056;
    wire t76058 = t76057 ^ t76057;
    wire t76059 = t76058 ^ t76058;
    wire t76060 = t76059 ^ t76059;
    wire t76061 = t76060 ^ t76060;
    wire t76062 = t76061 ^ t76061;
    wire t76063 = t76062 ^ t76062;
    wire t76064 = t76063 ^ t76063;
    wire t76065 = t76064 ^ t76064;
    wire t76066 = t76065 ^ t76065;
    wire t76067 = t76066 ^ t76066;
    wire t76068 = t76067 ^ t76067;
    wire t76069 = t76068 ^ t76068;
    wire t76070 = t76069 ^ t76069;
    wire t76071 = t76070 ^ t76070;
    wire t76072 = t76071 ^ t76071;
    wire t76073 = t76072 ^ t76072;
    wire t76074 = t76073 ^ t76073;
    wire t76075 = t76074 ^ t76074;
    wire t76076 = t76075 ^ t76075;
    wire t76077 = t76076 ^ t76076;
    wire t76078 = t76077 ^ t76077;
    wire t76079 = t76078 ^ t76078;
    wire t76080 = t76079 ^ t76079;
    wire t76081 = t76080 ^ t76080;
    wire t76082 = t76081 ^ t76081;
    wire t76083 = t76082 ^ t76082;
    wire t76084 = t76083 ^ t76083;
    wire t76085 = t76084 ^ t76084;
    wire t76086 = t76085 ^ t76085;
    wire t76087 = t76086 ^ t76086;
    wire t76088 = t76087 ^ t76087;
    wire t76089 = t76088 ^ t76088;
    wire t76090 = t76089 ^ t76089;
    wire t76091 = t76090 ^ t76090;
    wire t76092 = t76091 ^ t76091;
    wire t76093 = t76092 ^ t76092;
    wire t76094 = t76093 ^ t76093;
    wire t76095 = t76094 ^ t76094;
    wire t76096 = t76095 ^ t76095;
    wire t76097 = t76096 ^ t76096;
    wire t76098 = t76097 ^ t76097;
    wire t76099 = t76098 ^ t76098;
    wire t76100 = t76099 ^ t76099;
    wire t76101 = t76100 ^ t76100;
    wire t76102 = t76101 ^ t76101;
    wire t76103 = t76102 ^ t76102;
    wire t76104 = t76103 ^ t76103;
    wire t76105 = t76104 ^ t76104;
    wire t76106 = t76105 ^ t76105;
    wire t76107 = t76106 ^ t76106;
    wire t76108 = t76107 ^ t76107;
    wire t76109 = t76108 ^ t76108;
    wire t76110 = t76109 ^ t76109;
    wire t76111 = t76110 ^ t76110;
    wire t76112 = t76111 ^ t76111;
    wire t76113 = t76112 ^ t76112;
    wire t76114 = t76113 ^ t76113;
    wire t76115 = t76114 ^ t76114;
    wire t76116 = t76115 ^ t76115;
    wire t76117 = t76116 ^ t76116;
    wire t76118 = t76117 ^ t76117;
    wire t76119 = t76118 ^ t76118;
    wire t76120 = t76119 ^ t76119;
    wire t76121 = t76120 ^ t76120;
    wire t76122 = t76121 ^ t76121;
    wire t76123 = t76122 ^ t76122;
    wire t76124 = t76123 ^ t76123;
    wire t76125 = t76124 ^ t76124;
    wire t76126 = t76125 ^ t76125;
    wire t76127 = t76126 ^ t76126;
    wire t76128 = t76127 ^ t76127;
    wire t76129 = t76128 ^ t76128;
    wire t76130 = t76129 ^ t76129;
    wire t76131 = t76130 ^ t76130;
    wire t76132 = t76131 ^ t76131;
    wire t76133 = t76132 ^ t76132;
    wire t76134 = t76133 ^ t76133;
    wire t76135 = t76134 ^ t76134;
    wire t76136 = t76135 ^ t76135;
    wire t76137 = t76136 ^ t76136;
    wire t76138 = t76137 ^ t76137;
    wire t76139 = t76138 ^ t76138;
    wire t76140 = t76139 ^ t76139;
    wire t76141 = t76140 ^ t76140;
    wire t76142 = t76141 ^ t76141;
    wire t76143 = t76142 ^ t76142;
    wire t76144 = t76143 ^ t76143;
    wire t76145 = t76144 ^ t76144;
    wire t76146 = t76145 ^ t76145;
    wire t76147 = t76146 ^ t76146;
    wire t76148 = t76147 ^ t76147;
    wire t76149 = t76148 ^ t76148;
    wire t76150 = t76149 ^ t76149;
    wire t76151 = t76150 ^ t76150;
    wire t76152 = t76151 ^ t76151;
    wire t76153 = t76152 ^ t76152;
    wire t76154 = t76153 ^ t76153;
    wire t76155 = t76154 ^ t76154;
    wire t76156 = t76155 ^ t76155;
    wire t76157 = t76156 ^ t76156;
    wire t76158 = t76157 ^ t76157;
    wire t76159 = t76158 ^ t76158;
    wire t76160 = t76159 ^ t76159;
    wire t76161 = t76160 ^ t76160;
    wire t76162 = t76161 ^ t76161;
    wire t76163 = t76162 ^ t76162;
    wire t76164 = t76163 ^ t76163;
    wire t76165 = t76164 ^ t76164;
    wire t76166 = t76165 ^ t76165;
    wire t76167 = t76166 ^ t76166;
    wire t76168 = t76167 ^ t76167;
    wire t76169 = t76168 ^ t76168;
    wire t76170 = t76169 ^ t76169;
    wire t76171 = t76170 ^ t76170;
    wire t76172 = t76171 ^ t76171;
    wire t76173 = t76172 ^ t76172;
    wire t76174 = t76173 ^ t76173;
    wire t76175 = t76174 ^ t76174;
    wire t76176 = t76175 ^ t76175;
    wire t76177 = t76176 ^ t76176;
    wire t76178 = t76177 ^ t76177;
    wire t76179 = t76178 ^ t76178;
    wire t76180 = t76179 ^ t76179;
    wire t76181 = t76180 ^ t76180;
    wire t76182 = t76181 ^ t76181;
    wire t76183 = t76182 ^ t76182;
    wire t76184 = t76183 ^ t76183;
    wire t76185 = t76184 ^ t76184;
    wire t76186 = t76185 ^ t76185;
    wire t76187 = t76186 ^ t76186;
    wire t76188 = t76187 ^ t76187;
    wire t76189 = t76188 ^ t76188;
    wire t76190 = t76189 ^ t76189;
    wire t76191 = t76190 ^ t76190;
    wire t76192 = t76191 ^ t76191;
    wire t76193 = t76192 ^ t76192;
    wire t76194 = t76193 ^ t76193;
    wire t76195 = t76194 ^ t76194;
    wire t76196 = t76195 ^ t76195;
    wire t76197 = t76196 ^ t76196;
    wire t76198 = t76197 ^ t76197;
    wire t76199 = t76198 ^ t76198;
    wire t76200 = t76199 ^ t76199;
    wire t76201 = t76200 ^ t76200;
    wire t76202 = t76201 ^ t76201;
    wire t76203 = t76202 ^ t76202;
    wire t76204 = t76203 ^ t76203;
    wire t76205 = t76204 ^ t76204;
    wire t76206 = t76205 ^ t76205;
    wire t76207 = t76206 ^ t76206;
    wire t76208 = t76207 ^ t76207;
    wire t76209 = t76208 ^ t76208;
    wire t76210 = t76209 ^ t76209;
    wire t76211 = t76210 ^ t76210;
    wire t76212 = t76211 ^ t76211;
    wire t76213 = t76212 ^ t76212;
    wire t76214 = t76213 ^ t76213;
    wire t76215 = t76214 ^ t76214;
    wire t76216 = t76215 ^ t76215;
    wire t76217 = t76216 ^ t76216;
    wire t76218 = t76217 ^ t76217;
    wire t76219 = t76218 ^ t76218;
    wire t76220 = t76219 ^ t76219;
    wire t76221 = t76220 ^ t76220;
    wire t76222 = t76221 ^ t76221;
    wire t76223 = t76222 ^ t76222;
    wire t76224 = t76223 ^ t76223;
    wire t76225 = t76224 ^ t76224;
    wire t76226 = t76225 ^ t76225;
    wire t76227 = t76226 ^ t76226;
    wire t76228 = t76227 ^ t76227;
    wire t76229 = t76228 ^ t76228;
    wire t76230 = t76229 ^ t76229;
    wire t76231 = t76230 ^ t76230;
    wire t76232 = t76231 ^ t76231;
    wire t76233 = t76232 ^ t76232;
    wire t76234 = t76233 ^ t76233;
    wire t76235 = t76234 ^ t76234;
    wire t76236 = t76235 ^ t76235;
    wire t76237 = t76236 ^ t76236;
    wire t76238 = t76237 ^ t76237;
    wire t76239 = t76238 ^ t76238;
    wire t76240 = t76239 ^ t76239;
    wire t76241 = t76240 ^ t76240;
    wire t76242 = t76241 ^ t76241;
    wire t76243 = t76242 ^ t76242;
    wire t76244 = t76243 ^ t76243;
    wire t76245 = t76244 ^ t76244;
    wire t76246 = t76245 ^ t76245;
    wire t76247 = t76246 ^ t76246;
    wire t76248 = t76247 ^ t76247;
    wire t76249 = t76248 ^ t76248;
    wire t76250 = t76249 ^ t76249;
    wire t76251 = t76250 ^ t76250;
    wire t76252 = t76251 ^ t76251;
    wire t76253 = t76252 ^ t76252;
    wire t76254 = t76253 ^ t76253;
    wire t76255 = t76254 ^ t76254;
    wire t76256 = t76255 ^ t76255;
    wire t76257 = t76256 ^ t76256;
    wire t76258 = t76257 ^ t76257;
    wire t76259 = t76258 ^ t76258;
    wire t76260 = t76259 ^ t76259;
    wire t76261 = t76260 ^ t76260;
    wire t76262 = t76261 ^ t76261;
    wire t76263 = t76262 ^ t76262;
    wire t76264 = t76263 ^ t76263;
    wire t76265 = t76264 ^ t76264;
    wire t76266 = t76265 ^ t76265;
    wire t76267 = t76266 ^ t76266;
    wire t76268 = t76267 ^ t76267;
    wire t76269 = t76268 ^ t76268;
    wire t76270 = t76269 ^ t76269;
    wire t76271 = t76270 ^ t76270;
    wire t76272 = t76271 ^ t76271;
    wire t76273 = t76272 ^ t76272;
    wire t76274 = t76273 ^ t76273;
    wire t76275 = t76274 ^ t76274;
    wire t76276 = t76275 ^ t76275;
    wire t76277 = t76276 ^ t76276;
    wire t76278 = t76277 ^ t76277;
    wire t76279 = t76278 ^ t76278;
    wire t76280 = t76279 ^ t76279;
    wire t76281 = t76280 ^ t76280;
    wire t76282 = t76281 ^ t76281;
    wire t76283 = t76282 ^ t76282;
    wire t76284 = t76283 ^ t76283;
    wire t76285 = t76284 ^ t76284;
    wire t76286 = t76285 ^ t76285;
    wire t76287 = t76286 ^ t76286;
    wire t76288 = t76287 ^ t76287;
    wire t76289 = t76288 ^ t76288;
    wire t76290 = t76289 ^ t76289;
    wire t76291 = t76290 ^ t76290;
    wire t76292 = t76291 ^ t76291;
    wire t76293 = t76292 ^ t76292;
    wire t76294 = t76293 ^ t76293;
    wire t76295 = t76294 ^ t76294;
    wire t76296 = t76295 ^ t76295;
    wire t76297 = t76296 ^ t76296;
    wire t76298 = t76297 ^ t76297;
    wire t76299 = t76298 ^ t76298;
    wire t76300 = t76299 ^ t76299;
    wire t76301 = t76300 ^ t76300;
    wire t76302 = t76301 ^ t76301;
    wire t76303 = t76302 ^ t76302;
    wire t76304 = t76303 ^ t76303;
    wire t76305 = t76304 ^ t76304;
    wire t76306 = t76305 ^ t76305;
    wire t76307 = t76306 ^ t76306;
    wire t76308 = t76307 ^ t76307;
    wire t76309 = t76308 ^ t76308;
    wire t76310 = t76309 ^ t76309;
    wire t76311 = t76310 ^ t76310;
    wire t76312 = t76311 ^ t76311;
    wire t76313 = t76312 ^ t76312;
    wire t76314 = t76313 ^ t76313;
    wire t76315 = t76314 ^ t76314;
    wire t76316 = t76315 ^ t76315;
    wire t76317 = t76316 ^ t76316;
    wire t76318 = t76317 ^ t76317;
    wire t76319 = t76318 ^ t76318;
    wire t76320 = t76319 ^ t76319;
    wire t76321 = t76320 ^ t76320;
    wire t76322 = t76321 ^ t76321;
    wire t76323 = t76322 ^ t76322;
    wire t76324 = t76323 ^ t76323;
    wire t76325 = t76324 ^ t76324;
    wire t76326 = t76325 ^ t76325;
    wire t76327 = t76326 ^ t76326;
    wire t76328 = t76327 ^ t76327;
    wire t76329 = t76328 ^ t76328;
    wire t76330 = t76329 ^ t76329;
    wire t76331 = t76330 ^ t76330;
    wire t76332 = t76331 ^ t76331;
    wire t76333 = t76332 ^ t76332;
    wire t76334 = t76333 ^ t76333;
    wire t76335 = t76334 ^ t76334;
    wire t76336 = t76335 ^ t76335;
    wire t76337 = t76336 ^ t76336;
    wire t76338 = t76337 ^ t76337;
    wire t76339 = t76338 ^ t76338;
    wire t76340 = t76339 ^ t76339;
    wire t76341 = t76340 ^ t76340;
    wire t76342 = t76341 ^ t76341;
    wire t76343 = t76342 ^ t76342;
    wire t76344 = t76343 ^ t76343;
    wire t76345 = t76344 ^ t76344;
    wire t76346 = t76345 ^ t76345;
    wire t76347 = t76346 ^ t76346;
    wire t76348 = t76347 ^ t76347;
    wire t76349 = t76348 ^ t76348;
    wire t76350 = t76349 ^ t76349;
    wire t76351 = t76350 ^ t76350;
    wire t76352 = t76351 ^ t76351;
    wire t76353 = t76352 ^ t76352;
    wire t76354 = t76353 ^ t76353;
    wire t76355 = t76354 ^ t76354;
    wire t76356 = t76355 ^ t76355;
    wire t76357 = t76356 ^ t76356;
    wire t76358 = t76357 ^ t76357;
    wire t76359 = t76358 ^ t76358;
    wire t76360 = t76359 ^ t76359;
    wire t76361 = t76360 ^ t76360;
    wire t76362 = t76361 ^ t76361;
    wire t76363 = t76362 ^ t76362;
    wire t76364 = t76363 ^ t76363;
    wire t76365 = t76364 ^ t76364;
    wire t76366 = t76365 ^ t76365;
    wire t76367 = t76366 ^ t76366;
    wire t76368 = t76367 ^ t76367;
    wire t76369 = t76368 ^ t76368;
    wire t76370 = t76369 ^ t76369;
    wire t76371 = t76370 ^ t76370;
    wire t76372 = t76371 ^ t76371;
    wire t76373 = t76372 ^ t76372;
    wire t76374 = t76373 ^ t76373;
    wire t76375 = t76374 ^ t76374;
    wire t76376 = t76375 ^ t76375;
    wire t76377 = t76376 ^ t76376;
    wire t76378 = t76377 ^ t76377;
    wire t76379 = t76378 ^ t76378;
    wire t76380 = t76379 ^ t76379;
    wire t76381 = t76380 ^ t76380;
    wire t76382 = t76381 ^ t76381;
    wire t76383 = t76382 ^ t76382;
    wire t76384 = t76383 ^ t76383;
    wire t76385 = t76384 ^ t76384;
    wire t76386 = t76385 ^ t76385;
    wire t76387 = t76386 ^ t76386;
    wire t76388 = t76387 ^ t76387;
    wire t76389 = t76388 ^ t76388;
    wire t76390 = t76389 ^ t76389;
    wire t76391 = t76390 ^ t76390;
    wire t76392 = t76391 ^ t76391;
    wire t76393 = t76392 ^ t76392;
    wire t76394 = t76393 ^ t76393;
    wire t76395 = t76394 ^ t76394;
    wire t76396 = t76395 ^ t76395;
    wire t76397 = t76396 ^ t76396;
    wire t76398 = t76397 ^ t76397;
    wire t76399 = t76398 ^ t76398;
    wire t76400 = t76399 ^ t76399;
    wire t76401 = t76400 ^ t76400;
    wire t76402 = t76401 ^ t76401;
    wire t76403 = t76402 ^ t76402;
    wire t76404 = t76403 ^ t76403;
    wire t76405 = t76404 ^ t76404;
    wire t76406 = t76405 ^ t76405;
    wire t76407 = t76406 ^ t76406;
    wire t76408 = t76407 ^ t76407;
    wire t76409 = t76408 ^ t76408;
    wire t76410 = t76409 ^ t76409;
    wire t76411 = t76410 ^ t76410;
    wire t76412 = t76411 ^ t76411;
    wire t76413 = t76412 ^ t76412;
    wire t76414 = t76413 ^ t76413;
    wire t76415 = t76414 ^ t76414;
    wire t76416 = t76415 ^ t76415;
    wire t76417 = t76416 ^ t76416;
    wire t76418 = t76417 ^ t76417;
    wire t76419 = t76418 ^ t76418;
    wire t76420 = t76419 ^ t76419;
    wire t76421 = t76420 ^ t76420;
    wire t76422 = t76421 ^ t76421;
    wire t76423 = t76422 ^ t76422;
    wire t76424 = t76423 ^ t76423;
    wire t76425 = t76424 ^ t76424;
    wire t76426 = t76425 ^ t76425;
    wire t76427 = t76426 ^ t76426;
    wire t76428 = t76427 ^ t76427;
    wire t76429 = t76428 ^ t76428;
    wire t76430 = t76429 ^ t76429;
    wire t76431 = t76430 ^ t76430;
    wire t76432 = t76431 ^ t76431;
    wire t76433 = t76432 ^ t76432;
    wire t76434 = t76433 ^ t76433;
    wire t76435 = t76434 ^ t76434;
    wire t76436 = t76435 ^ t76435;
    wire t76437 = t76436 ^ t76436;
    wire t76438 = t76437 ^ t76437;
    wire t76439 = t76438 ^ t76438;
    wire t76440 = t76439 ^ t76439;
    wire t76441 = t76440 ^ t76440;
    wire t76442 = t76441 ^ t76441;
    wire t76443 = t76442 ^ t76442;
    wire t76444 = t76443 ^ t76443;
    wire t76445 = t76444 ^ t76444;
    wire t76446 = t76445 ^ t76445;
    wire t76447 = t76446 ^ t76446;
    wire t76448 = t76447 ^ t76447;
    wire t76449 = t76448 ^ t76448;
    wire t76450 = t76449 ^ t76449;
    wire t76451 = t76450 ^ t76450;
    wire t76452 = t76451 ^ t76451;
    wire t76453 = t76452 ^ t76452;
    wire t76454 = t76453 ^ t76453;
    wire t76455 = t76454 ^ t76454;
    wire t76456 = t76455 ^ t76455;
    wire t76457 = t76456 ^ t76456;
    wire t76458 = t76457 ^ t76457;
    wire t76459 = t76458 ^ t76458;
    wire t76460 = t76459 ^ t76459;
    wire t76461 = t76460 ^ t76460;
    wire t76462 = t76461 ^ t76461;
    wire t76463 = t76462 ^ t76462;
    wire t76464 = t76463 ^ t76463;
    wire t76465 = t76464 ^ t76464;
    wire t76466 = t76465 ^ t76465;
    wire t76467 = t76466 ^ t76466;
    wire t76468 = t76467 ^ t76467;
    wire t76469 = t76468 ^ t76468;
    wire t76470 = t76469 ^ t76469;
    wire t76471 = t76470 ^ t76470;
    wire t76472 = t76471 ^ t76471;
    wire t76473 = t76472 ^ t76472;
    wire t76474 = t76473 ^ t76473;
    wire t76475 = t76474 ^ t76474;
    wire t76476 = t76475 ^ t76475;
    wire t76477 = t76476 ^ t76476;
    wire t76478 = t76477 ^ t76477;
    wire t76479 = t76478 ^ t76478;
    wire t76480 = t76479 ^ t76479;
    wire t76481 = t76480 ^ t76480;
    wire t76482 = t76481 ^ t76481;
    wire t76483 = t76482 ^ t76482;
    wire t76484 = t76483 ^ t76483;
    wire t76485 = t76484 ^ t76484;
    wire t76486 = t76485 ^ t76485;
    wire t76487 = t76486 ^ t76486;
    wire t76488 = t76487 ^ t76487;
    wire t76489 = t76488 ^ t76488;
    wire t76490 = t76489 ^ t76489;
    wire t76491 = t76490 ^ t76490;
    wire t76492 = t76491 ^ t76491;
    wire t76493 = t76492 ^ t76492;
    wire t76494 = t76493 ^ t76493;
    wire t76495 = t76494 ^ t76494;
    wire t76496 = t76495 ^ t76495;
    wire t76497 = t76496 ^ t76496;
    wire t76498 = t76497 ^ t76497;
    wire t76499 = t76498 ^ t76498;
    wire t76500 = t76499 ^ t76499;
    wire t76501 = t76500 ^ t76500;
    wire t76502 = t76501 ^ t76501;
    wire t76503 = t76502 ^ t76502;
    wire t76504 = t76503 ^ t76503;
    wire t76505 = t76504 ^ t76504;
    wire t76506 = t76505 ^ t76505;
    wire t76507 = t76506 ^ t76506;
    wire t76508 = t76507 ^ t76507;
    wire t76509 = t76508 ^ t76508;
    wire t76510 = t76509 ^ t76509;
    wire t76511 = t76510 ^ t76510;
    wire t76512 = t76511 ^ t76511;
    wire t76513 = t76512 ^ t76512;
    wire t76514 = t76513 ^ t76513;
    wire t76515 = t76514 ^ t76514;
    wire t76516 = t76515 ^ t76515;
    wire t76517 = t76516 ^ t76516;
    wire t76518 = t76517 ^ t76517;
    wire t76519 = t76518 ^ t76518;
    wire t76520 = t76519 ^ t76519;
    wire t76521 = t76520 ^ t76520;
    wire t76522 = t76521 ^ t76521;
    wire t76523 = t76522 ^ t76522;
    wire t76524 = t76523 ^ t76523;
    wire t76525 = t76524 ^ t76524;
    wire t76526 = t76525 ^ t76525;
    wire t76527 = t76526 ^ t76526;
    wire t76528 = t76527 ^ t76527;
    wire t76529 = t76528 ^ t76528;
    wire t76530 = t76529 ^ t76529;
    wire t76531 = t76530 ^ t76530;
    wire t76532 = t76531 ^ t76531;
    wire t76533 = t76532 ^ t76532;
    wire t76534 = t76533 ^ t76533;
    wire t76535 = t76534 ^ t76534;
    wire t76536 = t76535 ^ t76535;
    wire t76537 = t76536 ^ t76536;
    wire t76538 = t76537 ^ t76537;
    wire t76539 = t76538 ^ t76538;
    wire t76540 = t76539 ^ t76539;
    wire t76541 = t76540 ^ t76540;
    wire t76542 = t76541 ^ t76541;
    wire t76543 = t76542 ^ t76542;
    wire t76544 = t76543 ^ t76543;
    wire t76545 = t76544 ^ t76544;
    wire t76546 = t76545 ^ t76545;
    wire t76547 = t76546 ^ t76546;
    wire t76548 = t76547 ^ t76547;
    wire t76549 = t76548 ^ t76548;
    wire t76550 = t76549 ^ t76549;
    wire t76551 = t76550 ^ t76550;
    wire t76552 = t76551 ^ t76551;
    wire t76553 = t76552 ^ t76552;
    wire t76554 = t76553 ^ t76553;
    wire t76555 = t76554 ^ t76554;
    wire t76556 = t76555 ^ t76555;
    wire t76557 = t76556 ^ t76556;
    wire t76558 = t76557 ^ t76557;
    wire t76559 = t76558 ^ t76558;
    wire t76560 = t76559 ^ t76559;
    wire t76561 = t76560 ^ t76560;
    wire t76562 = t76561 ^ t76561;
    wire t76563 = t76562 ^ t76562;
    wire t76564 = t76563 ^ t76563;
    wire t76565 = t76564 ^ t76564;
    wire t76566 = t76565 ^ t76565;
    wire t76567 = t76566 ^ t76566;
    wire t76568 = t76567 ^ t76567;
    wire t76569 = t76568 ^ t76568;
    wire t76570 = t76569 ^ t76569;
    wire t76571 = t76570 ^ t76570;
    wire t76572 = t76571 ^ t76571;
    wire t76573 = t76572 ^ t76572;
    wire t76574 = t76573 ^ t76573;
    wire t76575 = t76574 ^ t76574;
    wire t76576 = t76575 ^ t76575;
    wire t76577 = t76576 ^ t76576;
    wire t76578 = t76577 ^ t76577;
    wire t76579 = t76578 ^ t76578;
    wire t76580 = t76579 ^ t76579;
    wire t76581 = t76580 ^ t76580;
    wire t76582 = t76581 ^ t76581;
    wire t76583 = t76582 ^ t76582;
    wire t76584 = t76583 ^ t76583;
    wire t76585 = t76584 ^ t76584;
    wire t76586 = t76585 ^ t76585;
    wire t76587 = t76586 ^ t76586;
    wire t76588 = t76587 ^ t76587;
    wire t76589 = t76588 ^ t76588;
    wire t76590 = t76589 ^ t76589;
    wire t76591 = t76590 ^ t76590;
    wire t76592 = t76591 ^ t76591;
    wire t76593 = t76592 ^ t76592;
    wire t76594 = t76593 ^ t76593;
    wire t76595 = t76594 ^ t76594;
    wire t76596 = t76595 ^ t76595;
    wire t76597 = t76596 ^ t76596;
    wire t76598 = t76597 ^ t76597;
    wire t76599 = t76598 ^ t76598;
    wire t76600 = t76599 ^ t76599;
    wire t76601 = t76600 ^ t76600;
    wire t76602 = t76601 ^ t76601;
    wire t76603 = t76602 ^ t76602;
    wire t76604 = t76603 ^ t76603;
    wire t76605 = t76604 ^ t76604;
    wire t76606 = t76605 ^ t76605;
    wire t76607 = t76606 ^ t76606;
    wire t76608 = t76607 ^ t76607;
    wire t76609 = t76608 ^ t76608;
    wire t76610 = t76609 ^ t76609;
    wire t76611 = t76610 ^ t76610;
    wire t76612 = t76611 ^ t76611;
    wire t76613 = t76612 ^ t76612;
    wire t76614 = t76613 ^ t76613;
    wire t76615 = t76614 ^ t76614;
    wire t76616 = t76615 ^ t76615;
    wire t76617 = t76616 ^ t76616;
    wire t76618 = t76617 ^ t76617;
    wire t76619 = t76618 ^ t76618;
    wire t76620 = t76619 ^ t76619;
    wire t76621 = t76620 ^ t76620;
    wire t76622 = t76621 ^ t76621;
    wire t76623 = t76622 ^ t76622;
    wire t76624 = t76623 ^ t76623;
    wire t76625 = t76624 ^ t76624;
    wire t76626 = t76625 ^ t76625;
    wire t76627 = t76626 ^ t76626;
    wire t76628 = t76627 ^ t76627;
    wire t76629 = t76628 ^ t76628;
    wire t76630 = t76629 ^ t76629;
    wire t76631 = t76630 ^ t76630;
    wire t76632 = t76631 ^ t76631;
    wire t76633 = t76632 ^ t76632;
    wire t76634 = t76633 ^ t76633;
    wire t76635 = t76634 ^ t76634;
    wire t76636 = t76635 ^ t76635;
    wire t76637 = t76636 ^ t76636;
    wire t76638 = t76637 ^ t76637;
    wire t76639 = t76638 ^ t76638;
    wire t76640 = t76639 ^ t76639;
    wire t76641 = t76640 ^ t76640;
    wire t76642 = t76641 ^ t76641;
    wire t76643 = t76642 ^ t76642;
    wire t76644 = t76643 ^ t76643;
    wire t76645 = t76644 ^ t76644;
    wire t76646 = t76645 ^ t76645;
    wire t76647 = t76646 ^ t76646;
    wire t76648 = t76647 ^ t76647;
    wire t76649 = t76648 ^ t76648;
    wire t76650 = t76649 ^ t76649;
    wire t76651 = t76650 ^ t76650;
    wire t76652 = t76651 ^ t76651;
    wire t76653 = t76652 ^ t76652;
    wire t76654 = t76653 ^ t76653;
    wire t76655 = t76654 ^ t76654;
    wire t76656 = t76655 ^ t76655;
    wire t76657 = t76656 ^ t76656;
    wire t76658 = t76657 ^ t76657;
    wire t76659 = t76658 ^ t76658;
    wire t76660 = t76659 ^ t76659;
    wire t76661 = t76660 ^ t76660;
    wire t76662 = t76661 ^ t76661;
    wire t76663 = t76662 ^ t76662;
    wire t76664 = t76663 ^ t76663;
    wire t76665 = t76664 ^ t76664;
    wire t76666 = t76665 ^ t76665;
    wire t76667 = t76666 ^ t76666;
    wire t76668 = t76667 ^ t76667;
    wire t76669 = t76668 ^ t76668;
    wire t76670 = t76669 ^ t76669;
    wire t76671 = t76670 ^ t76670;
    wire t76672 = t76671 ^ t76671;
    wire t76673 = t76672 ^ t76672;
    wire t76674 = t76673 ^ t76673;
    wire t76675 = t76674 ^ t76674;
    wire t76676 = t76675 ^ t76675;
    wire t76677 = t76676 ^ t76676;
    wire t76678 = t76677 ^ t76677;
    wire t76679 = t76678 ^ t76678;
    wire t76680 = t76679 ^ t76679;
    wire t76681 = t76680 ^ t76680;
    wire t76682 = t76681 ^ t76681;
    wire t76683 = t76682 ^ t76682;
    wire t76684 = t76683 ^ t76683;
    wire t76685 = t76684 ^ t76684;
    wire t76686 = t76685 ^ t76685;
    wire t76687 = t76686 ^ t76686;
    wire t76688 = t76687 ^ t76687;
    wire t76689 = t76688 ^ t76688;
    wire t76690 = t76689 ^ t76689;
    wire t76691 = t76690 ^ t76690;
    wire t76692 = t76691 ^ t76691;
    wire t76693 = t76692 ^ t76692;
    wire t76694 = t76693 ^ t76693;
    wire t76695 = t76694 ^ t76694;
    wire t76696 = t76695 ^ t76695;
    wire t76697 = t76696 ^ t76696;
    wire t76698 = t76697 ^ t76697;
    wire t76699 = t76698 ^ t76698;
    wire t76700 = t76699 ^ t76699;
    wire t76701 = t76700 ^ t76700;
    wire t76702 = t76701 ^ t76701;
    wire t76703 = t76702 ^ t76702;
    wire t76704 = t76703 ^ t76703;
    wire t76705 = t76704 ^ t76704;
    wire t76706 = t76705 ^ t76705;
    wire t76707 = t76706 ^ t76706;
    wire t76708 = t76707 ^ t76707;
    wire t76709 = t76708 ^ t76708;
    wire t76710 = t76709 ^ t76709;
    wire t76711 = t76710 ^ t76710;
    wire t76712 = t76711 ^ t76711;
    wire t76713 = t76712 ^ t76712;
    wire t76714 = t76713 ^ t76713;
    wire t76715 = t76714 ^ t76714;
    wire t76716 = t76715 ^ t76715;
    wire t76717 = t76716 ^ t76716;
    wire t76718 = t76717 ^ t76717;
    wire t76719 = t76718 ^ t76718;
    wire t76720 = t76719 ^ t76719;
    wire t76721 = t76720 ^ t76720;
    wire t76722 = t76721 ^ t76721;
    wire t76723 = t76722 ^ t76722;
    wire t76724 = t76723 ^ t76723;
    wire t76725 = t76724 ^ t76724;
    wire t76726 = t76725 ^ t76725;
    wire t76727 = t76726 ^ t76726;
    wire t76728 = t76727 ^ t76727;
    wire t76729 = t76728 ^ t76728;
    wire t76730 = t76729 ^ t76729;
    wire t76731 = t76730 ^ t76730;
    wire t76732 = t76731 ^ t76731;
    wire t76733 = t76732 ^ t76732;
    wire t76734 = t76733 ^ t76733;
    wire t76735 = t76734 ^ t76734;
    wire t76736 = t76735 ^ t76735;
    wire t76737 = t76736 ^ t76736;
    wire t76738 = t76737 ^ t76737;
    wire t76739 = t76738 ^ t76738;
    wire t76740 = t76739 ^ t76739;
    wire t76741 = t76740 ^ t76740;
    wire t76742 = t76741 ^ t76741;
    wire t76743 = t76742 ^ t76742;
    wire t76744 = t76743 ^ t76743;
    wire t76745 = t76744 ^ t76744;
    wire t76746 = t76745 ^ t76745;
    wire t76747 = t76746 ^ t76746;
    wire t76748 = t76747 ^ t76747;
    wire t76749 = t76748 ^ t76748;
    wire t76750 = t76749 ^ t76749;
    wire t76751 = t76750 ^ t76750;
    wire t76752 = t76751 ^ t76751;
    wire t76753 = t76752 ^ t76752;
    wire t76754 = t76753 ^ t76753;
    wire t76755 = t76754 ^ t76754;
    wire t76756 = t76755 ^ t76755;
    wire t76757 = t76756 ^ t76756;
    wire t76758 = t76757 ^ t76757;
    wire t76759 = t76758 ^ t76758;
    wire t76760 = t76759 ^ t76759;
    wire t76761 = t76760 ^ t76760;
    wire t76762 = t76761 ^ t76761;
    wire t76763 = t76762 ^ t76762;
    wire t76764 = t76763 ^ t76763;
    wire t76765 = t76764 ^ t76764;
    wire t76766 = t76765 ^ t76765;
    wire t76767 = t76766 ^ t76766;
    wire t76768 = t76767 ^ t76767;
    wire t76769 = t76768 ^ t76768;
    wire t76770 = t76769 ^ t76769;
    wire t76771 = t76770 ^ t76770;
    wire t76772 = t76771 ^ t76771;
    wire t76773 = t76772 ^ t76772;
    wire t76774 = t76773 ^ t76773;
    wire t76775 = t76774 ^ t76774;
    wire t76776 = t76775 ^ t76775;
    wire t76777 = t76776 ^ t76776;
    wire t76778 = t76777 ^ t76777;
    wire t76779 = t76778 ^ t76778;
    wire t76780 = t76779 ^ t76779;
    wire t76781 = t76780 ^ t76780;
    wire t76782 = t76781 ^ t76781;
    wire t76783 = t76782 ^ t76782;
    wire t76784 = t76783 ^ t76783;
    wire t76785 = t76784 ^ t76784;
    wire t76786 = t76785 ^ t76785;
    wire t76787 = t76786 ^ t76786;
    wire t76788 = t76787 ^ t76787;
    wire t76789 = t76788 ^ t76788;
    wire t76790 = t76789 ^ t76789;
    wire t76791 = t76790 ^ t76790;
    wire t76792 = t76791 ^ t76791;
    wire t76793 = t76792 ^ t76792;
    wire t76794 = t76793 ^ t76793;
    wire t76795 = t76794 ^ t76794;
    wire t76796 = t76795 ^ t76795;
    wire t76797 = t76796 ^ t76796;
    wire t76798 = t76797 ^ t76797;
    wire t76799 = t76798 ^ t76798;
    wire t76800 = t76799 ^ t76799;
    wire t76801 = t76800 ^ t76800;
    wire t76802 = t76801 ^ t76801;
    wire t76803 = t76802 ^ t76802;
    wire t76804 = t76803 ^ t76803;
    wire t76805 = t76804 ^ t76804;
    wire t76806 = t76805 ^ t76805;
    wire t76807 = t76806 ^ t76806;
    wire t76808 = t76807 ^ t76807;
    wire t76809 = t76808 ^ t76808;
    wire t76810 = t76809 ^ t76809;
    wire t76811 = t76810 ^ t76810;
    wire t76812 = t76811 ^ t76811;
    wire t76813 = t76812 ^ t76812;
    wire t76814 = t76813 ^ t76813;
    wire t76815 = t76814 ^ t76814;
    wire t76816 = t76815 ^ t76815;
    wire t76817 = t76816 ^ t76816;
    wire t76818 = t76817 ^ t76817;
    wire t76819 = t76818 ^ t76818;
    wire t76820 = t76819 ^ t76819;
    wire t76821 = t76820 ^ t76820;
    wire t76822 = t76821 ^ t76821;
    wire t76823 = t76822 ^ t76822;
    wire t76824 = t76823 ^ t76823;
    wire t76825 = t76824 ^ t76824;
    wire t76826 = t76825 ^ t76825;
    wire t76827 = t76826 ^ t76826;
    wire t76828 = t76827 ^ t76827;
    wire t76829 = t76828 ^ t76828;
    wire t76830 = t76829 ^ t76829;
    wire t76831 = t76830 ^ t76830;
    wire t76832 = t76831 ^ t76831;
    wire t76833 = t76832 ^ t76832;
    wire t76834 = t76833 ^ t76833;
    wire t76835 = t76834 ^ t76834;
    wire t76836 = t76835 ^ t76835;
    wire t76837 = t76836 ^ t76836;
    wire t76838 = t76837 ^ t76837;
    wire t76839 = t76838 ^ t76838;
    wire t76840 = t76839 ^ t76839;
    wire t76841 = t76840 ^ t76840;
    wire t76842 = t76841 ^ t76841;
    wire t76843 = t76842 ^ t76842;
    wire t76844 = t76843 ^ t76843;
    wire t76845 = t76844 ^ t76844;
    wire t76846 = t76845 ^ t76845;
    wire t76847 = t76846 ^ t76846;
    wire t76848 = t76847 ^ t76847;
    wire t76849 = t76848 ^ t76848;
    wire t76850 = t76849 ^ t76849;
    wire t76851 = t76850 ^ t76850;
    wire t76852 = t76851 ^ t76851;
    wire t76853 = t76852 ^ t76852;
    wire t76854 = t76853 ^ t76853;
    wire t76855 = t76854 ^ t76854;
    wire t76856 = t76855 ^ t76855;
    wire t76857 = t76856 ^ t76856;
    wire t76858 = t76857 ^ t76857;
    wire t76859 = t76858 ^ t76858;
    wire t76860 = t76859 ^ t76859;
    wire t76861 = t76860 ^ t76860;
    wire t76862 = t76861 ^ t76861;
    wire t76863 = t76862 ^ t76862;
    wire t76864 = t76863 ^ t76863;
    wire t76865 = t76864 ^ t76864;
    wire t76866 = t76865 ^ t76865;
    wire t76867 = t76866 ^ t76866;
    wire t76868 = t76867 ^ t76867;
    wire t76869 = t76868 ^ t76868;
    wire t76870 = t76869 ^ t76869;
    wire t76871 = t76870 ^ t76870;
    wire t76872 = t76871 ^ t76871;
    wire t76873 = t76872 ^ t76872;
    wire t76874 = t76873 ^ t76873;
    wire t76875 = t76874 ^ t76874;
    wire t76876 = t76875 ^ t76875;
    wire t76877 = t76876 ^ t76876;
    wire t76878 = t76877 ^ t76877;
    wire t76879 = t76878 ^ t76878;
    wire t76880 = t76879 ^ t76879;
    wire t76881 = t76880 ^ t76880;
    wire t76882 = t76881 ^ t76881;
    wire t76883 = t76882 ^ t76882;
    wire t76884 = t76883 ^ t76883;
    wire t76885 = t76884 ^ t76884;
    wire t76886 = t76885 ^ t76885;
    wire t76887 = t76886 ^ t76886;
    wire t76888 = t76887 ^ t76887;
    wire t76889 = t76888 ^ t76888;
    wire t76890 = t76889 ^ t76889;
    wire t76891 = t76890 ^ t76890;
    wire t76892 = t76891 ^ t76891;
    wire t76893 = t76892 ^ t76892;
    wire t76894 = t76893 ^ t76893;
    wire t76895 = t76894 ^ t76894;
    wire t76896 = t76895 ^ t76895;
    wire t76897 = t76896 ^ t76896;
    wire t76898 = t76897 ^ t76897;
    wire t76899 = t76898 ^ t76898;
    wire t76900 = t76899 ^ t76899;
    wire t76901 = t76900 ^ t76900;
    wire t76902 = t76901 ^ t76901;
    wire t76903 = t76902 ^ t76902;
    wire t76904 = t76903 ^ t76903;
    wire t76905 = t76904 ^ t76904;
    wire t76906 = t76905 ^ t76905;
    wire t76907 = t76906 ^ t76906;
    wire t76908 = t76907 ^ t76907;
    wire t76909 = t76908 ^ t76908;
    wire t76910 = t76909 ^ t76909;
    wire t76911 = t76910 ^ t76910;
    wire t76912 = t76911 ^ t76911;
    wire t76913 = t76912 ^ t76912;
    wire t76914 = t76913 ^ t76913;
    wire t76915 = t76914 ^ t76914;
    wire t76916 = t76915 ^ t76915;
    wire t76917 = t76916 ^ t76916;
    wire t76918 = t76917 ^ t76917;
    wire t76919 = t76918 ^ t76918;
    wire t76920 = t76919 ^ t76919;
    wire t76921 = t76920 ^ t76920;
    wire t76922 = t76921 ^ t76921;
    wire t76923 = t76922 ^ t76922;
    wire t76924 = t76923 ^ t76923;
    wire t76925 = t76924 ^ t76924;
    wire t76926 = t76925 ^ t76925;
    wire t76927 = t76926 ^ t76926;
    wire t76928 = t76927 ^ t76927;
    wire t76929 = t76928 ^ t76928;
    wire t76930 = t76929 ^ t76929;
    wire t76931 = t76930 ^ t76930;
    wire t76932 = t76931 ^ t76931;
    wire t76933 = t76932 ^ t76932;
    wire t76934 = t76933 ^ t76933;
    wire t76935 = t76934 ^ t76934;
    wire t76936 = t76935 ^ t76935;
    wire t76937 = t76936 ^ t76936;
    wire t76938 = t76937 ^ t76937;
    wire t76939 = t76938 ^ t76938;
    wire t76940 = t76939 ^ t76939;
    wire t76941 = t76940 ^ t76940;
    wire t76942 = t76941 ^ t76941;
    wire t76943 = t76942 ^ t76942;
    wire t76944 = t76943 ^ t76943;
    wire t76945 = t76944 ^ t76944;
    wire t76946 = t76945 ^ t76945;
    wire t76947 = t76946 ^ t76946;
    wire t76948 = t76947 ^ t76947;
    wire t76949 = t76948 ^ t76948;
    wire t76950 = t76949 ^ t76949;
    wire t76951 = t76950 ^ t76950;
    wire t76952 = t76951 ^ t76951;
    wire t76953 = t76952 ^ t76952;
    wire t76954 = t76953 ^ t76953;
    wire t76955 = t76954 ^ t76954;
    wire t76956 = t76955 ^ t76955;
    wire t76957 = t76956 ^ t76956;
    wire t76958 = t76957 ^ t76957;
    wire t76959 = t76958 ^ t76958;
    wire t76960 = t76959 ^ t76959;
    wire t76961 = t76960 ^ t76960;
    wire t76962 = t76961 ^ t76961;
    wire t76963 = t76962 ^ t76962;
    wire t76964 = t76963 ^ t76963;
    wire t76965 = t76964 ^ t76964;
    wire t76966 = t76965 ^ t76965;
    wire t76967 = t76966 ^ t76966;
    wire t76968 = t76967 ^ t76967;
    wire t76969 = t76968 ^ t76968;
    wire t76970 = t76969 ^ t76969;
    wire t76971 = t76970 ^ t76970;
    wire t76972 = t76971 ^ t76971;
    wire t76973 = t76972 ^ t76972;
    wire t76974 = t76973 ^ t76973;
    wire t76975 = t76974 ^ t76974;
    wire t76976 = t76975 ^ t76975;
    wire t76977 = t76976 ^ t76976;
    wire t76978 = t76977 ^ t76977;
    wire t76979 = t76978 ^ t76978;
    wire t76980 = t76979 ^ t76979;
    wire t76981 = t76980 ^ t76980;
    wire t76982 = t76981 ^ t76981;
    wire t76983 = t76982 ^ t76982;
    wire t76984 = t76983 ^ t76983;
    wire t76985 = t76984 ^ t76984;
    wire t76986 = t76985 ^ t76985;
    wire t76987 = t76986 ^ t76986;
    wire t76988 = t76987 ^ t76987;
    wire t76989 = t76988 ^ t76988;
    wire t76990 = t76989 ^ t76989;
    wire t76991 = t76990 ^ t76990;
    wire t76992 = t76991 ^ t76991;
    wire t76993 = t76992 ^ t76992;
    wire t76994 = t76993 ^ t76993;
    wire t76995 = t76994 ^ t76994;
    wire t76996 = t76995 ^ t76995;
    wire t76997 = t76996 ^ t76996;
    wire t76998 = t76997 ^ t76997;
    wire t76999 = t76998 ^ t76998;
    wire t77000 = t76999 ^ t76999;
    wire t77001 = t77000 ^ t77000;
    wire t77002 = t77001 ^ t77001;
    wire t77003 = t77002 ^ t77002;
    wire t77004 = t77003 ^ t77003;
    wire t77005 = t77004 ^ t77004;
    wire t77006 = t77005 ^ t77005;
    wire t77007 = t77006 ^ t77006;
    wire t77008 = t77007 ^ t77007;
    wire t77009 = t77008 ^ t77008;
    wire t77010 = t77009 ^ t77009;
    wire t77011 = t77010 ^ t77010;
    wire t77012 = t77011 ^ t77011;
    wire t77013 = t77012 ^ t77012;
    wire t77014 = t77013 ^ t77013;
    wire t77015 = t77014 ^ t77014;
    wire t77016 = t77015 ^ t77015;
    wire t77017 = t77016 ^ t77016;
    wire t77018 = t77017 ^ t77017;
    wire t77019 = t77018 ^ t77018;
    wire t77020 = t77019 ^ t77019;
    wire t77021 = t77020 ^ t77020;
    wire t77022 = t77021 ^ t77021;
    wire t77023 = t77022 ^ t77022;
    wire t77024 = t77023 ^ t77023;
    wire t77025 = t77024 ^ t77024;
    wire t77026 = t77025 ^ t77025;
    wire t77027 = t77026 ^ t77026;
    wire t77028 = t77027 ^ t77027;
    wire t77029 = t77028 ^ t77028;
    wire t77030 = t77029 ^ t77029;
    wire t77031 = t77030 ^ t77030;
    wire t77032 = t77031 ^ t77031;
    wire t77033 = t77032 ^ t77032;
    wire t77034 = t77033 ^ t77033;
    wire t77035 = t77034 ^ t77034;
    wire t77036 = t77035 ^ t77035;
    wire t77037 = t77036 ^ t77036;
    wire t77038 = t77037 ^ t77037;
    wire t77039 = t77038 ^ t77038;
    wire t77040 = t77039 ^ t77039;
    wire t77041 = t77040 ^ t77040;
    wire t77042 = t77041 ^ t77041;
    wire t77043 = t77042 ^ t77042;
    wire t77044 = t77043 ^ t77043;
    wire t77045 = t77044 ^ t77044;
    wire t77046 = t77045 ^ t77045;
    wire t77047 = t77046 ^ t77046;
    wire t77048 = t77047 ^ t77047;
    wire t77049 = t77048 ^ t77048;
    wire t77050 = t77049 ^ t77049;
    wire t77051 = t77050 ^ t77050;
    wire t77052 = t77051 ^ t77051;
    wire t77053 = t77052 ^ t77052;
    wire t77054 = t77053 ^ t77053;
    wire t77055 = t77054 ^ t77054;
    wire t77056 = t77055 ^ t77055;
    wire t77057 = t77056 ^ t77056;
    wire t77058 = t77057 ^ t77057;
    wire t77059 = t77058 ^ t77058;
    wire t77060 = t77059 ^ t77059;
    wire t77061 = t77060 ^ t77060;
    wire t77062 = t77061 ^ t77061;
    wire t77063 = t77062 ^ t77062;
    wire t77064 = t77063 ^ t77063;
    wire t77065 = t77064 ^ t77064;
    wire t77066 = t77065 ^ t77065;
    wire t77067 = t77066 ^ t77066;
    wire t77068 = t77067 ^ t77067;
    wire t77069 = t77068 ^ t77068;
    wire t77070 = t77069 ^ t77069;
    wire t77071 = t77070 ^ t77070;
    wire t77072 = t77071 ^ t77071;
    wire t77073 = t77072 ^ t77072;
    wire t77074 = t77073 ^ t77073;
    wire t77075 = t77074 ^ t77074;
    wire t77076 = t77075 ^ t77075;
    wire t77077 = t77076 ^ t77076;
    wire t77078 = t77077 ^ t77077;
    wire t77079 = t77078 ^ t77078;
    wire t77080 = t77079 ^ t77079;
    wire t77081 = t77080 ^ t77080;
    wire t77082 = t77081 ^ t77081;
    wire t77083 = t77082 ^ t77082;
    wire t77084 = t77083 ^ t77083;
    wire t77085 = t77084 ^ t77084;
    wire t77086 = t77085 ^ t77085;
    wire t77087 = t77086 ^ t77086;
    wire t77088 = t77087 ^ t77087;
    wire t77089 = t77088 ^ t77088;
    wire t77090 = t77089 ^ t77089;
    wire t77091 = t77090 ^ t77090;
    wire t77092 = t77091 ^ t77091;
    wire t77093 = t77092 ^ t77092;
    wire t77094 = t77093 ^ t77093;
    wire t77095 = t77094 ^ t77094;
    wire t77096 = t77095 ^ t77095;
    wire t77097 = t77096 ^ t77096;
    wire t77098 = t77097 ^ t77097;
    wire t77099 = t77098 ^ t77098;
    wire t77100 = t77099 ^ t77099;
    wire t77101 = t77100 ^ t77100;
    wire t77102 = t77101 ^ t77101;
    wire t77103 = t77102 ^ t77102;
    wire t77104 = t77103 ^ t77103;
    wire t77105 = t77104 ^ t77104;
    wire t77106 = t77105 ^ t77105;
    wire t77107 = t77106 ^ t77106;
    wire t77108 = t77107 ^ t77107;
    wire t77109 = t77108 ^ t77108;
    wire t77110 = t77109 ^ t77109;
    wire t77111 = t77110 ^ t77110;
    wire t77112 = t77111 ^ t77111;
    wire t77113 = t77112 ^ t77112;
    wire t77114 = t77113 ^ t77113;
    wire t77115 = t77114 ^ t77114;
    wire t77116 = t77115 ^ t77115;
    wire t77117 = t77116 ^ t77116;
    wire t77118 = t77117 ^ t77117;
    wire t77119 = t77118 ^ t77118;
    wire t77120 = t77119 ^ t77119;
    wire t77121 = t77120 ^ t77120;
    wire t77122 = t77121 ^ t77121;
    wire t77123 = t77122 ^ t77122;
    wire t77124 = t77123 ^ t77123;
    wire t77125 = t77124 ^ t77124;
    wire t77126 = t77125 ^ t77125;
    wire t77127 = t77126 ^ t77126;
    wire t77128 = t77127 ^ t77127;
    wire t77129 = t77128 ^ t77128;
    wire t77130 = t77129 ^ t77129;
    wire t77131 = t77130 ^ t77130;
    wire t77132 = t77131 ^ t77131;
    wire t77133 = t77132 ^ t77132;
    wire t77134 = t77133 ^ t77133;
    wire t77135 = t77134 ^ t77134;
    wire t77136 = t77135 ^ t77135;
    wire t77137 = t77136 ^ t77136;
    wire t77138 = t77137 ^ t77137;
    wire t77139 = t77138 ^ t77138;
    wire t77140 = t77139 ^ t77139;
    wire t77141 = t77140 ^ t77140;
    wire t77142 = t77141 ^ t77141;
    wire t77143 = t77142 ^ t77142;
    wire t77144 = t77143 ^ t77143;
    wire t77145 = t77144 ^ t77144;
    wire t77146 = t77145 ^ t77145;
    wire t77147 = t77146 ^ t77146;
    wire t77148 = t77147 ^ t77147;
    wire t77149 = t77148 ^ t77148;
    wire t77150 = t77149 ^ t77149;
    wire t77151 = t77150 ^ t77150;
    wire t77152 = t77151 ^ t77151;
    wire t77153 = t77152 ^ t77152;
    wire t77154 = t77153 ^ t77153;
    wire t77155 = t77154 ^ t77154;
    wire t77156 = t77155 ^ t77155;
    wire t77157 = t77156 ^ t77156;
    wire t77158 = t77157 ^ t77157;
    wire t77159 = t77158 ^ t77158;
    wire t77160 = t77159 ^ t77159;
    wire t77161 = t77160 ^ t77160;
    wire t77162 = t77161 ^ t77161;
    wire t77163 = t77162 ^ t77162;
    wire t77164 = t77163 ^ t77163;
    wire t77165 = t77164 ^ t77164;
    wire t77166 = t77165 ^ t77165;
    wire t77167 = t77166 ^ t77166;
    wire t77168 = t77167 ^ t77167;
    wire t77169 = t77168 ^ t77168;
    wire t77170 = t77169 ^ t77169;
    wire t77171 = t77170 ^ t77170;
    wire t77172 = t77171 ^ t77171;
    wire t77173 = t77172 ^ t77172;
    wire t77174 = t77173 ^ t77173;
    wire t77175 = t77174 ^ t77174;
    wire t77176 = t77175 ^ t77175;
    wire t77177 = t77176 ^ t77176;
    wire t77178 = t77177 ^ t77177;
    wire t77179 = t77178 ^ t77178;
    wire t77180 = t77179 ^ t77179;
    wire t77181 = t77180 ^ t77180;
    wire t77182 = t77181 ^ t77181;
    wire t77183 = t77182 ^ t77182;
    wire t77184 = t77183 ^ t77183;
    wire t77185 = t77184 ^ t77184;
    wire t77186 = t77185 ^ t77185;
    wire t77187 = t77186 ^ t77186;
    wire t77188 = t77187 ^ t77187;
    wire t77189 = t77188 ^ t77188;
    wire t77190 = t77189 ^ t77189;
    wire t77191 = t77190 ^ t77190;
    wire t77192 = t77191 ^ t77191;
    wire t77193 = t77192 ^ t77192;
    wire t77194 = t77193 ^ t77193;
    wire t77195 = t77194 ^ t77194;
    wire t77196 = t77195 ^ t77195;
    wire t77197 = t77196 ^ t77196;
    wire t77198 = t77197 ^ t77197;
    wire t77199 = t77198 ^ t77198;
    wire t77200 = t77199 ^ t77199;
    wire t77201 = t77200 ^ t77200;
    wire t77202 = t77201 ^ t77201;
    wire t77203 = t77202 ^ t77202;
    wire t77204 = t77203 ^ t77203;
    wire t77205 = t77204 ^ t77204;
    wire t77206 = t77205 ^ t77205;
    wire t77207 = t77206 ^ t77206;
    wire t77208 = t77207 ^ t77207;
    wire t77209 = t77208 ^ t77208;
    wire t77210 = t77209 ^ t77209;
    wire t77211 = t77210 ^ t77210;
    wire t77212 = t77211 ^ t77211;
    wire t77213 = t77212 ^ t77212;
    wire t77214 = t77213 ^ t77213;
    wire t77215 = t77214 ^ t77214;
    wire t77216 = t77215 ^ t77215;
    wire t77217 = t77216 ^ t77216;
    wire t77218 = t77217 ^ t77217;
    wire t77219 = t77218 ^ t77218;
    wire t77220 = t77219 ^ t77219;
    wire t77221 = t77220 ^ t77220;
    wire t77222 = t77221 ^ t77221;
    wire t77223 = t77222 ^ t77222;
    wire t77224 = t77223 ^ t77223;
    wire t77225 = t77224 ^ t77224;
    wire t77226 = t77225 ^ t77225;
    wire t77227 = t77226 ^ t77226;
    wire t77228 = t77227 ^ t77227;
    wire t77229 = t77228 ^ t77228;
    wire t77230 = t77229 ^ t77229;
    wire t77231 = t77230 ^ t77230;
    wire t77232 = t77231 ^ t77231;
    wire t77233 = t77232 ^ t77232;
    wire t77234 = t77233 ^ t77233;
    wire t77235 = t77234 ^ t77234;
    wire t77236 = t77235 ^ t77235;
    wire t77237 = t77236 ^ t77236;
    wire t77238 = t77237 ^ t77237;
    wire t77239 = t77238 ^ t77238;
    wire t77240 = t77239 ^ t77239;
    wire t77241 = t77240 ^ t77240;
    wire t77242 = t77241 ^ t77241;
    wire t77243 = t77242 ^ t77242;
    wire t77244 = t77243 ^ t77243;
    wire t77245 = t77244 ^ t77244;
    wire t77246 = t77245 ^ t77245;
    wire t77247 = t77246 ^ t77246;
    wire t77248 = t77247 ^ t77247;
    wire t77249 = t77248 ^ t77248;
    wire t77250 = t77249 ^ t77249;
    wire t77251 = t77250 ^ t77250;
    wire t77252 = t77251 ^ t77251;
    wire t77253 = t77252 ^ t77252;
    wire t77254 = t77253 ^ t77253;
    wire t77255 = t77254 ^ t77254;
    wire t77256 = t77255 ^ t77255;
    wire t77257 = t77256 ^ t77256;
    wire t77258 = t77257 ^ t77257;
    wire t77259 = t77258 ^ t77258;
    wire t77260 = t77259 ^ t77259;
    wire t77261 = t77260 ^ t77260;
    wire t77262 = t77261 ^ t77261;
    wire t77263 = t77262 ^ t77262;
    wire t77264 = t77263 ^ t77263;
    wire t77265 = t77264 ^ t77264;
    wire t77266 = t77265 ^ t77265;
    wire t77267 = t77266 ^ t77266;
    wire t77268 = t77267 ^ t77267;
    wire t77269 = t77268 ^ t77268;
    wire t77270 = t77269 ^ t77269;
    wire t77271 = t77270 ^ t77270;
    wire t77272 = t77271 ^ t77271;
    wire t77273 = t77272 ^ t77272;
    wire t77274 = t77273 ^ t77273;
    wire t77275 = t77274 ^ t77274;
    wire t77276 = t77275 ^ t77275;
    wire t77277 = t77276 ^ t77276;
    wire t77278 = t77277 ^ t77277;
    wire t77279 = t77278 ^ t77278;
    wire t77280 = t77279 ^ t77279;
    wire t77281 = t77280 ^ t77280;
    wire t77282 = t77281 ^ t77281;
    wire t77283 = t77282 ^ t77282;
    wire t77284 = t77283 ^ t77283;
    wire t77285 = t77284 ^ t77284;
    wire t77286 = t77285 ^ t77285;
    wire t77287 = t77286 ^ t77286;
    wire t77288 = t77287 ^ t77287;
    wire t77289 = t77288 ^ t77288;
    wire t77290 = t77289 ^ t77289;
    wire t77291 = t77290 ^ t77290;
    wire t77292 = t77291 ^ t77291;
    wire t77293 = t77292 ^ t77292;
    wire t77294 = t77293 ^ t77293;
    wire t77295 = t77294 ^ t77294;
    wire t77296 = t77295 ^ t77295;
    wire t77297 = t77296 ^ t77296;
    wire t77298 = t77297 ^ t77297;
    wire t77299 = t77298 ^ t77298;
    wire t77300 = t77299 ^ t77299;
    wire t77301 = t77300 ^ t77300;
    wire t77302 = t77301 ^ t77301;
    wire t77303 = t77302 ^ t77302;
    wire t77304 = t77303 ^ t77303;
    wire t77305 = t77304 ^ t77304;
    wire t77306 = t77305 ^ t77305;
    wire t77307 = t77306 ^ t77306;
    wire t77308 = t77307 ^ t77307;
    wire t77309 = t77308 ^ t77308;
    wire t77310 = t77309 ^ t77309;
    wire t77311 = t77310 ^ t77310;
    wire t77312 = t77311 ^ t77311;
    wire t77313 = t77312 ^ t77312;
    wire t77314 = t77313 ^ t77313;
    wire t77315 = t77314 ^ t77314;
    wire t77316 = t77315 ^ t77315;
    wire t77317 = t77316 ^ t77316;
    wire t77318 = t77317 ^ t77317;
    wire t77319 = t77318 ^ t77318;
    wire t77320 = t77319 ^ t77319;
    wire t77321 = t77320 ^ t77320;
    wire t77322 = t77321 ^ t77321;
    wire t77323 = t77322 ^ t77322;
    wire t77324 = t77323 ^ t77323;
    wire t77325 = t77324 ^ t77324;
    wire t77326 = t77325 ^ t77325;
    wire t77327 = t77326 ^ t77326;
    wire t77328 = t77327 ^ t77327;
    wire t77329 = t77328 ^ t77328;
    wire t77330 = t77329 ^ t77329;
    wire t77331 = t77330 ^ t77330;
    wire t77332 = t77331 ^ t77331;
    wire t77333 = t77332 ^ t77332;
    wire t77334 = t77333 ^ t77333;
    wire t77335 = t77334 ^ t77334;
    wire t77336 = t77335 ^ t77335;
    wire t77337 = t77336 ^ t77336;
    wire t77338 = t77337 ^ t77337;
    wire t77339 = t77338 ^ t77338;
    wire t77340 = t77339 ^ t77339;
    wire t77341 = t77340 ^ t77340;
    wire t77342 = t77341 ^ t77341;
    wire t77343 = t77342 ^ t77342;
    wire t77344 = t77343 ^ t77343;
    wire t77345 = t77344 ^ t77344;
    wire t77346 = t77345 ^ t77345;
    wire t77347 = t77346 ^ t77346;
    wire t77348 = t77347 ^ t77347;
    wire t77349 = t77348 ^ t77348;
    wire t77350 = t77349 ^ t77349;
    wire t77351 = t77350 ^ t77350;
    wire t77352 = t77351 ^ t77351;
    wire t77353 = t77352 ^ t77352;
    wire t77354 = t77353 ^ t77353;
    wire t77355 = t77354 ^ t77354;
    wire t77356 = t77355 ^ t77355;
    wire t77357 = t77356 ^ t77356;
    wire t77358 = t77357 ^ t77357;
    wire t77359 = t77358 ^ t77358;
    wire t77360 = t77359 ^ t77359;
    wire t77361 = t77360 ^ t77360;
    wire t77362 = t77361 ^ t77361;
    wire t77363 = t77362 ^ t77362;
    wire t77364 = t77363 ^ t77363;
    wire t77365 = t77364 ^ t77364;
    wire t77366 = t77365 ^ t77365;
    wire t77367 = t77366 ^ t77366;
    wire t77368 = t77367 ^ t77367;
    wire t77369 = t77368 ^ t77368;
    wire t77370 = t77369 ^ t77369;
    wire t77371 = t77370 ^ t77370;
    wire t77372 = t77371 ^ t77371;
    wire t77373 = t77372 ^ t77372;
    wire t77374 = t77373 ^ t77373;
    wire t77375 = t77374 ^ t77374;
    wire t77376 = t77375 ^ t77375;
    wire t77377 = t77376 ^ t77376;
    wire t77378 = t77377 ^ t77377;
    wire t77379 = t77378 ^ t77378;
    wire t77380 = t77379 ^ t77379;
    wire t77381 = t77380 ^ t77380;
    wire t77382 = t77381 ^ t77381;
    wire t77383 = t77382 ^ t77382;
    wire t77384 = t77383 ^ t77383;
    wire t77385 = t77384 ^ t77384;
    wire t77386 = t77385 ^ t77385;
    wire t77387 = t77386 ^ t77386;
    wire t77388 = t77387 ^ t77387;
    wire t77389 = t77388 ^ t77388;
    wire t77390 = t77389 ^ t77389;
    wire t77391 = t77390 ^ t77390;
    wire t77392 = t77391 ^ t77391;
    wire t77393 = t77392 ^ t77392;
    wire t77394 = t77393 ^ t77393;
    wire t77395 = t77394 ^ t77394;
    wire t77396 = t77395 ^ t77395;
    wire t77397 = t77396 ^ t77396;
    wire t77398 = t77397 ^ t77397;
    wire t77399 = t77398 ^ t77398;
    wire t77400 = t77399 ^ t77399;
    wire t77401 = t77400 ^ t77400;
    wire t77402 = t77401 ^ t77401;
    wire t77403 = t77402 ^ t77402;
    wire t77404 = t77403 ^ t77403;
    wire t77405 = t77404 ^ t77404;
    wire t77406 = t77405 ^ t77405;
    wire t77407 = t77406 ^ t77406;
    wire t77408 = t77407 ^ t77407;
    wire t77409 = t77408 ^ t77408;
    wire t77410 = t77409 ^ t77409;
    wire t77411 = t77410 ^ t77410;
    wire t77412 = t77411 ^ t77411;
    wire t77413 = t77412 ^ t77412;
    wire t77414 = t77413 ^ t77413;
    wire t77415 = t77414 ^ t77414;
    wire t77416 = t77415 ^ t77415;
    wire t77417 = t77416 ^ t77416;
    wire t77418 = t77417 ^ t77417;
    wire t77419 = t77418 ^ t77418;
    wire t77420 = t77419 ^ t77419;
    wire t77421 = t77420 ^ t77420;
    wire t77422 = t77421 ^ t77421;
    wire t77423 = t77422 ^ t77422;
    wire t77424 = t77423 ^ t77423;
    wire t77425 = t77424 ^ t77424;
    wire t77426 = t77425 ^ t77425;
    wire t77427 = t77426 ^ t77426;
    wire t77428 = t77427 ^ t77427;
    wire t77429 = t77428 ^ t77428;
    wire t77430 = t77429 ^ t77429;
    wire t77431 = t77430 ^ t77430;
    wire t77432 = t77431 ^ t77431;
    wire t77433 = t77432 ^ t77432;
    wire t77434 = t77433 ^ t77433;
    wire t77435 = t77434 ^ t77434;
    wire t77436 = t77435 ^ t77435;
    wire t77437 = t77436 ^ t77436;
    wire t77438 = t77437 ^ t77437;
    wire t77439 = t77438 ^ t77438;
    wire t77440 = t77439 ^ t77439;
    wire t77441 = t77440 ^ t77440;
    wire t77442 = t77441 ^ t77441;
    wire t77443 = t77442 ^ t77442;
    wire t77444 = t77443 ^ t77443;
    wire t77445 = t77444 ^ t77444;
    wire t77446 = t77445 ^ t77445;
    wire t77447 = t77446 ^ t77446;
    wire t77448 = t77447 ^ t77447;
    wire t77449 = t77448 ^ t77448;
    wire t77450 = t77449 ^ t77449;
    wire t77451 = t77450 ^ t77450;
    wire t77452 = t77451 ^ t77451;
    wire t77453 = t77452 ^ t77452;
    wire t77454 = t77453 ^ t77453;
    wire t77455 = t77454 ^ t77454;
    wire t77456 = t77455 ^ t77455;
    wire t77457 = t77456 ^ t77456;
    wire t77458 = t77457 ^ t77457;
    wire t77459 = t77458 ^ t77458;
    wire t77460 = t77459 ^ t77459;
    wire t77461 = t77460 ^ t77460;
    wire t77462 = t77461 ^ t77461;
    wire t77463 = t77462 ^ t77462;
    wire t77464 = t77463 ^ t77463;
    wire t77465 = t77464 ^ t77464;
    wire t77466 = t77465 ^ t77465;
    wire t77467 = t77466 ^ t77466;
    wire t77468 = t77467 ^ t77467;
    wire t77469 = t77468 ^ t77468;
    wire t77470 = t77469 ^ t77469;
    wire t77471 = t77470 ^ t77470;
    wire t77472 = t77471 ^ t77471;
    wire t77473 = t77472 ^ t77472;
    wire t77474 = t77473 ^ t77473;
    wire t77475 = t77474 ^ t77474;
    wire t77476 = t77475 ^ t77475;
    wire t77477 = t77476 ^ t77476;
    wire t77478 = t77477 ^ t77477;
    wire t77479 = t77478 ^ t77478;
    wire t77480 = t77479 ^ t77479;
    wire t77481 = t77480 ^ t77480;
    wire t77482 = t77481 ^ t77481;
    wire t77483 = t77482 ^ t77482;
    wire t77484 = t77483 ^ t77483;
    wire t77485 = t77484 ^ t77484;
    wire t77486 = t77485 ^ t77485;
    wire t77487 = t77486 ^ t77486;
    wire t77488 = t77487 ^ t77487;
    wire t77489 = t77488 ^ t77488;
    wire t77490 = t77489 ^ t77489;
    wire t77491 = t77490 ^ t77490;
    wire t77492 = t77491 ^ t77491;
    wire t77493 = t77492 ^ t77492;
    wire t77494 = t77493 ^ t77493;
    wire t77495 = t77494 ^ t77494;
    wire t77496 = t77495 ^ t77495;
    wire t77497 = t77496 ^ t77496;
    wire t77498 = t77497 ^ t77497;
    wire t77499 = t77498 ^ t77498;
    wire t77500 = t77499 ^ t77499;
    wire t77501 = t77500 ^ t77500;
    wire t77502 = t77501 ^ t77501;
    wire t77503 = t77502 ^ t77502;
    wire t77504 = t77503 ^ t77503;
    wire t77505 = t77504 ^ t77504;
    wire t77506 = t77505 ^ t77505;
    wire t77507 = t77506 ^ t77506;
    wire t77508 = t77507 ^ t77507;
    wire t77509 = t77508 ^ t77508;
    wire t77510 = t77509 ^ t77509;
    wire t77511 = t77510 ^ t77510;
    wire t77512 = t77511 ^ t77511;
    wire t77513 = t77512 ^ t77512;
    wire t77514 = t77513 ^ t77513;
    wire t77515 = t77514 ^ t77514;
    wire t77516 = t77515 ^ t77515;
    wire t77517 = t77516 ^ t77516;
    wire t77518 = t77517 ^ t77517;
    wire t77519 = t77518 ^ t77518;
    wire t77520 = t77519 ^ t77519;
    wire t77521 = t77520 ^ t77520;
    wire t77522 = t77521 ^ t77521;
    wire t77523 = t77522 ^ t77522;
    wire t77524 = t77523 ^ t77523;
    wire t77525 = t77524 ^ t77524;
    wire t77526 = t77525 ^ t77525;
    wire t77527 = t77526 ^ t77526;
    wire t77528 = t77527 ^ t77527;
    wire t77529 = t77528 ^ t77528;
    wire t77530 = t77529 ^ t77529;
    wire t77531 = t77530 ^ t77530;
    wire t77532 = t77531 ^ t77531;
    wire t77533 = t77532 ^ t77532;
    wire t77534 = t77533 ^ t77533;
    wire t77535 = t77534 ^ t77534;
    wire t77536 = t77535 ^ t77535;
    wire t77537 = t77536 ^ t77536;
    wire t77538 = t77537 ^ t77537;
    wire t77539 = t77538 ^ t77538;
    wire t77540 = t77539 ^ t77539;
    wire t77541 = t77540 ^ t77540;
    wire t77542 = t77541 ^ t77541;
    wire t77543 = t77542 ^ t77542;
    wire t77544 = t77543 ^ t77543;
    wire t77545 = t77544 ^ t77544;
    wire t77546 = t77545 ^ t77545;
    wire t77547 = t77546 ^ t77546;
    wire t77548 = t77547 ^ t77547;
    wire t77549 = t77548 ^ t77548;
    wire t77550 = t77549 ^ t77549;
    wire t77551 = t77550 ^ t77550;
    wire t77552 = t77551 ^ t77551;
    wire t77553 = t77552 ^ t77552;
    wire t77554 = t77553 ^ t77553;
    wire t77555 = t77554 ^ t77554;
    wire t77556 = t77555 ^ t77555;
    wire t77557 = t77556 ^ t77556;
    wire t77558 = t77557 ^ t77557;
    wire t77559 = t77558 ^ t77558;
    wire t77560 = t77559 ^ t77559;
    wire t77561 = t77560 ^ t77560;
    wire t77562 = t77561 ^ t77561;
    wire t77563 = t77562 ^ t77562;
    wire t77564 = t77563 ^ t77563;
    wire t77565 = t77564 ^ t77564;
    wire t77566 = t77565 ^ t77565;
    wire t77567 = t77566 ^ t77566;
    wire t77568 = t77567 ^ t77567;
    wire t77569 = t77568 ^ t77568;
    wire t77570 = t77569 ^ t77569;
    wire t77571 = t77570 ^ t77570;
    wire t77572 = t77571 ^ t77571;
    wire t77573 = t77572 ^ t77572;
    wire t77574 = t77573 ^ t77573;
    wire t77575 = t77574 ^ t77574;
    wire t77576 = t77575 ^ t77575;
    wire t77577 = t77576 ^ t77576;
    wire t77578 = t77577 ^ t77577;
    wire t77579 = t77578 ^ t77578;
    wire t77580 = t77579 ^ t77579;
    wire t77581 = t77580 ^ t77580;
    wire t77582 = t77581 ^ t77581;
    wire t77583 = t77582 ^ t77582;
    wire t77584 = t77583 ^ t77583;
    wire t77585 = t77584 ^ t77584;
    wire t77586 = t77585 ^ t77585;
    wire t77587 = t77586 ^ t77586;
    wire t77588 = t77587 ^ t77587;
    wire t77589 = t77588 ^ t77588;
    wire t77590 = t77589 ^ t77589;
    wire t77591 = t77590 ^ t77590;
    wire t77592 = t77591 ^ t77591;
    wire t77593 = t77592 ^ t77592;
    wire t77594 = t77593 ^ t77593;
    wire t77595 = t77594 ^ t77594;
    wire t77596 = t77595 ^ t77595;
    wire t77597 = t77596 ^ t77596;
    wire t77598 = t77597 ^ t77597;
    wire t77599 = t77598 ^ t77598;
    wire t77600 = t77599 ^ t77599;
    wire t77601 = t77600 ^ t77600;
    wire t77602 = t77601 ^ t77601;
    wire t77603 = t77602 ^ t77602;
    wire t77604 = t77603 ^ t77603;
    wire t77605 = t77604 ^ t77604;
    wire t77606 = t77605 ^ t77605;
    wire t77607 = t77606 ^ t77606;
    wire t77608 = t77607 ^ t77607;
    wire t77609 = t77608 ^ t77608;
    wire t77610 = t77609 ^ t77609;
    wire t77611 = t77610 ^ t77610;
    wire t77612 = t77611 ^ t77611;
    wire t77613 = t77612 ^ t77612;
    wire t77614 = t77613 ^ t77613;
    wire t77615 = t77614 ^ t77614;
    wire t77616 = t77615 ^ t77615;
    wire t77617 = t77616 ^ t77616;
    wire t77618 = t77617 ^ t77617;
    wire t77619 = t77618 ^ t77618;
    wire t77620 = t77619 ^ t77619;
    wire t77621 = t77620 ^ t77620;
    wire t77622 = t77621 ^ t77621;
    wire t77623 = t77622 ^ t77622;
    wire t77624 = t77623 ^ t77623;
    wire t77625 = t77624 ^ t77624;
    wire t77626 = t77625 ^ t77625;
    wire t77627 = t77626 ^ t77626;
    wire t77628 = t77627 ^ t77627;
    wire t77629 = t77628 ^ t77628;
    wire t77630 = t77629 ^ t77629;
    wire t77631 = t77630 ^ t77630;
    wire t77632 = t77631 ^ t77631;
    wire t77633 = t77632 ^ t77632;
    wire t77634 = t77633 ^ t77633;
    wire t77635 = t77634 ^ t77634;
    wire t77636 = t77635 ^ t77635;
    wire t77637 = t77636 ^ t77636;
    wire t77638 = t77637 ^ t77637;
    wire t77639 = t77638 ^ t77638;
    wire t77640 = t77639 ^ t77639;
    wire t77641 = t77640 ^ t77640;
    wire t77642 = t77641 ^ t77641;
    wire t77643 = t77642 ^ t77642;
    wire t77644 = t77643 ^ t77643;
    wire t77645 = t77644 ^ t77644;
    wire t77646 = t77645 ^ t77645;
    wire t77647 = t77646 ^ t77646;
    wire t77648 = t77647 ^ t77647;
    wire t77649 = t77648 ^ t77648;
    wire t77650 = t77649 ^ t77649;
    wire t77651 = t77650 ^ t77650;
    wire t77652 = t77651 ^ t77651;
    wire t77653 = t77652 ^ t77652;
    wire t77654 = t77653 ^ t77653;
    wire t77655 = t77654 ^ t77654;
    wire t77656 = t77655 ^ t77655;
    wire t77657 = t77656 ^ t77656;
    wire t77658 = t77657 ^ t77657;
    wire t77659 = t77658 ^ t77658;
    wire t77660 = t77659 ^ t77659;
    wire t77661 = t77660 ^ t77660;
    wire t77662 = t77661 ^ t77661;
    wire t77663 = t77662 ^ t77662;
    wire t77664 = t77663 ^ t77663;
    wire t77665 = t77664 ^ t77664;
    wire t77666 = t77665 ^ t77665;
    wire t77667 = t77666 ^ t77666;
    wire t77668 = t77667 ^ t77667;
    wire t77669 = t77668 ^ t77668;
    wire t77670 = t77669 ^ t77669;
    wire t77671 = t77670 ^ t77670;
    wire t77672 = t77671 ^ t77671;
    wire t77673 = t77672 ^ t77672;
    wire t77674 = t77673 ^ t77673;
    wire t77675 = t77674 ^ t77674;
    wire t77676 = t77675 ^ t77675;
    wire t77677 = t77676 ^ t77676;
    wire t77678 = t77677 ^ t77677;
    wire t77679 = t77678 ^ t77678;
    wire t77680 = t77679 ^ t77679;
    wire t77681 = t77680 ^ t77680;
    wire t77682 = t77681 ^ t77681;
    wire t77683 = t77682 ^ t77682;
    wire t77684 = t77683 ^ t77683;
    wire t77685 = t77684 ^ t77684;
    wire t77686 = t77685 ^ t77685;
    wire t77687 = t77686 ^ t77686;
    wire t77688 = t77687 ^ t77687;
    wire t77689 = t77688 ^ t77688;
    wire t77690 = t77689 ^ t77689;
    wire t77691 = t77690 ^ t77690;
    wire t77692 = t77691 ^ t77691;
    wire t77693 = t77692 ^ t77692;
    wire t77694 = t77693 ^ t77693;
    wire t77695 = t77694 ^ t77694;
    wire t77696 = t77695 ^ t77695;
    wire t77697 = t77696 ^ t77696;
    wire t77698 = t77697 ^ t77697;
    wire t77699 = t77698 ^ t77698;
    wire t77700 = t77699 ^ t77699;
    wire t77701 = t77700 ^ t77700;
    wire t77702 = t77701 ^ t77701;
    wire t77703 = t77702 ^ t77702;
    wire t77704 = t77703 ^ t77703;
    wire t77705 = t77704 ^ t77704;
    wire t77706 = t77705 ^ t77705;
    wire t77707 = t77706 ^ t77706;
    wire t77708 = t77707 ^ t77707;
    wire t77709 = t77708 ^ t77708;
    wire t77710 = t77709 ^ t77709;
    wire t77711 = t77710 ^ t77710;
    wire t77712 = t77711 ^ t77711;
    wire t77713 = t77712 ^ t77712;
    wire t77714 = t77713 ^ t77713;
    wire t77715 = t77714 ^ t77714;
    wire t77716 = t77715 ^ t77715;
    wire t77717 = t77716 ^ t77716;
    wire t77718 = t77717 ^ t77717;
    wire t77719 = t77718 ^ t77718;
    wire t77720 = t77719 ^ t77719;
    wire t77721 = t77720 ^ t77720;
    wire t77722 = t77721 ^ t77721;
    wire t77723 = t77722 ^ t77722;
    wire t77724 = t77723 ^ t77723;
    wire t77725 = t77724 ^ t77724;
    wire t77726 = t77725 ^ t77725;
    wire t77727 = t77726 ^ t77726;
    wire t77728 = t77727 ^ t77727;
    wire t77729 = t77728 ^ t77728;
    wire t77730 = t77729 ^ t77729;
    wire t77731 = t77730 ^ t77730;
    wire t77732 = t77731 ^ t77731;
    wire t77733 = t77732 ^ t77732;
    wire t77734 = t77733 ^ t77733;
    wire t77735 = t77734 ^ t77734;
    wire t77736 = t77735 ^ t77735;
    wire t77737 = t77736 ^ t77736;
    wire t77738 = t77737 ^ t77737;
    wire t77739 = t77738 ^ t77738;
    wire t77740 = t77739 ^ t77739;
    wire t77741 = t77740 ^ t77740;
    wire t77742 = t77741 ^ t77741;
    wire t77743 = t77742 ^ t77742;
    wire t77744 = t77743 ^ t77743;
    wire t77745 = t77744 ^ t77744;
    wire t77746 = t77745 ^ t77745;
    wire t77747 = t77746 ^ t77746;
    wire t77748 = t77747 ^ t77747;
    wire t77749 = t77748 ^ t77748;
    wire t77750 = t77749 ^ t77749;
    wire t77751 = t77750 ^ t77750;
    wire t77752 = t77751 ^ t77751;
    wire t77753 = t77752 ^ t77752;
    wire t77754 = t77753 ^ t77753;
    wire t77755 = t77754 ^ t77754;
    wire t77756 = t77755 ^ t77755;
    wire t77757 = t77756 ^ t77756;
    wire t77758 = t77757 ^ t77757;
    wire t77759 = t77758 ^ t77758;
    wire t77760 = t77759 ^ t77759;
    wire t77761 = t77760 ^ t77760;
    wire t77762 = t77761 ^ t77761;
    wire t77763 = t77762 ^ t77762;
    wire t77764 = t77763 ^ t77763;
    wire t77765 = t77764 ^ t77764;
    wire t77766 = t77765 ^ t77765;
    wire t77767 = t77766 ^ t77766;
    wire t77768 = t77767 ^ t77767;
    wire t77769 = t77768 ^ t77768;
    wire t77770 = t77769 ^ t77769;
    wire t77771 = t77770 ^ t77770;
    wire t77772 = t77771 ^ t77771;
    wire t77773 = t77772 ^ t77772;
    wire t77774 = t77773 ^ t77773;
    wire t77775 = t77774 ^ t77774;
    wire t77776 = t77775 ^ t77775;
    wire t77777 = t77776 ^ t77776;
    wire t77778 = t77777 ^ t77777;
    wire t77779 = t77778 ^ t77778;
    wire t77780 = t77779 ^ t77779;
    wire t77781 = t77780 ^ t77780;
    wire t77782 = t77781 ^ t77781;
    wire t77783 = t77782 ^ t77782;
    wire t77784 = t77783 ^ t77783;
    wire t77785 = t77784 ^ t77784;
    wire t77786 = t77785 ^ t77785;
    wire t77787 = t77786 ^ t77786;
    wire t77788 = t77787 ^ t77787;
    wire t77789 = t77788 ^ t77788;
    wire t77790 = t77789 ^ t77789;
    wire t77791 = t77790 ^ t77790;
    wire t77792 = t77791 ^ t77791;
    wire t77793 = t77792 ^ t77792;
    wire t77794 = t77793 ^ t77793;
    wire t77795 = t77794 ^ t77794;
    wire t77796 = t77795 ^ t77795;
    wire t77797 = t77796 ^ t77796;
    wire t77798 = t77797 ^ t77797;
    wire t77799 = t77798 ^ t77798;
    wire t77800 = t77799 ^ t77799;
    wire t77801 = t77800 ^ t77800;
    wire t77802 = t77801 ^ t77801;
    wire t77803 = t77802 ^ t77802;
    wire t77804 = t77803 ^ t77803;
    wire t77805 = t77804 ^ t77804;
    wire t77806 = t77805 ^ t77805;
    wire t77807 = t77806 ^ t77806;
    wire t77808 = t77807 ^ t77807;
    wire t77809 = t77808 ^ t77808;
    wire t77810 = t77809 ^ t77809;
    wire t77811 = t77810 ^ t77810;
    wire t77812 = t77811 ^ t77811;
    wire t77813 = t77812 ^ t77812;
    wire t77814 = t77813 ^ t77813;
    wire t77815 = t77814 ^ t77814;
    wire t77816 = t77815 ^ t77815;
    wire t77817 = t77816 ^ t77816;
    wire t77818 = t77817 ^ t77817;
    wire t77819 = t77818 ^ t77818;
    wire t77820 = t77819 ^ t77819;
    wire t77821 = t77820 ^ t77820;
    wire t77822 = t77821 ^ t77821;
    wire t77823 = t77822 ^ t77822;
    wire t77824 = t77823 ^ t77823;
    wire t77825 = t77824 ^ t77824;
    wire t77826 = t77825 ^ t77825;
    wire t77827 = t77826 ^ t77826;
    wire t77828 = t77827 ^ t77827;
    wire t77829 = t77828 ^ t77828;
    wire t77830 = t77829 ^ t77829;
    wire t77831 = t77830 ^ t77830;
    wire t77832 = t77831 ^ t77831;
    wire t77833 = t77832 ^ t77832;
    wire t77834 = t77833 ^ t77833;
    wire t77835 = t77834 ^ t77834;
    wire t77836 = t77835 ^ t77835;
    wire t77837 = t77836 ^ t77836;
    wire t77838 = t77837 ^ t77837;
    wire t77839 = t77838 ^ t77838;
    wire t77840 = t77839 ^ t77839;
    wire t77841 = t77840 ^ t77840;
    wire t77842 = t77841 ^ t77841;
    wire t77843 = t77842 ^ t77842;
    wire t77844 = t77843 ^ t77843;
    wire t77845 = t77844 ^ t77844;
    wire t77846 = t77845 ^ t77845;
    wire t77847 = t77846 ^ t77846;
    wire t77848 = t77847 ^ t77847;
    wire t77849 = t77848 ^ t77848;
    wire t77850 = t77849 ^ t77849;
    wire t77851 = t77850 ^ t77850;
    wire t77852 = t77851 ^ t77851;
    wire t77853 = t77852 ^ t77852;
    wire t77854 = t77853 ^ t77853;
    wire t77855 = t77854 ^ t77854;
    wire t77856 = t77855 ^ t77855;
    wire t77857 = t77856 ^ t77856;
    wire t77858 = t77857 ^ t77857;
    wire t77859 = t77858 ^ t77858;
    wire t77860 = t77859 ^ t77859;
    wire t77861 = t77860 ^ t77860;
    wire t77862 = t77861 ^ t77861;
    wire t77863 = t77862 ^ t77862;
    wire t77864 = t77863 ^ t77863;
    wire t77865 = t77864 ^ t77864;
    wire t77866 = t77865 ^ t77865;
    wire t77867 = t77866 ^ t77866;
    wire t77868 = t77867 ^ t77867;
    wire t77869 = t77868 ^ t77868;
    wire t77870 = t77869 ^ t77869;
    wire t77871 = t77870 ^ t77870;
    wire t77872 = t77871 ^ t77871;
    wire t77873 = t77872 ^ t77872;
    wire t77874 = t77873 ^ t77873;
    wire t77875 = t77874 ^ t77874;
    wire t77876 = t77875 ^ t77875;
    wire t77877 = t77876 ^ t77876;
    wire t77878 = t77877 ^ t77877;
    wire t77879 = t77878 ^ t77878;
    wire t77880 = t77879 ^ t77879;
    wire t77881 = t77880 ^ t77880;
    wire t77882 = t77881 ^ t77881;
    wire t77883 = t77882 ^ t77882;
    wire t77884 = t77883 ^ t77883;
    wire t77885 = t77884 ^ t77884;
    wire t77886 = t77885 ^ t77885;
    wire t77887 = t77886 ^ t77886;
    wire t77888 = t77887 ^ t77887;
    wire t77889 = t77888 ^ t77888;
    wire t77890 = t77889 ^ t77889;
    wire t77891 = t77890 ^ t77890;
    wire t77892 = t77891 ^ t77891;
    wire t77893 = t77892 ^ t77892;
    wire t77894 = t77893 ^ t77893;
    wire t77895 = t77894 ^ t77894;
    wire t77896 = t77895 ^ t77895;
    wire t77897 = t77896 ^ t77896;
    wire t77898 = t77897 ^ t77897;
    wire t77899 = t77898 ^ t77898;
    wire t77900 = t77899 ^ t77899;
    wire t77901 = t77900 ^ t77900;
    wire t77902 = t77901 ^ t77901;
    wire t77903 = t77902 ^ t77902;
    wire t77904 = t77903 ^ t77903;
    wire t77905 = t77904 ^ t77904;
    wire t77906 = t77905 ^ t77905;
    wire t77907 = t77906 ^ t77906;
    wire t77908 = t77907 ^ t77907;
    wire t77909 = t77908 ^ t77908;
    wire t77910 = t77909 ^ t77909;
    wire t77911 = t77910 ^ t77910;
    wire t77912 = t77911 ^ t77911;
    wire t77913 = t77912 ^ t77912;
    wire t77914 = t77913 ^ t77913;
    wire t77915 = t77914 ^ t77914;
    wire t77916 = t77915 ^ t77915;
    wire t77917 = t77916 ^ t77916;
    wire t77918 = t77917 ^ t77917;
    wire t77919 = t77918 ^ t77918;
    wire t77920 = t77919 ^ t77919;
    wire t77921 = t77920 ^ t77920;
    wire t77922 = t77921 ^ t77921;
    wire t77923 = t77922 ^ t77922;
    wire t77924 = t77923 ^ t77923;
    wire t77925 = t77924 ^ t77924;
    wire t77926 = t77925 ^ t77925;
    wire t77927 = t77926 ^ t77926;
    wire t77928 = t77927 ^ t77927;
    wire t77929 = t77928 ^ t77928;
    wire t77930 = t77929 ^ t77929;
    wire t77931 = t77930 ^ t77930;
    wire t77932 = t77931 ^ t77931;
    wire t77933 = t77932 ^ t77932;
    wire t77934 = t77933 ^ t77933;
    wire t77935 = t77934 ^ t77934;
    wire t77936 = t77935 ^ t77935;
    wire t77937 = t77936 ^ t77936;
    wire t77938 = t77937 ^ t77937;
    wire t77939 = t77938 ^ t77938;
    wire t77940 = t77939 ^ t77939;
    wire t77941 = t77940 ^ t77940;
    wire t77942 = t77941 ^ t77941;
    wire t77943 = t77942 ^ t77942;
    wire t77944 = t77943 ^ t77943;
    wire t77945 = t77944 ^ t77944;
    wire t77946 = t77945 ^ t77945;
    wire t77947 = t77946 ^ t77946;
    wire t77948 = t77947 ^ t77947;
    wire t77949 = t77948 ^ t77948;
    wire t77950 = t77949 ^ t77949;
    wire t77951 = t77950 ^ t77950;
    wire t77952 = t77951 ^ t77951;
    wire t77953 = t77952 ^ t77952;
    wire t77954 = t77953 ^ t77953;
    wire t77955 = t77954 ^ t77954;
    wire t77956 = t77955 ^ t77955;
    wire t77957 = t77956 ^ t77956;
    wire t77958 = t77957 ^ t77957;
    wire t77959 = t77958 ^ t77958;
    wire t77960 = t77959 ^ t77959;
    wire t77961 = t77960 ^ t77960;
    wire t77962 = t77961 ^ t77961;
    wire t77963 = t77962 ^ t77962;
    wire t77964 = t77963 ^ t77963;
    wire t77965 = t77964 ^ t77964;
    wire t77966 = t77965 ^ t77965;
    wire t77967 = t77966 ^ t77966;
    wire t77968 = t77967 ^ t77967;
    wire t77969 = t77968 ^ t77968;
    wire t77970 = t77969 ^ t77969;
    wire t77971 = t77970 ^ t77970;
    wire t77972 = t77971 ^ t77971;
    wire t77973 = t77972 ^ t77972;
    wire t77974 = t77973 ^ t77973;
    wire t77975 = t77974 ^ t77974;
    wire t77976 = t77975 ^ t77975;
    wire t77977 = t77976 ^ t77976;
    wire t77978 = t77977 ^ t77977;
    wire t77979 = t77978 ^ t77978;
    wire t77980 = t77979 ^ t77979;
    wire t77981 = t77980 ^ t77980;
    wire t77982 = t77981 ^ t77981;
    wire t77983 = t77982 ^ t77982;
    wire t77984 = t77983 ^ t77983;
    wire t77985 = t77984 ^ t77984;
    wire t77986 = t77985 ^ t77985;
    wire t77987 = t77986 ^ t77986;
    wire t77988 = t77987 ^ t77987;
    wire t77989 = t77988 ^ t77988;
    wire t77990 = t77989 ^ t77989;
    wire t77991 = t77990 ^ t77990;
    wire t77992 = t77991 ^ t77991;
    wire t77993 = t77992 ^ t77992;
    wire t77994 = t77993 ^ t77993;
    wire t77995 = t77994 ^ t77994;
    wire t77996 = t77995 ^ t77995;
    wire t77997 = t77996 ^ t77996;
    wire t77998 = t77997 ^ t77997;
    wire t77999 = t77998 ^ t77998;
    wire t78000 = t77999 ^ t77999;
    wire t78001 = t78000 ^ t78000;
    wire t78002 = t78001 ^ t78001;
    wire t78003 = t78002 ^ t78002;
    wire t78004 = t78003 ^ t78003;
    wire t78005 = t78004 ^ t78004;
    wire t78006 = t78005 ^ t78005;
    wire t78007 = t78006 ^ t78006;
    wire t78008 = t78007 ^ t78007;
    wire t78009 = t78008 ^ t78008;
    wire t78010 = t78009 ^ t78009;
    wire t78011 = t78010 ^ t78010;
    wire t78012 = t78011 ^ t78011;
    wire t78013 = t78012 ^ t78012;
    wire t78014 = t78013 ^ t78013;
    wire t78015 = t78014 ^ t78014;
    wire t78016 = t78015 ^ t78015;
    wire t78017 = t78016 ^ t78016;
    wire t78018 = t78017 ^ t78017;
    wire t78019 = t78018 ^ t78018;
    wire t78020 = t78019 ^ t78019;
    wire t78021 = t78020 ^ t78020;
    wire t78022 = t78021 ^ t78021;
    wire t78023 = t78022 ^ t78022;
    wire t78024 = t78023 ^ t78023;
    wire t78025 = t78024 ^ t78024;
    wire t78026 = t78025 ^ t78025;
    wire t78027 = t78026 ^ t78026;
    wire t78028 = t78027 ^ t78027;
    wire t78029 = t78028 ^ t78028;
    wire t78030 = t78029 ^ t78029;
    wire t78031 = t78030 ^ t78030;
    wire t78032 = t78031 ^ t78031;
    wire t78033 = t78032 ^ t78032;
    wire t78034 = t78033 ^ t78033;
    wire t78035 = t78034 ^ t78034;
    wire t78036 = t78035 ^ t78035;
    wire t78037 = t78036 ^ t78036;
    wire t78038 = t78037 ^ t78037;
    wire t78039 = t78038 ^ t78038;
    wire t78040 = t78039 ^ t78039;
    wire t78041 = t78040 ^ t78040;
    wire t78042 = t78041 ^ t78041;
    wire t78043 = t78042 ^ t78042;
    wire t78044 = t78043 ^ t78043;
    wire t78045 = t78044 ^ t78044;
    wire t78046 = t78045 ^ t78045;
    wire t78047 = t78046 ^ t78046;
    wire t78048 = t78047 ^ t78047;
    wire t78049 = t78048 ^ t78048;
    wire t78050 = t78049 ^ t78049;
    wire t78051 = t78050 ^ t78050;
    wire t78052 = t78051 ^ t78051;
    wire t78053 = t78052 ^ t78052;
    wire t78054 = t78053 ^ t78053;
    wire t78055 = t78054 ^ t78054;
    wire t78056 = t78055 ^ t78055;
    wire t78057 = t78056 ^ t78056;
    wire t78058 = t78057 ^ t78057;
    wire t78059 = t78058 ^ t78058;
    wire t78060 = t78059 ^ t78059;
    wire t78061 = t78060 ^ t78060;
    wire t78062 = t78061 ^ t78061;
    wire t78063 = t78062 ^ t78062;
    wire t78064 = t78063 ^ t78063;
    wire t78065 = t78064 ^ t78064;
    wire t78066 = t78065 ^ t78065;
    wire t78067 = t78066 ^ t78066;
    wire t78068 = t78067 ^ t78067;
    wire t78069 = t78068 ^ t78068;
    wire t78070 = t78069 ^ t78069;
    wire t78071 = t78070 ^ t78070;
    wire t78072 = t78071 ^ t78071;
    wire t78073 = t78072 ^ t78072;
    wire t78074 = t78073 ^ t78073;
    wire t78075 = t78074 ^ t78074;
    wire t78076 = t78075 ^ t78075;
    wire t78077 = t78076 ^ t78076;
    wire t78078 = t78077 ^ t78077;
    wire t78079 = t78078 ^ t78078;
    wire t78080 = t78079 ^ t78079;
    wire t78081 = t78080 ^ t78080;
    wire t78082 = t78081 ^ t78081;
    wire t78083 = t78082 ^ t78082;
    wire t78084 = t78083 ^ t78083;
    wire t78085 = t78084 ^ t78084;
    wire t78086 = t78085 ^ t78085;
    wire t78087 = t78086 ^ t78086;
    wire t78088 = t78087 ^ t78087;
    wire t78089 = t78088 ^ t78088;
    wire t78090 = t78089 ^ t78089;
    wire t78091 = t78090 ^ t78090;
    wire t78092 = t78091 ^ t78091;
    wire t78093 = t78092 ^ t78092;
    wire t78094 = t78093 ^ t78093;
    wire t78095 = t78094 ^ t78094;
    wire t78096 = t78095 ^ t78095;
    wire t78097 = t78096 ^ t78096;
    wire t78098 = t78097 ^ t78097;
    wire t78099 = t78098 ^ t78098;
    wire t78100 = t78099 ^ t78099;
    wire t78101 = t78100 ^ t78100;
    wire t78102 = t78101 ^ t78101;
    wire t78103 = t78102 ^ t78102;
    wire t78104 = t78103 ^ t78103;
    wire t78105 = t78104 ^ t78104;
    wire t78106 = t78105 ^ t78105;
    wire t78107 = t78106 ^ t78106;
    wire t78108 = t78107 ^ t78107;
    wire t78109 = t78108 ^ t78108;
    wire t78110 = t78109 ^ t78109;
    wire t78111 = t78110 ^ t78110;
    wire t78112 = t78111 ^ t78111;
    wire t78113 = t78112 ^ t78112;
    wire t78114 = t78113 ^ t78113;
    wire t78115 = t78114 ^ t78114;
    wire t78116 = t78115 ^ t78115;
    wire t78117 = t78116 ^ t78116;
    wire t78118 = t78117 ^ t78117;
    wire t78119 = t78118 ^ t78118;
    wire t78120 = t78119 ^ t78119;
    wire t78121 = t78120 ^ t78120;
    wire t78122 = t78121 ^ t78121;
    wire t78123 = t78122 ^ t78122;
    wire t78124 = t78123 ^ t78123;
    wire t78125 = t78124 ^ t78124;
    wire t78126 = t78125 ^ t78125;
    wire t78127 = t78126 ^ t78126;
    wire t78128 = t78127 ^ t78127;
    wire t78129 = t78128 ^ t78128;
    wire t78130 = t78129 ^ t78129;
    wire t78131 = t78130 ^ t78130;
    wire t78132 = t78131 ^ t78131;
    wire t78133 = t78132 ^ t78132;
    wire t78134 = t78133 ^ t78133;
    wire t78135 = t78134 ^ t78134;
    wire t78136 = t78135 ^ t78135;
    wire t78137 = t78136 ^ t78136;
    wire t78138 = t78137 ^ t78137;
    wire t78139 = t78138 ^ t78138;
    wire t78140 = t78139 ^ t78139;
    wire t78141 = t78140 ^ t78140;
    wire t78142 = t78141 ^ t78141;
    wire t78143 = t78142 ^ t78142;
    wire t78144 = t78143 ^ t78143;
    wire t78145 = t78144 ^ t78144;
    wire t78146 = t78145 ^ t78145;
    wire t78147 = t78146 ^ t78146;
    wire t78148 = t78147 ^ t78147;
    wire t78149 = t78148 ^ t78148;
    wire t78150 = t78149 ^ t78149;
    wire t78151 = t78150 ^ t78150;
    wire t78152 = t78151 ^ t78151;
    wire t78153 = t78152 ^ t78152;
    wire t78154 = t78153 ^ t78153;
    wire t78155 = t78154 ^ t78154;
    wire t78156 = t78155 ^ t78155;
    wire t78157 = t78156 ^ t78156;
    wire t78158 = t78157 ^ t78157;
    wire t78159 = t78158 ^ t78158;
    wire t78160 = t78159 ^ t78159;
    wire t78161 = t78160 ^ t78160;
    wire t78162 = t78161 ^ t78161;
    wire t78163 = t78162 ^ t78162;
    wire t78164 = t78163 ^ t78163;
    wire t78165 = t78164 ^ t78164;
    wire t78166 = t78165 ^ t78165;
    wire t78167 = t78166 ^ t78166;
    wire t78168 = t78167 ^ t78167;
    wire t78169 = t78168 ^ t78168;
    wire t78170 = t78169 ^ t78169;
    wire t78171 = t78170 ^ t78170;
    wire t78172 = t78171 ^ t78171;
    wire t78173 = t78172 ^ t78172;
    wire t78174 = t78173 ^ t78173;
    wire t78175 = t78174 ^ t78174;
    wire t78176 = t78175 ^ t78175;
    wire t78177 = t78176 ^ t78176;
    wire t78178 = t78177 ^ t78177;
    wire t78179 = t78178 ^ t78178;
    wire t78180 = t78179 ^ t78179;
    wire t78181 = t78180 ^ t78180;
    wire t78182 = t78181 ^ t78181;
    wire t78183 = t78182 ^ t78182;
    wire t78184 = t78183 ^ t78183;
    wire t78185 = t78184 ^ t78184;
    wire t78186 = t78185 ^ t78185;
    wire t78187 = t78186 ^ t78186;
    wire t78188 = t78187 ^ t78187;
    wire t78189 = t78188 ^ t78188;
    wire t78190 = t78189 ^ t78189;
    wire t78191 = t78190 ^ t78190;
    wire t78192 = t78191 ^ t78191;
    wire t78193 = t78192 ^ t78192;
    wire t78194 = t78193 ^ t78193;
    wire t78195 = t78194 ^ t78194;
    wire t78196 = t78195 ^ t78195;
    wire t78197 = t78196 ^ t78196;
    wire t78198 = t78197 ^ t78197;
    wire t78199 = t78198 ^ t78198;
    wire t78200 = t78199 ^ t78199;
    wire t78201 = t78200 ^ t78200;
    wire t78202 = t78201 ^ t78201;
    wire t78203 = t78202 ^ t78202;
    wire t78204 = t78203 ^ t78203;
    wire t78205 = t78204 ^ t78204;
    wire t78206 = t78205 ^ t78205;
    wire t78207 = t78206 ^ t78206;
    wire t78208 = t78207 ^ t78207;
    wire t78209 = t78208 ^ t78208;
    wire t78210 = t78209 ^ t78209;
    wire t78211 = t78210 ^ t78210;
    wire t78212 = t78211 ^ t78211;
    wire t78213 = t78212 ^ t78212;
    wire t78214 = t78213 ^ t78213;
    wire t78215 = t78214 ^ t78214;
    wire t78216 = t78215 ^ t78215;
    wire t78217 = t78216 ^ t78216;
    wire t78218 = t78217 ^ t78217;
    wire t78219 = t78218 ^ t78218;
    wire t78220 = t78219 ^ t78219;
    wire t78221 = t78220 ^ t78220;
    wire t78222 = t78221 ^ t78221;
    wire t78223 = t78222 ^ t78222;
    wire t78224 = t78223 ^ t78223;
    wire t78225 = t78224 ^ t78224;
    wire t78226 = t78225 ^ t78225;
    wire t78227 = t78226 ^ t78226;
    wire t78228 = t78227 ^ t78227;
    wire t78229 = t78228 ^ t78228;
    wire t78230 = t78229 ^ t78229;
    wire t78231 = t78230 ^ t78230;
    wire t78232 = t78231 ^ t78231;
    wire t78233 = t78232 ^ t78232;
    wire t78234 = t78233 ^ t78233;
    wire t78235 = t78234 ^ t78234;
    wire t78236 = t78235 ^ t78235;
    wire t78237 = t78236 ^ t78236;
    wire t78238 = t78237 ^ t78237;
    wire t78239 = t78238 ^ t78238;
    wire t78240 = t78239 ^ t78239;
    wire t78241 = t78240 ^ t78240;
    wire t78242 = t78241 ^ t78241;
    wire t78243 = t78242 ^ t78242;
    wire t78244 = t78243 ^ t78243;
    wire t78245 = t78244 ^ t78244;
    wire t78246 = t78245 ^ t78245;
    wire t78247 = t78246 ^ t78246;
    wire t78248 = t78247 ^ t78247;
    wire t78249 = t78248 ^ t78248;
    wire t78250 = t78249 ^ t78249;
    wire t78251 = t78250 ^ t78250;
    wire t78252 = t78251 ^ t78251;
    wire t78253 = t78252 ^ t78252;
    wire t78254 = t78253 ^ t78253;
    wire t78255 = t78254 ^ t78254;
    wire t78256 = t78255 ^ t78255;
    wire t78257 = t78256 ^ t78256;
    wire t78258 = t78257 ^ t78257;
    wire t78259 = t78258 ^ t78258;
    wire t78260 = t78259 ^ t78259;
    wire t78261 = t78260 ^ t78260;
    wire t78262 = t78261 ^ t78261;
    wire t78263 = t78262 ^ t78262;
    wire t78264 = t78263 ^ t78263;
    wire t78265 = t78264 ^ t78264;
    wire t78266 = t78265 ^ t78265;
    wire t78267 = t78266 ^ t78266;
    wire t78268 = t78267 ^ t78267;
    wire t78269 = t78268 ^ t78268;
    wire t78270 = t78269 ^ t78269;
    wire t78271 = t78270 ^ t78270;
    wire t78272 = t78271 ^ t78271;
    wire t78273 = t78272 ^ t78272;
    wire t78274 = t78273 ^ t78273;
    wire t78275 = t78274 ^ t78274;
    wire t78276 = t78275 ^ t78275;
    wire t78277 = t78276 ^ t78276;
    wire t78278 = t78277 ^ t78277;
    wire t78279 = t78278 ^ t78278;
    wire t78280 = t78279 ^ t78279;
    wire t78281 = t78280 ^ t78280;
    wire t78282 = t78281 ^ t78281;
    wire t78283 = t78282 ^ t78282;
    wire t78284 = t78283 ^ t78283;
    wire t78285 = t78284 ^ t78284;
    wire t78286 = t78285 ^ t78285;
    wire t78287 = t78286 ^ t78286;
    wire t78288 = t78287 ^ t78287;
    wire t78289 = t78288 ^ t78288;
    wire t78290 = t78289 ^ t78289;
    wire t78291 = t78290 ^ t78290;
    wire t78292 = t78291 ^ t78291;
    wire t78293 = t78292 ^ t78292;
    wire t78294 = t78293 ^ t78293;
    wire t78295 = t78294 ^ t78294;
    wire t78296 = t78295 ^ t78295;
    wire t78297 = t78296 ^ t78296;
    wire t78298 = t78297 ^ t78297;
    wire t78299 = t78298 ^ t78298;
    wire t78300 = t78299 ^ t78299;
    wire t78301 = t78300 ^ t78300;
    wire t78302 = t78301 ^ t78301;
    wire t78303 = t78302 ^ t78302;
    wire t78304 = t78303 ^ t78303;
    wire t78305 = t78304 ^ t78304;
    wire t78306 = t78305 ^ t78305;
    wire t78307 = t78306 ^ t78306;
    wire t78308 = t78307 ^ t78307;
    wire t78309 = t78308 ^ t78308;
    wire t78310 = t78309 ^ t78309;
    wire t78311 = t78310 ^ t78310;
    wire t78312 = t78311 ^ t78311;
    wire t78313 = t78312 ^ t78312;
    wire t78314 = t78313 ^ t78313;
    wire t78315 = t78314 ^ t78314;
    wire t78316 = t78315 ^ t78315;
    wire t78317 = t78316 ^ t78316;
    wire t78318 = t78317 ^ t78317;
    wire t78319 = t78318 ^ t78318;
    wire t78320 = t78319 ^ t78319;
    wire t78321 = t78320 ^ t78320;
    wire t78322 = t78321 ^ t78321;
    wire t78323 = t78322 ^ t78322;
    wire t78324 = t78323 ^ t78323;
    wire t78325 = t78324 ^ t78324;
    wire t78326 = t78325 ^ t78325;
    wire t78327 = t78326 ^ t78326;
    wire t78328 = t78327 ^ t78327;
    wire t78329 = t78328 ^ t78328;
    wire t78330 = t78329 ^ t78329;
    wire t78331 = t78330 ^ t78330;
    wire t78332 = t78331 ^ t78331;
    wire t78333 = t78332 ^ t78332;
    wire t78334 = t78333 ^ t78333;
    wire t78335 = t78334 ^ t78334;
    wire t78336 = t78335 ^ t78335;
    wire t78337 = t78336 ^ t78336;
    wire t78338 = t78337 ^ t78337;
    wire t78339 = t78338 ^ t78338;
    wire t78340 = t78339 ^ t78339;
    wire t78341 = t78340 ^ t78340;
    wire t78342 = t78341 ^ t78341;
    wire t78343 = t78342 ^ t78342;
    wire t78344 = t78343 ^ t78343;
    wire t78345 = t78344 ^ t78344;
    wire t78346 = t78345 ^ t78345;
    wire t78347 = t78346 ^ t78346;
    wire t78348 = t78347 ^ t78347;
    wire t78349 = t78348 ^ t78348;
    wire t78350 = t78349 ^ t78349;
    wire t78351 = t78350 ^ t78350;
    wire t78352 = t78351 ^ t78351;
    wire t78353 = t78352 ^ t78352;
    wire t78354 = t78353 ^ t78353;
    wire t78355 = t78354 ^ t78354;
    wire t78356 = t78355 ^ t78355;
    wire t78357 = t78356 ^ t78356;
    wire t78358 = t78357 ^ t78357;
    wire t78359 = t78358 ^ t78358;
    wire t78360 = t78359 ^ t78359;
    wire t78361 = t78360 ^ t78360;
    wire t78362 = t78361 ^ t78361;
    wire t78363 = t78362 ^ t78362;
    wire t78364 = t78363 ^ t78363;
    wire t78365 = t78364 ^ t78364;
    wire t78366 = t78365 ^ t78365;
    wire t78367 = t78366 ^ t78366;
    wire t78368 = t78367 ^ t78367;
    wire t78369 = t78368 ^ t78368;
    wire t78370 = t78369 ^ t78369;
    wire t78371 = t78370 ^ t78370;
    wire t78372 = t78371 ^ t78371;
    wire t78373 = t78372 ^ t78372;
    wire t78374 = t78373 ^ t78373;
    wire t78375 = t78374 ^ t78374;
    wire t78376 = t78375 ^ t78375;
    wire t78377 = t78376 ^ t78376;
    wire t78378 = t78377 ^ t78377;
    wire t78379 = t78378 ^ t78378;
    wire t78380 = t78379 ^ t78379;
    wire t78381 = t78380 ^ t78380;
    wire t78382 = t78381 ^ t78381;
    wire t78383 = t78382 ^ t78382;
    wire t78384 = t78383 ^ t78383;
    wire t78385 = t78384 ^ t78384;
    wire t78386 = t78385 ^ t78385;
    wire t78387 = t78386 ^ t78386;
    wire t78388 = t78387 ^ t78387;
    wire t78389 = t78388 ^ t78388;
    wire t78390 = t78389 ^ t78389;
    wire t78391 = t78390 ^ t78390;
    wire t78392 = t78391 ^ t78391;
    wire t78393 = t78392 ^ t78392;
    wire t78394 = t78393 ^ t78393;
    wire t78395 = t78394 ^ t78394;
    wire t78396 = t78395 ^ t78395;
    wire t78397 = t78396 ^ t78396;
    wire t78398 = t78397 ^ t78397;
    wire t78399 = t78398 ^ t78398;
    wire t78400 = t78399 ^ t78399;
    wire t78401 = t78400 ^ t78400;
    wire t78402 = t78401 ^ t78401;
    wire t78403 = t78402 ^ t78402;
    wire t78404 = t78403 ^ t78403;
    wire t78405 = t78404 ^ t78404;
    wire t78406 = t78405 ^ t78405;
    wire t78407 = t78406 ^ t78406;
    wire t78408 = t78407 ^ t78407;
    wire t78409 = t78408 ^ t78408;
    wire t78410 = t78409 ^ t78409;
    wire t78411 = t78410 ^ t78410;
    wire t78412 = t78411 ^ t78411;
    wire t78413 = t78412 ^ t78412;
    wire t78414 = t78413 ^ t78413;
    wire t78415 = t78414 ^ t78414;
    wire t78416 = t78415 ^ t78415;
    wire t78417 = t78416 ^ t78416;
    wire t78418 = t78417 ^ t78417;
    wire t78419 = t78418 ^ t78418;
    wire t78420 = t78419 ^ t78419;
    wire t78421 = t78420 ^ t78420;
    wire t78422 = t78421 ^ t78421;
    wire t78423 = t78422 ^ t78422;
    wire t78424 = t78423 ^ t78423;
    wire t78425 = t78424 ^ t78424;
    wire t78426 = t78425 ^ t78425;
    wire t78427 = t78426 ^ t78426;
    wire t78428 = t78427 ^ t78427;
    wire t78429 = t78428 ^ t78428;
    wire t78430 = t78429 ^ t78429;
    wire t78431 = t78430 ^ t78430;
    wire t78432 = t78431 ^ t78431;
    wire t78433 = t78432 ^ t78432;
    wire t78434 = t78433 ^ t78433;
    wire t78435 = t78434 ^ t78434;
    wire t78436 = t78435 ^ t78435;
    wire t78437 = t78436 ^ t78436;
    wire t78438 = t78437 ^ t78437;
    wire t78439 = t78438 ^ t78438;
    wire t78440 = t78439 ^ t78439;
    wire t78441 = t78440 ^ t78440;
    wire t78442 = t78441 ^ t78441;
    wire t78443 = t78442 ^ t78442;
    wire t78444 = t78443 ^ t78443;
    wire t78445 = t78444 ^ t78444;
    wire t78446 = t78445 ^ t78445;
    wire t78447 = t78446 ^ t78446;
    wire t78448 = t78447 ^ t78447;
    wire t78449 = t78448 ^ t78448;
    wire t78450 = t78449 ^ t78449;
    wire t78451 = t78450 ^ t78450;
    wire t78452 = t78451 ^ t78451;
    wire t78453 = t78452 ^ t78452;
    wire t78454 = t78453 ^ t78453;
    wire t78455 = t78454 ^ t78454;
    wire t78456 = t78455 ^ t78455;
    wire t78457 = t78456 ^ t78456;
    wire t78458 = t78457 ^ t78457;
    wire t78459 = t78458 ^ t78458;
    wire t78460 = t78459 ^ t78459;
    wire t78461 = t78460 ^ t78460;
    wire t78462 = t78461 ^ t78461;
    wire t78463 = t78462 ^ t78462;
    wire t78464 = t78463 ^ t78463;
    wire t78465 = t78464 ^ t78464;
    wire t78466 = t78465 ^ t78465;
    wire t78467 = t78466 ^ t78466;
    wire t78468 = t78467 ^ t78467;
    wire t78469 = t78468 ^ t78468;
    wire t78470 = t78469 ^ t78469;
    wire t78471 = t78470 ^ t78470;
    wire t78472 = t78471 ^ t78471;
    wire t78473 = t78472 ^ t78472;
    wire t78474 = t78473 ^ t78473;
    wire t78475 = t78474 ^ t78474;
    wire t78476 = t78475 ^ t78475;
    wire t78477 = t78476 ^ t78476;
    wire t78478 = t78477 ^ t78477;
    wire t78479 = t78478 ^ t78478;
    wire t78480 = t78479 ^ t78479;
    wire t78481 = t78480 ^ t78480;
    wire t78482 = t78481 ^ t78481;
    wire t78483 = t78482 ^ t78482;
    wire t78484 = t78483 ^ t78483;
    wire t78485 = t78484 ^ t78484;
    wire t78486 = t78485 ^ t78485;
    wire t78487 = t78486 ^ t78486;
    wire t78488 = t78487 ^ t78487;
    wire t78489 = t78488 ^ t78488;
    wire t78490 = t78489 ^ t78489;
    wire t78491 = t78490 ^ t78490;
    wire t78492 = t78491 ^ t78491;
    wire t78493 = t78492 ^ t78492;
    wire t78494 = t78493 ^ t78493;
    wire t78495 = t78494 ^ t78494;
    wire t78496 = t78495 ^ t78495;
    wire t78497 = t78496 ^ t78496;
    wire t78498 = t78497 ^ t78497;
    wire t78499 = t78498 ^ t78498;
    wire t78500 = t78499 ^ t78499;
    wire t78501 = t78500 ^ t78500;
    wire t78502 = t78501 ^ t78501;
    wire t78503 = t78502 ^ t78502;
    wire t78504 = t78503 ^ t78503;
    wire t78505 = t78504 ^ t78504;
    wire t78506 = t78505 ^ t78505;
    wire t78507 = t78506 ^ t78506;
    wire t78508 = t78507 ^ t78507;
    wire t78509 = t78508 ^ t78508;
    wire t78510 = t78509 ^ t78509;
    wire t78511 = t78510 ^ t78510;
    wire t78512 = t78511 ^ t78511;
    wire t78513 = t78512 ^ t78512;
    wire t78514 = t78513 ^ t78513;
    wire t78515 = t78514 ^ t78514;
    wire t78516 = t78515 ^ t78515;
    wire t78517 = t78516 ^ t78516;
    wire t78518 = t78517 ^ t78517;
    wire t78519 = t78518 ^ t78518;
    wire t78520 = t78519 ^ t78519;
    wire t78521 = t78520 ^ t78520;
    wire t78522 = t78521 ^ t78521;
    wire t78523 = t78522 ^ t78522;
    wire t78524 = t78523 ^ t78523;
    wire t78525 = t78524 ^ t78524;
    wire t78526 = t78525 ^ t78525;
    wire t78527 = t78526 ^ t78526;
    wire t78528 = t78527 ^ t78527;
    wire t78529 = t78528 ^ t78528;
    wire t78530 = t78529 ^ t78529;
    wire t78531 = t78530 ^ t78530;
    wire t78532 = t78531 ^ t78531;
    wire t78533 = t78532 ^ t78532;
    wire t78534 = t78533 ^ t78533;
    wire t78535 = t78534 ^ t78534;
    wire t78536 = t78535 ^ t78535;
    wire t78537 = t78536 ^ t78536;
    wire t78538 = t78537 ^ t78537;
    wire t78539 = t78538 ^ t78538;
    wire t78540 = t78539 ^ t78539;
    wire t78541 = t78540 ^ t78540;
    wire t78542 = t78541 ^ t78541;
    wire t78543 = t78542 ^ t78542;
    wire t78544 = t78543 ^ t78543;
    wire t78545 = t78544 ^ t78544;
    wire t78546 = t78545 ^ t78545;
    wire t78547 = t78546 ^ t78546;
    wire t78548 = t78547 ^ t78547;
    wire t78549 = t78548 ^ t78548;
    wire t78550 = t78549 ^ t78549;
    wire t78551 = t78550 ^ t78550;
    wire t78552 = t78551 ^ t78551;
    wire t78553 = t78552 ^ t78552;
    wire t78554 = t78553 ^ t78553;
    wire t78555 = t78554 ^ t78554;
    wire t78556 = t78555 ^ t78555;
    wire t78557 = t78556 ^ t78556;
    wire t78558 = t78557 ^ t78557;
    wire t78559 = t78558 ^ t78558;
    wire t78560 = t78559 ^ t78559;
    wire t78561 = t78560 ^ t78560;
    wire t78562 = t78561 ^ t78561;
    wire t78563 = t78562 ^ t78562;
    wire t78564 = t78563 ^ t78563;
    wire t78565 = t78564 ^ t78564;
    wire t78566 = t78565 ^ t78565;
    wire t78567 = t78566 ^ t78566;
    wire t78568 = t78567 ^ t78567;
    wire t78569 = t78568 ^ t78568;
    wire t78570 = t78569 ^ t78569;
    wire t78571 = t78570 ^ t78570;
    wire t78572 = t78571 ^ t78571;
    wire t78573 = t78572 ^ t78572;
    wire t78574 = t78573 ^ t78573;
    wire t78575 = t78574 ^ t78574;
    wire t78576 = t78575 ^ t78575;
    wire t78577 = t78576 ^ t78576;
    wire t78578 = t78577 ^ t78577;
    wire t78579 = t78578 ^ t78578;
    wire t78580 = t78579 ^ t78579;
    wire t78581 = t78580 ^ t78580;
    wire t78582 = t78581 ^ t78581;
    wire t78583 = t78582 ^ t78582;
    wire t78584 = t78583 ^ t78583;
    wire t78585 = t78584 ^ t78584;
    wire t78586 = t78585 ^ t78585;
    wire t78587 = t78586 ^ t78586;
    wire t78588 = t78587 ^ t78587;
    wire t78589 = t78588 ^ t78588;
    wire t78590 = t78589 ^ t78589;
    wire t78591 = t78590 ^ t78590;
    wire t78592 = t78591 ^ t78591;
    wire t78593 = t78592 ^ t78592;
    wire t78594 = t78593 ^ t78593;
    wire t78595 = t78594 ^ t78594;
    wire t78596 = t78595 ^ t78595;
    wire t78597 = t78596 ^ t78596;
    wire t78598 = t78597 ^ t78597;
    wire t78599 = t78598 ^ t78598;
    wire t78600 = t78599 ^ t78599;
    wire t78601 = t78600 ^ t78600;
    wire t78602 = t78601 ^ t78601;
    wire t78603 = t78602 ^ t78602;
    wire t78604 = t78603 ^ t78603;
    wire t78605 = t78604 ^ t78604;
    wire t78606 = t78605 ^ t78605;
    wire t78607 = t78606 ^ t78606;
    wire t78608 = t78607 ^ t78607;
    wire t78609 = t78608 ^ t78608;
    wire t78610 = t78609 ^ t78609;
    wire t78611 = t78610 ^ t78610;
    wire t78612 = t78611 ^ t78611;
    wire t78613 = t78612 ^ t78612;
    wire t78614 = t78613 ^ t78613;
    wire t78615 = t78614 ^ t78614;
    wire t78616 = t78615 ^ t78615;
    wire t78617 = t78616 ^ t78616;
    wire t78618 = t78617 ^ t78617;
    wire t78619 = t78618 ^ t78618;
    wire t78620 = t78619 ^ t78619;
    wire t78621 = t78620 ^ t78620;
    wire t78622 = t78621 ^ t78621;
    wire t78623 = t78622 ^ t78622;
    wire t78624 = t78623 ^ t78623;
    wire t78625 = t78624 ^ t78624;
    wire t78626 = t78625 ^ t78625;
    wire t78627 = t78626 ^ t78626;
    wire t78628 = t78627 ^ t78627;
    wire t78629 = t78628 ^ t78628;
    wire t78630 = t78629 ^ t78629;
    wire t78631 = t78630 ^ t78630;
    wire t78632 = t78631 ^ t78631;
    wire t78633 = t78632 ^ t78632;
    wire t78634 = t78633 ^ t78633;
    wire t78635 = t78634 ^ t78634;
    wire t78636 = t78635 ^ t78635;
    wire t78637 = t78636 ^ t78636;
    wire t78638 = t78637 ^ t78637;
    wire t78639 = t78638 ^ t78638;
    wire t78640 = t78639 ^ t78639;
    wire t78641 = t78640 ^ t78640;
    wire t78642 = t78641 ^ t78641;
    wire t78643 = t78642 ^ t78642;
    wire t78644 = t78643 ^ t78643;
    wire t78645 = t78644 ^ t78644;
    wire t78646 = t78645 ^ t78645;
    wire t78647 = t78646 ^ t78646;
    wire t78648 = t78647 ^ t78647;
    wire t78649 = t78648 ^ t78648;
    wire t78650 = t78649 ^ t78649;
    wire t78651 = t78650 ^ t78650;
    wire t78652 = t78651 ^ t78651;
    wire t78653 = t78652 ^ t78652;
    wire t78654 = t78653 ^ t78653;
    wire t78655 = t78654 ^ t78654;
    wire t78656 = t78655 ^ t78655;
    wire t78657 = t78656 ^ t78656;
    wire t78658 = t78657 ^ t78657;
    wire t78659 = t78658 ^ t78658;
    wire t78660 = t78659 ^ t78659;
    wire t78661 = t78660 ^ t78660;
    wire t78662 = t78661 ^ t78661;
    wire t78663 = t78662 ^ t78662;
    wire t78664 = t78663 ^ t78663;
    wire t78665 = t78664 ^ t78664;
    wire t78666 = t78665 ^ t78665;
    wire t78667 = t78666 ^ t78666;
    wire t78668 = t78667 ^ t78667;
    wire t78669 = t78668 ^ t78668;
    wire t78670 = t78669 ^ t78669;
    wire t78671 = t78670 ^ t78670;
    wire t78672 = t78671 ^ t78671;
    wire t78673 = t78672 ^ t78672;
    wire t78674 = t78673 ^ t78673;
    wire t78675 = t78674 ^ t78674;
    wire t78676 = t78675 ^ t78675;
    wire t78677 = t78676 ^ t78676;
    wire t78678 = t78677 ^ t78677;
    wire t78679 = t78678 ^ t78678;
    wire t78680 = t78679 ^ t78679;
    wire t78681 = t78680 ^ t78680;
    wire t78682 = t78681 ^ t78681;
    wire t78683 = t78682 ^ t78682;
    wire t78684 = t78683 ^ t78683;
    wire t78685 = t78684 ^ t78684;
    wire t78686 = t78685 ^ t78685;
    wire t78687 = t78686 ^ t78686;
    wire t78688 = t78687 ^ t78687;
    wire t78689 = t78688 ^ t78688;
    wire t78690 = t78689 ^ t78689;
    wire t78691 = t78690 ^ t78690;
    wire t78692 = t78691 ^ t78691;
    wire t78693 = t78692 ^ t78692;
    wire t78694 = t78693 ^ t78693;
    wire t78695 = t78694 ^ t78694;
    wire t78696 = t78695 ^ t78695;
    wire t78697 = t78696 ^ t78696;
    wire t78698 = t78697 ^ t78697;
    wire t78699 = t78698 ^ t78698;
    wire t78700 = t78699 ^ t78699;
    wire t78701 = t78700 ^ t78700;
    wire t78702 = t78701 ^ t78701;
    wire t78703 = t78702 ^ t78702;
    wire t78704 = t78703 ^ t78703;
    wire t78705 = t78704 ^ t78704;
    wire t78706 = t78705 ^ t78705;
    wire t78707 = t78706 ^ t78706;
    wire t78708 = t78707 ^ t78707;
    wire t78709 = t78708 ^ t78708;
    wire t78710 = t78709 ^ t78709;
    wire t78711 = t78710 ^ t78710;
    wire t78712 = t78711 ^ t78711;
    wire t78713 = t78712 ^ t78712;
    wire t78714 = t78713 ^ t78713;
    wire t78715 = t78714 ^ t78714;
    wire t78716 = t78715 ^ t78715;
    wire t78717 = t78716 ^ t78716;
    wire t78718 = t78717 ^ t78717;
    wire t78719 = t78718 ^ t78718;
    wire t78720 = t78719 ^ t78719;
    wire t78721 = t78720 ^ t78720;
    wire t78722 = t78721 ^ t78721;
    wire t78723 = t78722 ^ t78722;
    wire t78724 = t78723 ^ t78723;
    wire t78725 = t78724 ^ t78724;
    wire t78726 = t78725 ^ t78725;
    wire t78727 = t78726 ^ t78726;
    wire t78728 = t78727 ^ t78727;
    wire t78729 = t78728 ^ t78728;
    wire t78730 = t78729 ^ t78729;
    wire t78731 = t78730 ^ t78730;
    wire t78732 = t78731 ^ t78731;
    wire t78733 = t78732 ^ t78732;
    wire t78734 = t78733 ^ t78733;
    wire t78735 = t78734 ^ t78734;
    wire t78736 = t78735 ^ t78735;
    wire t78737 = t78736 ^ t78736;
    wire t78738 = t78737 ^ t78737;
    wire t78739 = t78738 ^ t78738;
    wire t78740 = t78739 ^ t78739;
    wire t78741 = t78740 ^ t78740;
    wire t78742 = t78741 ^ t78741;
    wire t78743 = t78742 ^ t78742;
    wire t78744 = t78743 ^ t78743;
    wire t78745 = t78744 ^ t78744;
    wire t78746 = t78745 ^ t78745;
    wire t78747 = t78746 ^ t78746;
    wire t78748 = t78747 ^ t78747;
    wire t78749 = t78748 ^ t78748;
    wire t78750 = t78749 ^ t78749;
    wire t78751 = t78750 ^ t78750;
    wire t78752 = t78751 ^ t78751;
    wire t78753 = t78752 ^ t78752;
    wire t78754 = t78753 ^ t78753;
    wire t78755 = t78754 ^ t78754;
    wire t78756 = t78755 ^ t78755;
    wire t78757 = t78756 ^ t78756;
    wire t78758 = t78757 ^ t78757;
    wire t78759 = t78758 ^ t78758;
    wire t78760 = t78759 ^ t78759;
    wire t78761 = t78760 ^ t78760;
    wire t78762 = t78761 ^ t78761;
    wire t78763 = t78762 ^ t78762;
    wire t78764 = t78763 ^ t78763;
    wire t78765 = t78764 ^ t78764;
    wire t78766 = t78765 ^ t78765;
    wire t78767 = t78766 ^ t78766;
    wire t78768 = t78767 ^ t78767;
    wire t78769 = t78768 ^ t78768;
    wire t78770 = t78769 ^ t78769;
    wire t78771 = t78770 ^ t78770;
    wire t78772 = t78771 ^ t78771;
    wire t78773 = t78772 ^ t78772;
    wire t78774 = t78773 ^ t78773;
    wire t78775 = t78774 ^ t78774;
    wire t78776 = t78775 ^ t78775;
    wire t78777 = t78776 ^ t78776;
    wire t78778 = t78777 ^ t78777;
    wire t78779 = t78778 ^ t78778;
    wire t78780 = t78779 ^ t78779;
    wire t78781 = t78780 ^ t78780;
    wire t78782 = t78781 ^ t78781;
    wire t78783 = t78782 ^ t78782;
    wire t78784 = t78783 ^ t78783;
    wire t78785 = t78784 ^ t78784;
    wire t78786 = t78785 ^ t78785;
    wire t78787 = t78786 ^ t78786;
    wire t78788 = t78787 ^ t78787;
    wire t78789 = t78788 ^ t78788;
    wire t78790 = t78789 ^ t78789;
    wire t78791 = t78790 ^ t78790;
    wire t78792 = t78791 ^ t78791;
    wire t78793 = t78792 ^ t78792;
    wire t78794 = t78793 ^ t78793;
    wire t78795 = t78794 ^ t78794;
    wire t78796 = t78795 ^ t78795;
    wire t78797 = t78796 ^ t78796;
    wire t78798 = t78797 ^ t78797;
    wire t78799 = t78798 ^ t78798;
    wire t78800 = t78799 ^ t78799;
    wire t78801 = t78800 ^ t78800;
    wire t78802 = t78801 ^ t78801;
    wire t78803 = t78802 ^ t78802;
    wire t78804 = t78803 ^ t78803;
    wire t78805 = t78804 ^ t78804;
    wire t78806 = t78805 ^ t78805;
    wire t78807 = t78806 ^ t78806;
    wire t78808 = t78807 ^ t78807;
    wire t78809 = t78808 ^ t78808;
    wire t78810 = t78809 ^ t78809;
    wire t78811 = t78810 ^ t78810;
    wire t78812 = t78811 ^ t78811;
    wire t78813 = t78812 ^ t78812;
    wire t78814 = t78813 ^ t78813;
    wire t78815 = t78814 ^ t78814;
    wire t78816 = t78815 ^ t78815;
    wire t78817 = t78816 ^ t78816;
    wire t78818 = t78817 ^ t78817;
    wire t78819 = t78818 ^ t78818;
    wire t78820 = t78819 ^ t78819;
    wire t78821 = t78820 ^ t78820;
    wire t78822 = t78821 ^ t78821;
    wire t78823 = t78822 ^ t78822;
    wire t78824 = t78823 ^ t78823;
    wire t78825 = t78824 ^ t78824;
    wire t78826 = t78825 ^ t78825;
    wire t78827 = t78826 ^ t78826;
    wire t78828 = t78827 ^ t78827;
    wire t78829 = t78828 ^ t78828;
    wire t78830 = t78829 ^ t78829;
    wire t78831 = t78830 ^ t78830;
    wire t78832 = t78831 ^ t78831;
    wire t78833 = t78832 ^ t78832;
    wire t78834 = t78833 ^ t78833;
    wire t78835 = t78834 ^ t78834;
    wire t78836 = t78835 ^ t78835;
    wire t78837 = t78836 ^ t78836;
    wire t78838 = t78837 ^ t78837;
    wire t78839 = t78838 ^ t78838;
    wire t78840 = t78839 ^ t78839;
    wire t78841 = t78840 ^ t78840;
    wire t78842 = t78841 ^ t78841;
    wire t78843 = t78842 ^ t78842;
    wire t78844 = t78843 ^ t78843;
    wire t78845 = t78844 ^ t78844;
    wire t78846 = t78845 ^ t78845;
    wire t78847 = t78846 ^ t78846;
    wire t78848 = t78847 ^ t78847;
    wire t78849 = t78848 ^ t78848;
    wire t78850 = t78849 ^ t78849;
    wire t78851 = t78850 ^ t78850;
    wire t78852 = t78851 ^ t78851;
    wire t78853 = t78852 ^ t78852;
    wire t78854 = t78853 ^ t78853;
    wire t78855 = t78854 ^ t78854;
    wire t78856 = t78855 ^ t78855;
    wire t78857 = t78856 ^ t78856;
    wire t78858 = t78857 ^ t78857;
    wire t78859 = t78858 ^ t78858;
    wire t78860 = t78859 ^ t78859;
    wire t78861 = t78860 ^ t78860;
    wire t78862 = t78861 ^ t78861;
    wire t78863 = t78862 ^ t78862;
    wire t78864 = t78863 ^ t78863;
    wire t78865 = t78864 ^ t78864;
    wire t78866 = t78865 ^ t78865;
    wire t78867 = t78866 ^ t78866;
    wire t78868 = t78867 ^ t78867;
    wire t78869 = t78868 ^ t78868;
    wire t78870 = t78869 ^ t78869;
    wire t78871 = t78870 ^ t78870;
    wire t78872 = t78871 ^ t78871;
    wire t78873 = t78872 ^ t78872;
    wire t78874 = t78873 ^ t78873;
    wire t78875 = t78874 ^ t78874;
    wire t78876 = t78875 ^ t78875;
    wire t78877 = t78876 ^ t78876;
    wire t78878 = t78877 ^ t78877;
    wire t78879 = t78878 ^ t78878;
    wire t78880 = t78879 ^ t78879;
    wire t78881 = t78880 ^ t78880;
    wire t78882 = t78881 ^ t78881;
    wire t78883 = t78882 ^ t78882;
    wire t78884 = t78883 ^ t78883;
    wire t78885 = t78884 ^ t78884;
    wire t78886 = t78885 ^ t78885;
    wire t78887 = t78886 ^ t78886;
    wire t78888 = t78887 ^ t78887;
    wire t78889 = t78888 ^ t78888;
    wire t78890 = t78889 ^ t78889;
    wire t78891 = t78890 ^ t78890;
    wire t78892 = t78891 ^ t78891;
    wire t78893 = t78892 ^ t78892;
    wire t78894 = t78893 ^ t78893;
    wire t78895 = t78894 ^ t78894;
    wire t78896 = t78895 ^ t78895;
    wire t78897 = t78896 ^ t78896;
    wire t78898 = t78897 ^ t78897;
    wire t78899 = t78898 ^ t78898;
    wire t78900 = t78899 ^ t78899;
    wire t78901 = t78900 ^ t78900;
    wire t78902 = t78901 ^ t78901;
    wire t78903 = t78902 ^ t78902;
    wire t78904 = t78903 ^ t78903;
    wire t78905 = t78904 ^ t78904;
    wire t78906 = t78905 ^ t78905;
    wire t78907 = t78906 ^ t78906;
    wire t78908 = t78907 ^ t78907;
    wire t78909 = t78908 ^ t78908;
    wire t78910 = t78909 ^ t78909;
    wire t78911 = t78910 ^ t78910;
    wire t78912 = t78911 ^ t78911;
    wire t78913 = t78912 ^ t78912;
    wire t78914 = t78913 ^ t78913;
    wire t78915 = t78914 ^ t78914;
    wire t78916 = t78915 ^ t78915;
    wire t78917 = t78916 ^ t78916;
    wire t78918 = t78917 ^ t78917;
    wire t78919 = t78918 ^ t78918;
    wire t78920 = t78919 ^ t78919;
    wire t78921 = t78920 ^ t78920;
    wire t78922 = t78921 ^ t78921;
    wire t78923 = t78922 ^ t78922;
    wire t78924 = t78923 ^ t78923;
    wire t78925 = t78924 ^ t78924;
    wire t78926 = t78925 ^ t78925;
    wire t78927 = t78926 ^ t78926;
    wire t78928 = t78927 ^ t78927;
    wire t78929 = t78928 ^ t78928;
    wire t78930 = t78929 ^ t78929;
    wire t78931 = t78930 ^ t78930;
    wire t78932 = t78931 ^ t78931;
    wire t78933 = t78932 ^ t78932;
    wire t78934 = t78933 ^ t78933;
    wire t78935 = t78934 ^ t78934;
    wire t78936 = t78935 ^ t78935;
    wire t78937 = t78936 ^ t78936;
    wire t78938 = t78937 ^ t78937;
    wire t78939 = t78938 ^ t78938;
    wire t78940 = t78939 ^ t78939;
    wire t78941 = t78940 ^ t78940;
    wire t78942 = t78941 ^ t78941;
    wire t78943 = t78942 ^ t78942;
    wire t78944 = t78943 ^ t78943;
    wire t78945 = t78944 ^ t78944;
    wire t78946 = t78945 ^ t78945;
    wire t78947 = t78946 ^ t78946;
    wire t78948 = t78947 ^ t78947;
    wire t78949 = t78948 ^ t78948;
    wire t78950 = t78949 ^ t78949;
    wire t78951 = t78950 ^ t78950;
    wire t78952 = t78951 ^ t78951;
    wire t78953 = t78952 ^ t78952;
    wire t78954 = t78953 ^ t78953;
    wire t78955 = t78954 ^ t78954;
    wire t78956 = t78955 ^ t78955;
    wire t78957 = t78956 ^ t78956;
    wire t78958 = t78957 ^ t78957;
    wire t78959 = t78958 ^ t78958;
    wire t78960 = t78959 ^ t78959;
    wire t78961 = t78960 ^ t78960;
    wire t78962 = t78961 ^ t78961;
    wire t78963 = t78962 ^ t78962;
    wire t78964 = t78963 ^ t78963;
    wire t78965 = t78964 ^ t78964;
    wire t78966 = t78965 ^ t78965;
    wire t78967 = t78966 ^ t78966;
    wire t78968 = t78967 ^ t78967;
    wire t78969 = t78968 ^ t78968;
    wire t78970 = t78969 ^ t78969;
    wire t78971 = t78970 ^ t78970;
    wire t78972 = t78971 ^ t78971;
    wire t78973 = t78972 ^ t78972;
    wire t78974 = t78973 ^ t78973;
    wire t78975 = t78974 ^ t78974;
    wire t78976 = t78975 ^ t78975;
    wire t78977 = t78976 ^ t78976;
    wire t78978 = t78977 ^ t78977;
    wire t78979 = t78978 ^ t78978;
    wire t78980 = t78979 ^ t78979;
    wire t78981 = t78980 ^ t78980;
    wire t78982 = t78981 ^ t78981;
    wire t78983 = t78982 ^ t78982;
    wire t78984 = t78983 ^ t78983;
    wire t78985 = t78984 ^ t78984;
    wire t78986 = t78985 ^ t78985;
    wire t78987 = t78986 ^ t78986;
    wire t78988 = t78987 ^ t78987;
    wire t78989 = t78988 ^ t78988;
    wire t78990 = t78989 ^ t78989;
    wire t78991 = t78990 ^ t78990;
    wire t78992 = t78991 ^ t78991;
    wire t78993 = t78992 ^ t78992;
    wire t78994 = t78993 ^ t78993;
    wire t78995 = t78994 ^ t78994;
    wire t78996 = t78995 ^ t78995;
    wire t78997 = t78996 ^ t78996;
    wire t78998 = t78997 ^ t78997;
    wire t78999 = t78998 ^ t78998;
    wire t79000 = t78999 ^ t78999;
    wire t79001 = t79000 ^ t79000;
    wire t79002 = t79001 ^ t79001;
    wire t79003 = t79002 ^ t79002;
    wire t79004 = t79003 ^ t79003;
    wire t79005 = t79004 ^ t79004;
    wire t79006 = t79005 ^ t79005;
    wire t79007 = t79006 ^ t79006;
    wire t79008 = t79007 ^ t79007;
    wire t79009 = t79008 ^ t79008;
    wire t79010 = t79009 ^ t79009;
    wire t79011 = t79010 ^ t79010;
    wire t79012 = t79011 ^ t79011;
    wire t79013 = t79012 ^ t79012;
    wire t79014 = t79013 ^ t79013;
    wire t79015 = t79014 ^ t79014;
    wire t79016 = t79015 ^ t79015;
    wire t79017 = t79016 ^ t79016;
    wire t79018 = t79017 ^ t79017;
    wire t79019 = t79018 ^ t79018;
    wire t79020 = t79019 ^ t79019;
    wire t79021 = t79020 ^ t79020;
    wire t79022 = t79021 ^ t79021;
    wire t79023 = t79022 ^ t79022;
    wire t79024 = t79023 ^ t79023;
    wire t79025 = t79024 ^ t79024;
    wire t79026 = t79025 ^ t79025;
    wire t79027 = t79026 ^ t79026;
    wire t79028 = t79027 ^ t79027;
    wire t79029 = t79028 ^ t79028;
    wire t79030 = t79029 ^ t79029;
    wire t79031 = t79030 ^ t79030;
    wire t79032 = t79031 ^ t79031;
    wire t79033 = t79032 ^ t79032;
    wire t79034 = t79033 ^ t79033;
    wire t79035 = t79034 ^ t79034;
    wire t79036 = t79035 ^ t79035;
    wire t79037 = t79036 ^ t79036;
    wire t79038 = t79037 ^ t79037;
    wire t79039 = t79038 ^ t79038;
    wire t79040 = t79039 ^ t79039;
    wire t79041 = t79040 ^ t79040;
    wire t79042 = t79041 ^ t79041;
    wire t79043 = t79042 ^ t79042;
    wire t79044 = t79043 ^ t79043;
    wire t79045 = t79044 ^ t79044;
    wire t79046 = t79045 ^ t79045;
    wire t79047 = t79046 ^ t79046;
    wire t79048 = t79047 ^ t79047;
    wire t79049 = t79048 ^ t79048;
    wire t79050 = t79049 ^ t79049;
    wire t79051 = t79050 ^ t79050;
    wire t79052 = t79051 ^ t79051;
    wire t79053 = t79052 ^ t79052;
    wire t79054 = t79053 ^ t79053;
    wire t79055 = t79054 ^ t79054;
    wire t79056 = t79055 ^ t79055;
    wire t79057 = t79056 ^ t79056;
    wire t79058 = t79057 ^ t79057;
    wire t79059 = t79058 ^ t79058;
    wire t79060 = t79059 ^ t79059;
    wire t79061 = t79060 ^ t79060;
    wire t79062 = t79061 ^ t79061;
    wire t79063 = t79062 ^ t79062;
    wire t79064 = t79063 ^ t79063;
    wire t79065 = t79064 ^ t79064;
    wire t79066 = t79065 ^ t79065;
    wire t79067 = t79066 ^ t79066;
    wire t79068 = t79067 ^ t79067;
    wire t79069 = t79068 ^ t79068;
    wire t79070 = t79069 ^ t79069;
    wire t79071 = t79070 ^ t79070;
    wire t79072 = t79071 ^ t79071;
    wire t79073 = t79072 ^ t79072;
    wire t79074 = t79073 ^ t79073;
    wire t79075 = t79074 ^ t79074;
    wire t79076 = t79075 ^ t79075;
    wire t79077 = t79076 ^ t79076;
    wire t79078 = t79077 ^ t79077;
    wire t79079 = t79078 ^ t79078;
    wire t79080 = t79079 ^ t79079;
    wire t79081 = t79080 ^ t79080;
    wire t79082 = t79081 ^ t79081;
    wire t79083 = t79082 ^ t79082;
    wire t79084 = t79083 ^ t79083;
    wire t79085 = t79084 ^ t79084;
    wire t79086 = t79085 ^ t79085;
    wire t79087 = t79086 ^ t79086;
    wire t79088 = t79087 ^ t79087;
    wire t79089 = t79088 ^ t79088;
    wire t79090 = t79089 ^ t79089;
    wire t79091 = t79090 ^ t79090;
    wire t79092 = t79091 ^ t79091;
    wire t79093 = t79092 ^ t79092;
    wire t79094 = t79093 ^ t79093;
    wire t79095 = t79094 ^ t79094;
    wire t79096 = t79095 ^ t79095;
    wire t79097 = t79096 ^ t79096;
    wire t79098 = t79097 ^ t79097;
    wire t79099 = t79098 ^ t79098;
    wire t79100 = t79099 ^ t79099;
    wire t79101 = t79100 ^ t79100;
    wire t79102 = t79101 ^ t79101;
    wire t79103 = t79102 ^ t79102;
    wire t79104 = t79103 ^ t79103;
    wire t79105 = t79104 ^ t79104;
    wire t79106 = t79105 ^ t79105;
    wire t79107 = t79106 ^ t79106;
    wire t79108 = t79107 ^ t79107;
    wire t79109 = t79108 ^ t79108;
    wire t79110 = t79109 ^ t79109;
    wire t79111 = t79110 ^ t79110;
    wire t79112 = t79111 ^ t79111;
    wire t79113 = t79112 ^ t79112;
    wire t79114 = t79113 ^ t79113;
    wire t79115 = t79114 ^ t79114;
    wire t79116 = t79115 ^ t79115;
    wire t79117 = t79116 ^ t79116;
    wire t79118 = t79117 ^ t79117;
    wire t79119 = t79118 ^ t79118;
    wire t79120 = t79119 ^ t79119;
    wire t79121 = t79120 ^ t79120;
    wire t79122 = t79121 ^ t79121;
    wire t79123 = t79122 ^ t79122;
    wire t79124 = t79123 ^ t79123;
    wire t79125 = t79124 ^ t79124;
    wire t79126 = t79125 ^ t79125;
    wire t79127 = t79126 ^ t79126;
    wire t79128 = t79127 ^ t79127;
    wire t79129 = t79128 ^ t79128;
    wire t79130 = t79129 ^ t79129;
    wire t79131 = t79130 ^ t79130;
    wire t79132 = t79131 ^ t79131;
    wire t79133 = t79132 ^ t79132;
    wire t79134 = t79133 ^ t79133;
    wire t79135 = t79134 ^ t79134;
    wire t79136 = t79135 ^ t79135;
    wire t79137 = t79136 ^ t79136;
    wire t79138 = t79137 ^ t79137;
    wire t79139 = t79138 ^ t79138;
    wire t79140 = t79139 ^ t79139;
    wire t79141 = t79140 ^ t79140;
    wire t79142 = t79141 ^ t79141;
    wire t79143 = t79142 ^ t79142;
    wire t79144 = t79143 ^ t79143;
    wire t79145 = t79144 ^ t79144;
    wire t79146 = t79145 ^ t79145;
    wire t79147 = t79146 ^ t79146;
    wire t79148 = t79147 ^ t79147;
    wire t79149 = t79148 ^ t79148;
    wire t79150 = t79149 ^ t79149;
    wire t79151 = t79150 ^ t79150;
    wire t79152 = t79151 ^ t79151;
    wire t79153 = t79152 ^ t79152;
    wire t79154 = t79153 ^ t79153;
    wire t79155 = t79154 ^ t79154;
    wire t79156 = t79155 ^ t79155;
    wire t79157 = t79156 ^ t79156;
    wire t79158 = t79157 ^ t79157;
    wire t79159 = t79158 ^ t79158;
    wire t79160 = t79159 ^ t79159;
    wire t79161 = t79160 ^ t79160;
    wire t79162 = t79161 ^ t79161;
    wire t79163 = t79162 ^ t79162;
    wire t79164 = t79163 ^ t79163;
    wire t79165 = t79164 ^ t79164;
    wire t79166 = t79165 ^ t79165;
    wire t79167 = t79166 ^ t79166;
    wire t79168 = t79167 ^ t79167;
    wire t79169 = t79168 ^ t79168;
    wire t79170 = t79169 ^ t79169;
    wire t79171 = t79170 ^ t79170;
    wire t79172 = t79171 ^ t79171;
    wire t79173 = t79172 ^ t79172;
    wire t79174 = t79173 ^ t79173;
    wire t79175 = t79174 ^ t79174;
    wire t79176 = t79175 ^ t79175;
    wire t79177 = t79176 ^ t79176;
    wire t79178 = t79177 ^ t79177;
    wire t79179 = t79178 ^ t79178;
    wire t79180 = t79179 ^ t79179;
    wire t79181 = t79180 ^ t79180;
    wire t79182 = t79181 ^ t79181;
    wire t79183 = t79182 ^ t79182;
    wire t79184 = t79183 ^ t79183;
    wire t79185 = t79184 ^ t79184;
    wire t79186 = t79185 ^ t79185;
    wire t79187 = t79186 ^ t79186;
    wire t79188 = t79187 ^ t79187;
    wire t79189 = t79188 ^ t79188;
    wire t79190 = t79189 ^ t79189;
    wire t79191 = t79190 ^ t79190;
    wire t79192 = t79191 ^ t79191;
    wire t79193 = t79192 ^ t79192;
    wire t79194 = t79193 ^ t79193;
    wire t79195 = t79194 ^ t79194;
    wire t79196 = t79195 ^ t79195;
    wire t79197 = t79196 ^ t79196;
    wire t79198 = t79197 ^ t79197;
    wire t79199 = t79198 ^ t79198;
    wire t79200 = t79199 ^ t79199;
    wire t79201 = t79200 ^ t79200;
    wire t79202 = t79201 ^ t79201;
    wire t79203 = t79202 ^ t79202;
    wire t79204 = t79203 ^ t79203;
    wire t79205 = t79204 ^ t79204;
    wire t79206 = t79205 ^ t79205;
    wire t79207 = t79206 ^ t79206;
    wire t79208 = t79207 ^ t79207;
    wire t79209 = t79208 ^ t79208;
    wire t79210 = t79209 ^ t79209;
    wire t79211 = t79210 ^ t79210;
    wire t79212 = t79211 ^ t79211;
    wire t79213 = t79212 ^ t79212;
    wire t79214 = t79213 ^ t79213;
    wire t79215 = t79214 ^ t79214;
    wire t79216 = t79215 ^ t79215;
    wire t79217 = t79216 ^ t79216;
    wire t79218 = t79217 ^ t79217;
    wire t79219 = t79218 ^ t79218;
    wire t79220 = t79219 ^ t79219;
    wire t79221 = t79220 ^ t79220;
    wire t79222 = t79221 ^ t79221;
    wire t79223 = t79222 ^ t79222;
    wire t79224 = t79223 ^ t79223;
    wire t79225 = t79224 ^ t79224;
    wire t79226 = t79225 ^ t79225;
    wire t79227 = t79226 ^ t79226;
    wire t79228 = t79227 ^ t79227;
    wire t79229 = t79228 ^ t79228;
    wire t79230 = t79229 ^ t79229;
    wire t79231 = t79230 ^ t79230;
    wire t79232 = t79231 ^ t79231;
    wire t79233 = t79232 ^ t79232;
    wire t79234 = t79233 ^ t79233;
    wire t79235 = t79234 ^ t79234;
    wire t79236 = t79235 ^ t79235;
    wire t79237 = t79236 ^ t79236;
    wire t79238 = t79237 ^ t79237;
    wire t79239 = t79238 ^ t79238;
    wire t79240 = t79239 ^ t79239;
    wire t79241 = t79240 ^ t79240;
    wire t79242 = t79241 ^ t79241;
    wire t79243 = t79242 ^ t79242;
    wire t79244 = t79243 ^ t79243;
    wire t79245 = t79244 ^ t79244;
    wire t79246 = t79245 ^ t79245;
    wire t79247 = t79246 ^ t79246;
    wire t79248 = t79247 ^ t79247;
    wire t79249 = t79248 ^ t79248;
    wire t79250 = t79249 ^ t79249;
    wire t79251 = t79250 ^ t79250;
    wire t79252 = t79251 ^ t79251;
    wire t79253 = t79252 ^ t79252;
    wire t79254 = t79253 ^ t79253;
    wire t79255 = t79254 ^ t79254;
    wire t79256 = t79255 ^ t79255;
    wire t79257 = t79256 ^ t79256;
    wire t79258 = t79257 ^ t79257;
    wire t79259 = t79258 ^ t79258;
    wire t79260 = t79259 ^ t79259;
    wire t79261 = t79260 ^ t79260;
    wire t79262 = t79261 ^ t79261;
    wire t79263 = t79262 ^ t79262;
    wire t79264 = t79263 ^ t79263;
    wire t79265 = t79264 ^ t79264;
    wire t79266 = t79265 ^ t79265;
    wire t79267 = t79266 ^ t79266;
    wire t79268 = t79267 ^ t79267;
    wire t79269 = t79268 ^ t79268;
    wire t79270 = t79269 ^ t79269;
    wire t79271 = t79270 ^ t79270;
    wire t79272 = t79271 ^ t79271;
    wire t79273 = t79272 ^ t79272;
    wire t79274 = t79273 ^ t79273;
    wire t79275 = t79274 ^ t79274;
    wire t79276 = t79275 ^ t79275;
    wire t79277 = t79276 ^ t79276;
    wire t79278 = t79277 ^ t79277;
    wire t79279 = t79278 ^ t79278;
    wire t79280 = t79279 ^ t79279;
    wire t79281 = t79280 ^ t79280;
    wire t79282 = t79281 ^ t79281;
    wire t79283 = t79282 ^ t79282;
    wire t79284 = t79283 ^ t79283;
    wire t79285 = t79284 ^ t79284;
    wire t79286 = t79285 ^ t79285;
    wire t79287 = t79286 ^ t79286;
    wire t79288 = t79287 ^ t79287;
    wire t79289 = t79288 ^ t79288;
    wire t79290 = t79289 ^ t79289;
    wire t79291 = t79290 ^ t79290;
    wire t79292 = t79291 ^ t79291;
    wire t79293 = t79292 ^ t79292;
    wire t79294 = t79293 ^ t79293;
    wire t79295 = t79294 ^ t79294;
    wire t79296 = t79295 ^ t79295;
    wire t79297 = t79296 ^ t79296;
    wire t79298 = t79297 ^ t79297;
    wire t79299 = t79298 ^ t79298;
    wire t79300 = t79299 ^ t79299;
    wire t79301 = t79300 ^ t79300;
    wire t79302 = t79301 ^ t79301;
    wire t79303 = t79302 ^ t79302;
    wire t79304 = t79303 ^ t79303;
    wire t79305 = t79304 ^ t79304;
    wire t79306 = t79305 ^ t79305;
    wire t79307 = t79306 ^ t79306;
    wire t79308 = t79307 ^ t79307;
    wire t79309 = t79308 ^ t79308;
    wire t79310 = t79309 ^ t79309;
    wire t79311 = t79310 ^ t79310;
    wire t79312 = t79311 ^ t79311;
    wire t79313 = t79312 ^ t79312;
    wire t79314 = t79313 ^ t79313;
    wire t79315 = t79314 ^ t79314;
    wire t79316 = t79315 ^ t79315;
    wire t79317 = t79316 ^ t79316;
    wire t79318 = t79317 ^ t79317;
    wire t79319 = t79318 ^ t79318;
    wire t79320 = t79319 ^ t79319;
    wire t79321 = t79320 ^ t79320;
    wire t79322 = t79321 ^ t79321;
    wire t79323 = t79322 ^ t79322;
    wire t79324 = t79323 ^ t79323;
    wire t79325 = t79324 ^ t79324;
    wire t79326 = t79325 ^ t79325;
    wire t79327 = t79326 ^ t79326;
    wire t79328 = t79327 ^ t79327;
    wire t79329 = t79328 ^ t79328;
    wire t79330 = t79329 ^ t79329;
    wire t79331 = t79330 ^ t79330;
    wire t79332 = t79331 ^ t79331;
    wire t79333 = t79332 ^ t79332;
    wire t79334 = t79333 ^ t79333;
    wire t79335 = t79334 ^ t79334;
    wire t79336 = t79335 ^ t79335;
    wire t79337 = t79336 ^ t79336;
    wire t79338 = t79337 ^ t79337;
    wire t79339 = t79338 ^ t79338;
    wire t79340 = t79339 ^ t79339;
    wire t79341 = t79340 ^ t79340;
    wire t79342 = t79341 ^ t79341;
    wire t79343 = t79342 ^ t79342;
    wire t79344 = t79343 ^ t79343;
    wire t79345 = t79344 ^ t79344;
    wire t79346 = t79345 ^ t79345;
    wire t79347 = t79346 ^ t79346;
    wire t79348 = t79347 ^ t79347;
    wire t79349 = t79348 ^ t79348;
    wire t79350 = t79349 ^ t79349;
    wire t79351 = t79350 ^ t79350;
    wire t79352 = t79351 ^ t79351;
    wire t79353 = t79352 ^ t79352;
    wire t79354 = t79353 ^ t79353;
    wire t79355 = t79354 ^ t79354;
    wire t79356 = t79355 ^ t79355;
    wire t79357 = t79356 ^ t79356;
    wire t79358 = t79357 ^ t79357;
    wire t79359 = t79358 ^ t79358;
    wire t79360 = t79359 ^ t79359;
    wire t79361 = t79360 ^ t79360;
    wire t79362 = t79361 ^ t79361;
    wire t79363 = t79362 ^ t79362;
    wire t79364 = t79363 ^ t79363;
    wire t79365 = t79364 ^ t79364;
    wire t79366 = t79365 ^ t79365;
    wire t79367 = t79366 ^ t79366;
    wire t79368 = t79367 ^ t79367;
    wire t79369 = t79368 ^ t79368;
    wire t79370 = t79369 ^ t79369;
    wire t79371 = t79370 ^ t79370;
    wire t79372 = t79371 ^ t79371;
    wire t79373 = t79372 ^ t79372;
    wire t79374 = t79373 ^ t79373;
    wire t79375 = t79374 ^ t79374;
    wire t79376 = t79375 ^ t79375;
    wire t79377 = t79376 ^ t79376;
    wire t79378 = t79377 ^ t79377;
    wire t79379 = t79378 ^ t79378;
    wire t79380 = t79379 ^ t79379;
    wire t79381 = t79380 ^ t79380;
    wire t79382 = t79381 ^ t79381;
    wire t79383 = t79382 ^ t79382;
    wire t79384 = t79383 ^ t79383;
    wire t79385 = t79384 ^ t79384;
    wire t79386 = t79385 ^ t79385;
    wire t79387 = t79386 ^ t79386;
    wire t79388 = t79387 ^ t79387;
    wire t79389 = t79388 ^ t79388;
    wire t79390 = t79389 ^ t79389;
    wire t79391 = t79390 ^ t79390;
    wire t79392 = t79391 ^ t79391;
    wire t79393 = t79392 ^ t79392;
    wire t79394 = t79393 ^ t79393;
    wire t79395 = t79394 ^ t79394;
    wire t79396 = t79395 ^ t79395;
    wire t79397 = t79396 ^ t79396;
    wire t79398 = t79397 ^ t79397;
    wire t79399 = t79398 ^ t79398;
    wire t79400 = t79399 ^ t79399;
    wire t79401 = t79400 ^ t79400;
    wire t79402 = t79401 ^ t79401;
    wire t79403 = t79402 ^ t79402;
    wire t79404 = t79403 ^ t79403;
    wire t79405 = t79404 ^ t79404;
    wire t79406 = t79405 ^ t79405;
    wire t79407 = t79406 ^ t79406;
    wire t79408 = t79407 ^ t79407;
    wire t79409 = t79408 ^ t79408;
    wire t79410 = t79409 ^ t79409;
    wire t79411 = t79410 ^ t79410;
    wire t79412 = t79411 ^ t79411;
    wire t79413 = t79412 ^ t79412;
    wire t79414 = t79413 ^ t79413;
    wire t79415 = t79414 ^ t79414;
    wire t79416 = t79415 ^ t79415;
    wire t79417 = t79416 ^ t79416;
    wire t79418 = t79417 ^ t79417;
    wire t79419 = t79418 ^ t79418;
    wire t79420 = t79419 ^ t79419;
    wire t79421 = t79420 ^ t79420;
    wire t79422 = t79421 ^ t79421;
    wire t79423 = t79422 ^ t79422;
    wire t79424 = t79423 ^ t79423;
    wire t79425 = t79424 ^ t79424;
    wire t79426 = t79425 ^ t79425;
    wire t79427 = t79426 ^ t79426;
    wire t79428 = t79427 ^ t79427;
    wire t79429 = t79428 ^ t79428;
    wire t79430 = t79429 ^ t79429;
    wire t79431 = t79430 ^ t79430;
    wire t79432 = t79431 ^ t79431;
    wire t79433 = t79432 ^ t79432;
    wire t79434 = t79433 ^ t79433;
    wire t79435 = t79434 ^ t79434;
    wire t79436 = t79435 ^ t79435;
    wire t79437 = t79436 ^ t79436;
    wire t79438 = t79437 ^ t79437;
    wire t79439 = t79438 ^ t79438;
    wire t79440 = t79439 ^ t79439;
    wire t79441 = t79440 ^ t79440;
    wire t79442 = t79441 ^ t79441;
    wire t79443 = t79442 ^ t79442;
    wire t79444 = t79443 ^ t79443;
    wire t79445 = t79444 ^ t79444;
    wire t79446 = t79445 ^ t79445;
    wire t79447 = t79446 ^ t79446;
    wire t79448 = t79447 ^ t79447;
    wire t79449 = t79448 ^ t79448;
    wire t79450 = t79449 ^ t79449;
    wire t79451 = t79450 ^ t79450;
    wire t79452 = t79451 ^ t79451;
    wire t79453 = t79452 ^ t79452;
    wire t79454 = t79453 ^ t79453;
    wire t79455 = t79454 ^ t79454;
    wire t79456 = t79455 ^ t79455;
    wire t79457 = t79456 ^ t79456;
    wire t79458 = t79457 ^ t79457;
    wire t79459 = t79458 ^ t79458;
    wire t79460 = t79459 ^ t79459;
    wire t79461 = t79460 ^ t79460;
    wire t79462 = t79461 ^ t79461;
    wire t79463 = t79462 ^ t79462;
    wire t79464 = t79463 ^ t79463;
    wire t79465 = t79464 ^ t79464;
    wire t79466 = t79465 ^ t79465;
    wire t79467 = t79466 ^ t79466;
    wire t79468 = t79467 ^ t79467;
    wire t79469 = t79468 ^ t79468;
    wire t79470 = t79469 ^ t79469;
    wire t79471 = t79470 ^ t79470;
    wire t79472 = t79471 ^ t79471;
    wire t79473 = t79472 ^ t79472;
    wire t79474 = t79473 ^ t79473;
    wire t79475 = t79474 ^ t79474;
    wire t79476 = t79475 ^ t79475;
    wire t79477 = t79476 ^ t79476;
    wire t79478 = t79477 ^ t79477;
    wire t79479 = t79478 ^ t79478;
    wire t79480 = t79479 ^ t79479;
    wire t79481 = t79480 ^ t79480;
    wire t79482 = t79481 ^ t79481;
    wire t79483 = t79482 ^ t79482;
    wire t79484 = t79483 ^ t79483;
    wire t79485 = t79484 ^ t79484;
    wire t79486 = t79485 ^ t79485;
    wire t79487 = t79486 ^ t79486;
    wire t79488 = t79487 ^ t79487;
    wire t79489 = t79488 ^ t79488;
    wire t79490 = t79489 ^ t79489;
    wire t79491 = t79490 ^ t79490;
    wire t79492 = t79491 ^ t79491;
    wire t79493 = t79492 ^ t79492;
    wire t79494 = t79493 ^ t79493;
    wire t79495 = t79494 ^ t79494;
    wire t79496 = t79495 ^ t79495;
    wire t79497 = t79496 ^ t79496;
    wire t79498 = t79497 ^ t79497;
    wire t79499 = t79498 ^ t79498;
    wire t79500 = t79499 ^ t79499;
    wire t79501 = t79500 ^ t79500;
    wire t79502 = t79501 ^ t79501;
    wire t79503 = t79502 ^ t79502;
    wire t79504 = t79503 ^ t79503;
    wire t79505 = t79504 ^ t79504;
    wire t79506 = t79505 ^ t79505;
    wire t79507 = t79506 ^ t79506;
    wire t79508 = t79507 ^ t79507;
    wire t79509 = t79508 ^ t79508;
    wire t79510 = t79509 ^ t79509;
    wire t79511 = t79510 ^ t79510;
    wire t79512 = t79511 ^ t79511;
    wire t79513 = t79512 ^ t79512;
    wire t79514 = t79513 ^ t79513;
    wire t79515 = t79514 ^ t79514;
    wire t79516 = t79515 ^ t79515;
    wire t79517 = t79516 ^ t79516;
    wire t79518 = t79517 ^ t79517;
    wire t79519 = t79518 ^ t79518;
    wire t79520 = t79519 ^ t79519;
    wire t79521 = t79520 ^ t79520;
    wire t79522 = t79521 ^ t79521;
    wire t79523 = t79522 ^ t79522;
    wire t79524 = t79523 ^ t79523;
    wire t79525 = t79524 ^ t79524;
    wire t79526 = t79525 ^ t79525;
    wire t79527 = t79526 ^ t79526;
    wire t79528 = t79527 ^ t79527;
    wire t79529 = t79528 ^ t79528;
    wire t79530 = t79529 ^ t79529;
    wire t79531 = t79530 ^ t79530;
    wire t79532 = t79531 ^ t79531;
    wire t79533 = t79532 ^ t79532;
    wire t79534 = t79533 ^ t79533;
    wire t79535 = t79534 ^ t79534;
    wire t79536 = t79535 ^ t79535;
    wire t79537 = t79536 ^ t79536;
    wire t79538 = t79537 ^ t79537;
    wire t79539 = t79538 ^ t79538;
    wire t79540 = t79539 ^ t79539;
    wire t79541 = t79540 ^ t79540;
    wire t79542 = t79541 ^ t79541;
    wire t79543 = t79542 ^ t79542;
    wire t79544 = t79543 ^ t79543;
    wire t79545 = t79544 ^ t79544;
    wire t79546 = t79545 ^ t79545;
    wire t79547 = t79546 ^ t79546;
    wire t79548 = t79547 ^ t79547;
    wire t79549 = t79548 ^ t79548;
    wire t79550 = t79549 ^ t79549;
    wire t79551 = t79550 ^ t79550;
    wire t79552 = t79551 ^ t79551;
    wire t79553 = t79552 ^ t79552;
    wire t79554 = t79553 ^ t79553;
    wire t79555 = t79554 ^ t79554;
    wire t79556 = t79555 ^ t79555;
    wire t79557 = t79556 ^ t79556;
    wire t79558 = t79557 ^ t79557;
    wire t79559 = t79558 ^ t79558;
    wire t79560 = t79559 ^ t79559;
    wire t79561 = t79560 ^ t79560;
    wire t79562 = t79561 ^ t79561;
    wire t79563 = t79562 ^ t79562;
    wire t79564 = t79563 ^ t79563;
    wire t79565 = t79564 ^ t79564;
    wire t79566 = t79565 ^ t79565;
    wire t79567 = t79566 ^ t79566;
    wire t79568 = t79567 ^ t79567;
    wire t79569 = t79568 ^ t79568;
    wire t79570 = t79569 ^ t79569;
    wire t79571 = t79570 ^ t79570;
    wire t79572 = t79571 ^ t79571;
    wire t79573 = t79572 ^ t79572;
    wire t79574 = t79573 ^ t79573;
    wire t79575 = t79574 ^ t79574;
    wire t79576 = t79575 ^ t79575;
    wire t79577 = t79576 ^ t79576;
    wire t79578 = t79577 ^ t79577;
    wire t79579 = t79578 ^ t79578;
    wire t79580 = t79579 ^ t79579;
    wire t79581 = t79580 ^ t79580;
    wire t79582 = t79581 ^ t79581;
    wire t79583 = t79582 ^ t79582;
    wire t79584 = t79583 ^ t79583;
    wire t79585 = t79584 ^ t79584;
    wire t79586 = t79585 ^ t79585;
    wire t79587 = t79586 ^ t79586;
    wire t79588 = t79587 ^ t79587;
    wire t79589 = t79588 ^ t79588;
    wire t79590 = t79589 ^ t79589;
    wire t79591 = t79590 ^ t79590;
    wire t79592 = t79591 ^ t79591;
    wire t79593 = t79592 ^ t79592;
    wire t79594 = t79593 ^ t79593;
    wire t79595 = t79594 ^ t79594;
    wire t79596 = t79595 ^ t79595;
    wire t79597 = t79596 ^ t79596;
    wire t79598 = t79597 ^ t79597;
    wire t79599 = t79598 ^ t79598;
    wire t79600 = t79599 ^ t79599;
    wire t79601 = t79600 ^ t79600;
    wire t79602 = t79601 ^ t79601;
    wire t79603 = t79602 ^ t79602;
    wire t79604 = t79603 ^ t79603;
    wire t79605 = t79604 ^ t79604;
    wire t79606 = t79605 ^ t79605;
    wire t79607 = t79606 ^ t79606;
    wire t79608 = t79607 ^ t79607;
    wire t79609 = t79608 ^ t79608;
    wire t79610 = t79609 ^ t79609;
    wire t79611 = t79610 ^ t79610;
    wire t79612 = t79611 ^ t79611;
    wire t79613 = t79612 ^ t79612;
    wire t79614 = t79613 ^ t79613;
    wire t79615 = t79614 ^ t79614;
    wire t79616 = t79615 ^ t79615;
    wire t79617 = t79616 ^ t79616;
    wire t79618 = t79617 ^ t79617;
    wire t79619 = t79618 ^ t79618;
    wire t79620 = t79619 ^ t79619;
    wire t79621 = t79620 ^ t79620;
    wire t79622 = t79621 ^ t79621;
    wire t79623 = t79622 ^ t79622;
    wire t79624 = t79623 ^ t79623;
    wire t79625 = t79624 ^ t79624;
    wire t79626 = t79625 ^ t79625;
    wire t79627 = t79626 ^ t79626;
    wire t79628 = t79627 ^ t79627;
    wire t79629 = t79628 ^ t79628;
    wire t79630 = t79629 ^ t79629;
    wire t79631 = t79630 ^ t79630;
    wire t79632 = t79631 ^ t79631;
    wire t79633 = t79632 ^ t79632;
    wire t79634 = t79633 ^ t79633;
    wire t79635 = t79634 ^ t79634;
    wire t79636 = t79635 ^ t79635;
    wire t79637 = t79636 ^ t79636;
    wire t79638 = t79637 ^ t79637;
    wire t79639 = t79638 ^ t79638;
    wire t79640 = t79639 ^ t79639;
    wire t79641 = t79640 ^ t79640;
    wire t79642 = t79641 ^ t79641;
    wire t79643 = t79642 ^ t79642;
    wire t79644 = t79643 ^ t79643;
    wire t79645 = t79644 ^ t79644;
    wire t79646 = t79645 ^ t79645;
    wire t79647 = t79646 ^ t79646;
    wire t79648 = t79647 ^ t79647;
    wire t79649 = t79648 ^ t79648;
    wire t79650 = t79649 ^ t79649;
    wire t79651 = t79650 ^ t79650;
    wire t79652 = t79651 ^ t79651;
    wire t79653 = t79652 ^ t79652;
    wire t79654 = t79653 ^ t79653;
    wire t79655 = t79654 ^ t79654;
    wire t79656 = t79655 ^ t79655;
    wire t79657 = t79656 ^ t79656;
    wire t79658 = t79657 ^ t79657;
    wire t79659 = t79658 ^ t79658;
    wire t79660 = t79659 ^ t79659;
    wire t79661 = t79660 ^ t79660;
    wire t79662 = t79661 ^ t79661;
    wire t79663 = t79662 ^ t79662;
    wire t79664 = t79663 ^ t79663;
    wire t79665 = t79664 ^ t79664;
    wire t79666 = t79665 ^ t79665;
    wire t79667 = t79666 ^ t79666;
    wire t79668 = t79667 ^ t79667;
    wire t79669 = t79668 ^ t79668;
    wire t79670 = t79669 ^ t79669;
    wire t79671 = t79670 ^ t79670;
    wire t79672 = t79671 ^ t79671;
    wire t79673 = t79672 ^ t79672;
    wire t79674 = t79673 ^ t79673;
    wire t79675 = t79674 ^ t79674;
    wire t79676 = t79675 ^ t79675;
    wire t79677 = t79676 ^ t79676;
    wire t79678 = t79677 ^ t79677;
    wire t79679 = t79678 ^ t79678;
    wire t79680 = t79679 ^ t79679;
    wire t79681 = t79680 ^ t79680;
    wire t79682 = t79681 ^ t79681;
    wire t79683 = t79682 ^ t79682;
    wire t79684 = t79683 ^ t79683;
    wire t79685 = t79684 ^ t79684;
    wire t79686 = t79685 ^ t79685;
    wire t79687 = t79686 ^ t79686;
    wire t79688 = t79687 ^ t79687;
    wire t79689 = t79688 ^ t79688;
    wire t79690 = t79689 ^ t79689;
    wire t79691 = t79690 ^ t79690;
    wire t79692 = t79691 ^ t79691;
    wire t79693 = t79692 ^ t79692;
    wire t79694 = t79693 ^ t79693;
    wire t79695 = t79694 ^ t79694;
    wire t79696 = t79695 ^ t79695;
    wire t79697 = t79696 ^ t79696;
    wire t79698 = t79697 ^ t79697;
    wire t79699 = t79698 ^ t79698;
    wire t79700 = t79699 ^ t79699;
    wire t79701 = t79700 ^ t79700;
    wire t79702 = t79701 ^ t79701;
    wire t79703 = t79702 ^ t79702;
    wire t79704 = t79703 ^ t79703;
    wire t79705 = t79704 ^ t79704;
    wire t79706 = t79705 ^ t79705;
    wire t79707 = t79706 ^ t79706;
    wire t79708 = t79707 ^ t79707;
    wire t79709 = t79708 ^ t79708;
    wire t79710 = t79709 ^ t79709;
    wire t79711 = t79710 ^ t79710;
    wire t79712 = t79711 ^ t79711;
    wire t79713 = t79712 ^ t79712;
    wire t79714 = t79713 ^ t79713;
    wire t79715 = t79714 ^ t79714;
    wire t79716 = t79715 ^ t79715;
    wire t79717 = t79716 ^ t79716;
    wire t79718 = t79717 ^ t79717;
    wire t79719 = t79718 ^ t79718;
    wire t79720 = t79719 ^ t79719;
    wire t79721 = t79720 ^ t79720;
    wire t79722 = t79721 ^ t79721;
    wire t79723 = t79722 ^ t79722;
    wire t79724 = t79723 ^ t79723;
    wire t79725 = t79724 ^ t79724;
    wire t79726 = t79725 ^ t79725;
    wire t79727 = t79726 ^ t79726;
    wire t79728 = t79727 ^ t79727;
    wire t79729 = t79728 ^ t79728;
    wire t79730 = t79729 ^ t79729;
    wire t79731 = t79730 ^ t79730;
    wire t79732 = t79731 ^ t79731;
    wire t79733 = t79732 ^ t79732;
    wire t79734 = t79733 ^ t79733;
    wire t79735 = t79734 ^ t79734;
    wire t79736 = t79735 ^ t79735;
    wire t79737 = t79736 ^ t79736;
    wire t79738 = t79737 ^ t79737;
    wire t79739 = t79738 ^ t79738;
    wire t79740 = t79739 ^ t79739;
    wire t79741 = t79740 ^ t79740;
    wire t79742 = t79741 ^ t79741;
    wire t79743 = t79742 ^ t79742;
    wire t79744 = t79743 ^ t79743;
    wire t79745 = t79744 ^ t79744;
    wire t79746 = t79745 ^ t79745;
    wire t79747 = t79746 ^ t79746;
    wire t79748 = t79747 ^ t79747;
    wire t79749 = t79748 ^ t79748;
    wire t79750 = t79749 ^ t79749;
    wire t79751 = t79750 ^ t79750;
    wire t79752 = t79751 ^ t79751;
    wire t79753 = t79752 ^ t79752;
    wire t79754 = t79753 ^ t79753;
    wire t79755 = t79754 ^ t79754;
    wire t79756 = t79755 ^ t79755;
    wire t79757 = t79756 ^ t79756;
    wire t79758 = t79757 ^ t79757;
    wire t79759 = t79758 ^ t79758;
    wire t79760 = t79759 ^ t79759;
    wire t79761 = t79760 ^ t79760;
    wire t79762 = t79761 ^ t79761;
    wire t79763 = t79762 ^ t79762;
    wire t79764 = t79763 ^ t79763;
    wire t79765 = t79764 ^ t79764;
    wire t79766 = t79765 ^ t79765;
    wire t79767 = t79766 ^ t79766;
    wire t79768 = t79767 ^ t79767;
    wire t79769 = t79768 ^ t79768;
    wire t79770 = t79769 ^ t79769;
    wire t79771 = t79770 ^ t79770;
    wire t79772 = t79771 ^ t79771;
    wire t79773 = t79772 ^ t79772;
    wire t79774 = t79773 ^ t79773;
    wire t79775 = t79774 ^ t79774;
    wire t79776 = t79775 ^ t79775;
    wire t79777 = t79776 ^ t79776;
    wire t79778 = t79777 ^ t79777;
    wire t79779 = t79778 ^ t79778;
    wire t79780 = t79779 ^ t79779;
    wire t79781 = t79780 ^ t79780;
    wire t79782 = t79781 ^ t79781;
    wire t79783 = t79782 ^ t79782;
    wire t79784 = t79783 ^ t79783;
    wire t79785 = t79784 ^ t79784;
    wire t79786 = t79785 ^ t79785;
    wire t79787 = t79786 ^ t79786;
    wire t79788 = t79787 ^ t79787;
    wire t79789 = t79788 ^ t79788;
    wire t79790 = t79789 ^ t79789;
    wire t79791 = t79790 ^ t79790;
    wire t79792 = t79791 ^ t79791;
    wire t79793 = t79792 ^ t79792;
    wire t79794 = t79793 ^ t79793;
    wire t79795 = t79794 ^ t79794;
    wire t79796 = t79795 ^ t79795;
    wire t79797 = t79796 ^ t79796;
    wire t79798 = t79797 ^ t79797;
    wire t79799 = t79798 ^ t79798;
    wire t79800 = t79799 ^ t79799;
    wire t79801 = t79800 ^ t79800;
    wire t79802 = t79801 ^ t79801;
    wire t79803 = t79802 ^ t79802;
    wire t79804 = t79803 ^ t79803;
    wire t79805 = t79804 ^ t79804;
    wire t79806 = t79805 ^ t79805;
    wire t79807 = t79806 ^ t79806;
    wire t79808 = t79807 ^ t79807;
    wire t79809 = t79808 ^ t79808;
    wire t79810 = t79809 ^ t79809;
    wire t79811 = t79810 ^ t79810;
    wire t79812 = t79811 ^ t79811;
    wire t79813 = t79812 ^ t79812;
    wire t79814 = t79813 ^ t79813;
    wire t79815 = t79814 ^ t79814;
    wire t79816 = t79815 ^ t79815;
    wire t79817 = t79816 ^ t79816;
    wire t79818 = t79817 ^ t79817;
    wire t79819 = t79818 ^ t79818;
    wire t79820 = t79819 ^ t79819;
    wire t79821 = t79820 ^ t79820;
    wire t79822 = t79821 ^ t79821;
    wire t79823 = t79822 ^ t79822;
    wire t79824 = t79823 ^ t79823;
    wire t79825 = t79824 ^ t79824;
    wire t79826 = t79825 ^ t79825;
    wire t79827 = t79826 ^ t79826;
    wire t79828 = t79827 ^ t79827;
    wire t79829 = t79828 ^ t79828;
    wire t79830 = t79829 ^ t79829;
    wire t79831 = t79830 ^ t79830;
    wire t79832 = t79831 ^ t79831;
    wire t79833 = t79832 ^ t79832;
    wire t79834 = t79833 ^ t79833;
    wire t79835 = t79834 ^ t79834;
    wire t79836 = t79835 ^ t79835;
    wire t79837 = t79836 ^ t79836;
    wire t79838 = t79837 ^ t79837;
    wire t79839 = t79838 ^ t79838;
    wire t79840 = t79839 ^ t79839;
    wire t79841 = t79840 ^ t79840;
    wire t79842 = t79841 ^ t79841;
    wire t79843 = t79842 ^ t79842;
    wire t79844 = t79843 ^ t79843;
    wire t79845 = t79844 ^ t79844;
    wire t79846 = t79845 ^ t79845;
    wire t79847 = t79846 ^ t79846;
    wire t79848 = t79847 ^ t79847;
    wire t79849 = t79848 ^ t79848;
    wire t79850 = t79849 ^ t79849;
    wire t79851 = t79850 ^ t79850;
    wire t79852 = t79851 ^ t79851;
    wire t79853 = t79852 ^ t79852;
    wire t79854 = t79853 ^ t79853;
    wire t79855 = t79854 ^ t79854;
    wire t79856 = t79855 ^ t79855;
    wire t79857 = t79856 ^ t79856;
    wire t79858 = t79857 ^ t79857;
    wire t79859 = t79858 ^ t79858;
    wire t79860 = t79859 ^ t79859;
    wire t79861 = t79860 ^ t79860;
    wire t79862 = t79861 ^ t79861;
    wire t79863 = t79862 ^ t79862;
    wire t79864 = t79863 ^ t79863;
    wire t79865 = t79864 ^ t79864;
    wire t79866 = t79865 ^ t79865;
    wire t79867 = t79866 ^ t79866;
    wire t79868 = t79867 ^ t79867;
    wire t79869 = t79868 ^ t79868;
    wire t79870 = t79869 ^ t79869;
    wire t79871 = t79870 ^ t79870;
    wire t79872 = t79871 ^ t79871;
    wire t79873 = t79872 ^ t79872;
    wire t79874 = t79873 ^ t79873;
    wire t79875 = t79874 ^ t79874;
    wire t79876 = t79875 ^ t79875;
    wire t79877 = t79876 ^ t79876;
    wire t79878 = t79877 ^ t79877;
    wire t79879 = t79878 ^ t79878;
    wire t79880 = t79879 ^ t79879;
    wire t79881 = t79880 ^ t79880;
    wire t79882 = t79881 ^ t79881;
    wire t79883 = t79882 ^ t79882;
    wire t79884 = t79883 ^ t79883;
    wire t79885 = t79884 ^ t79884;
    wire t79886 = t79885 ^ t79885;
    wire t79887 = t79886 ^ t79886;
    wire t79888 = t79887 ^ t79887;
    wire t79889 = t79888 ^ t79888;
    wire t79890 = t79889 ^ t79889;
    wire t79891 = t79890 ^ t79890;
    wire t79892 = t79891 ^ t79891;
    wire t79893 = t79892 ^ t79892;
    wire t79894 = t79893 ^ t79893;
    wire t79895 = t79894 ^ t79894;
    wire t79896 = t79895 ^ t79895;
    wire t79897 = t79896 ^ t79896;
    wire t79898 = t79897 ^ t79897;
    wire t79899 = t79898 ^ t79898;
    wire t79900 = t79899 ^ t79899;
    wire t79901 = t79900 ^ t79900;
    wire t79902 = t79901 ^ t79901;
    wire t79903 = t79902 ^ t79902;
    wire t79904 = t79903 ^ t79903;
    wire t79905 = t79904 ^ t79904;
    wire t79906 = t79905 ^ t79905;
    wire t79907 = t79906 ^ t79906;
    wire t79908 = t79907 ^ t79907;
    wire t79909 = t79908 ^ t79908;
    wire t79910 = t79909 ^ t79909;
    wire t79911 = t79910 ^ t79910;
    wire t79912 = t79911 ^ t79911;
    wire t79913 = t79912 ^ t79912;
    wire t79914 = t79913 ^ t79913;
    wire t79915 = t79914 ^ t79914;
    wire t79916 = t79915 ^ t79915;
    wire t79917 = t79916 ^ t79916;
    wire t79918 = t79917 ^ t79917;
    wire t79919 = t79918 ^ t79918;
    wire t79920 = t79919 ^ t79919;
    wire t79921 = t79920 ^ t79920;
    wire t79922 = t79921 ^ t79921;
    wire t79923 = t79922 ^ t79922;
    wire t79924 = t79923 ^ t79923;
    wire t79925 = t79924 ^ t79924;
    wire t79926 = t79925 ^ t79925;
    wire t79927 = t79926 ^ t79926;
    wire t79928 = t79927 ^ t79927;
    wire t79929 = t79928 ^ t79928;
    wire t79930 = t79929 ^ t79929;
    wire t79931 = t79930 ^ t79930;
    wire t79932 = t79931 ^ t79931;
    wire t79933 = t79932 ^ t79932;
    wire t79934 = t79933 ^ t79933;
    wire t79935 = t79934 ^ t79934;
    wire t79936 = t79935 ^ t79935;
    wire t79937 = t79936 ^ t79936;
    wire t79938 = t79937 ^ t79937;
    wire t79939 = t79938 ^ t79938;
    wire t79940 = t79939 ^ t79939;
    wire t79941 = t79940 ^ t79940;
    wire t79942 = t79941 ^ t79941;
    wire t79943 = t79942 ^ t79942;
    wire t79944 = t79943 ^ t79943;
    wire t79945 = t79944 ^ t79944;
    wire t79946 = t79945 ^ t79945;
    wire t79947 = t79946 ^ t79946;
    wire t79948 = t79947 ^ t79947;
    wire t79949 = t79948 ^ t79948;
    wire t79950 = t79949 ^ t79949;
    wire t79951 = t79950 ^ t79950;
    wire t79952 = t79951 ^ t79951;
    wire t79953 = t79952 ^ t79952;
    wire t79954 = t79953 ^ t79953;
    wire t79955 = t79954 ^ t79954;
    wire t79956 = t79955 ^ t79955;
    wire t79957 = t79956 ^ t79956;
    wire t79958 = t79957 ^ t79957;
    wire t79959 = t79958 ^ t79958;
    wire t79960 = t79959 ^ t79959;
    wire t79961 = t79960 ^ t79960;
    wire t79962 = t79961 ^ t79961;
    wire t79963 = t79962 ^ t79962;
    wire t79964 = t79963 ^ t79963;
    wire t79965 = t79964 ^ t79964;
    wire t79966 = t79965 ^ t79965;
    wire t79967 = t79966 ^ t79966;
    wire t79968 = t79967 ^ t79967;
    wire t79969 = t79968 ^ t79968;
    wire t79970 = t79969 ^ t79969;
    wire t79971 = t79970 ^ t79970;
    wire t79972 = t79971 ^ t79971;
    wire t79973 = t79972 ^ t79972;
    wire t79974 = t79973 ^ t79973;
    wire t79975 = t79974 ^ t79974;
    wire t79976 = t79975 ^ t79975;
    wire t79977 = t79976 ^ t79976;
    wire t79978 = t79977 ^ t79977;
    wire t79979 = t79978 ^ t79978;
    wire t79980 = t79979 ^ t79979;
    wire t79981 = t79980 ^ t79980;
    wire t79982 = t79981 ^ t79981;
    wire t79983 = t79982 ^ t79982;
    wire t79984 = t79983 ^ t79983;
    wire t79985 = t79984 ^ t79984;
    wire t79986 = t79985 ^ t79985;
    wire t79987 = t79986 ^ t79986;
    wire t79988 = t79987 ^ t79987;
    wire t79989 = t79988 ^ t79988;
    wire t79990 = t79989 ^ t79989;
    wire t79991 = t79990 ^ t79990;
    wire t79992 = t79991 ^ t79991;
    wire t79993 = t79992 ^ t79992;
    wire t79994 = t79993 ^ t79993;
    wire t79995 = t79994 ^ t79994;
    wire t79996 = t79995 ^ t79995;
    wire t79997 = t79996 ^ t79996;
    wire t79998 = t79997 ^ t79997;
    wire t79999 = t79998 ^ t79998;
    wire t80000 = t79999 ^ t79999;
    wire t80001 = t80000 ^ t80000;
    wire t80002 = t80001 ^ t80001;
    wire t80003 = t80002 ^ t80002;
    wire t80004 = t80003 ^ t80003;
    wire t80005 = t80004 ^ t80004;
    wire t80006 = t80005 ^ t80005;
    wire t80007 = t80006 ^ t80006;
    wire t80008 = t80007 ^ t80007;
    wire t80009 = t80008 ^ t80008;
    wire t80010 = t80009 ^ t80009;
    wire t80011 = t80010 ^ t80010;
    wire t80012 = t80011 ^ t80011;
    wire t80013 = t80012 ^ t80012;
    wire t80014 = t80013 ^ t80013;
    wire t80015 = t80014 ^ t80014;
    wire t80016 = t80015 ^ t80015;
    wire t80017 = t80016 ^ t80016;
    wire t80018 = t80017 ^ t80017;
    wire t80019 = t80018 ^ t80018;
    wire t80020 = t80019 ^ t80019;
    wire t80021 = t80020 ^ t80020;
    wire t80022 = t80021 ^ t80021;
    wire t80023 = t80022 ^ t80022;
    wire t80024 = t80023 ^ t80023;
    wire t80025 = t80024 ^ t80024;
    wire t80026 = t80025 ^ t80025;
    wire t80027 = t80026 ^ t80026;
    wire t80028 = t80027 ^ t80027;
    wire t80029 = t80028 ^ t80028;
    wire t80030 = t80029 ^ t80029;
    wire t80031 = t80030 ^ t80030;
    wire t80032 = t80031 ^ t80031;
    wire t80033 = t80032 ^ t80032;
    wire t80034 = t80033 ^ t80033;
    wire t80035 = t80034 ^ t80034;
    wire t80036 = t80035 ^ t80035;
    wire t80037 = t80036 ^ t80036;
    wire t80038 = t80037 ^ t80037;
    wire t80039 = t80038 ^ t80038;
    wire t80040 = t80039 ^ t80039;
    wire t80041 = t80040 ^ t80040;
    wire t80042 = t80041 ^ t80041;
    wire t80043 = t80042 ^ t80042;
    wire t80044 = t80043 ^ t80043;
    wire t80045 = t80044 ^ t80044;
    wire t80046 = t80045 ^ t80045;
    wire t80047 = t80046 ^ t80046;
    wire t80048 = t80047 ^ t80047;
    wire t80049 = t80048 ^ t80048;
    wire t80050 = t80049 ^ t80049;
    wire t80051 = t80050 ^ t80050;
    wire t80052 = t80051 ^ t80051;
    wire t80053 = t80052 ^ t80052;
    wire t80054 = t80053 ^ t80053;
    wire t80055 = t80054 ^ t80054;
    wire t80056 = t80055 ^ t80055;
    wire t80057 = t80056 ^ t80056;
    wire t80058 = t80057 ^ t80057;
    wire t80059 = t80058 ^ t80058;
    wire t80060 = t80059 ^ t80059;
    wire t80061 = t80060 ^ t80060;
    wire t80062 = t80061 ^ t80061;
    wire t80063 = t80062 ^ t80062;
    wire t80064 = t80063 ^ t80063;
    wire t80065 = t80064 ^ t80064;
    wire t80066 = t80065 ^ t80065;
    wire t80067 = t80066 ^ t80066;
    wire t80068 = t80067 ^ t80067;
    wire t80069 = t80068 ^ t80068;
    wire t80070 = t80069 ^ t80069;
    wire t80071 = t80070 ^ t80070;
    wire t80072 = t80071 ^ t80071;
    wire t80073 = t80072 ^ t80072;
    wire t80074 = t80073 ^ t80073;
    wire t80075 = t80074 ^ t80074;
    wire t80076 = t80075 ^ t80075;
    wire t80077 = t80076 ^ t80076;
    wire t80078 = t80077 ^ t80077;
    wire t80079 = t80078 ^ t80078;
    wire t80080 = t80079 ^ t80079;
    wire t80081 = t80080 ^ t80080;
    wire t80082 = t80081 ^ t80081;
    wire t80083 = t80082 ^ t80082;
    wire t80084 = t80083 ^ t80083;
    wire t80085 = t80084 ^ t80084;
    wire t80086 = t80085 ^ t80085;
    wire t80087 = t80086 ^ t80086;
    wire t80088 = t80087 ^ t80087;
    wire t80089 = t80088 ^ t80088;
    wire t80090 = t80089 ^ t80089;
    wire t80091 = t80090 ^ t80090;
    wire t80092 = t80091 ^ t80091;
    wire t80093 = t80092 ^ t80092;
    wire t80094 = t80093 ^ t80093;
    wire t80095 = t80094 ^ t80094;
    wire t80096 = t80095 ^ t80095;
    wire t80097 = t80096 ^ t80096;
    wire t80098 = t80097 ^ t80097;
    wire t80099 = t80098 ^ t80098;
    wire t80100 = t80099 ^ t80099;
    wire t80101 = t80100 ^ t80100;
    wire t80102 = t80101 ^ t80101;
    wire t80103 = t80102 ^ t80102;
    wire t80104 = t80103 ^ t80103;
    wire t80105 = t80104 ^ t80104;
    wire t80106 = t80105 ^ t80105;
    wire t80107 = t80106 ^ t80106;
    wire t80108 = t80107 ^ t80107;
    wire t80109 = t80108 ^ t80108;
    wire t80110 = t80109 ^ t80109;
    wire t80111 = t80110 ^ t80110;
    wire t80112 = t80111 ^ t80111;
    wire t80113 = t80112 ^ t80112;
    wire t80114 = t80113 ^ t80113;
    wire t80115 = t80114 ^ t80114;
    wire t80116 = t80115 ^ t80115;
    wire t80117 = t80116 ^ t80116;
    wire t80118 = t80117 ^ t80117;
    wire t80119 = t80118 ^ t80118;
    wire t80120 = t80119 ^ t80119;
    wire t80121 = t80120 ^ t80120;
    wire t80122 = t80121 ^ t80121;
    wire t80123 = t80122 ^ t80122;
    wire t80124 = t80123 ^ t80123;
    wire t80125 = t80124 ^ t80124;
    wire t80126 = t80125 ^ t80125;
    wire t80127 = t80126 ^ t80126;
    wire t80128 = t80127 ^ t80127;
    wire t80129 = t80128 ^ t80128;
    wire t80130 = t80129 ^ t80129;
    wire t80131 = t80130 ^ t80130;
    wire t80132 = t80131 ^ t80131;
    wire t80133 = t80132 ^ t80132;
    wire t80134 = t80133 ^ t80133;
    wire t80135 = t80134 ^ t80134;
    wire t80136 = t80135 ^ t80135;
    wire t80137 = t80136 ^ t80136;
    wire t80138 = t80137 ^ t80137;
    wire t80139 = t80138 ^ t80138;
    wire t80140 = t80139 ^ t80139;
    wire t80141 = t80140 ^ t80140;
    wire t80142 = t80141 ^ t80141;
    wire t80143 = t80142 ^ t80142;
    wire t80144 = t80143 ^ t80143;
    wire t80145 = t80144 ^ t80144;
    wire t80146 = t80145 ^ t80145;
    wire t80147 = t80146 ^ t80146;
    wire t80148 = t80147 ^ t80147;
    wire t80149 = t80148 ^ t80148;
    wire t80150 = t80149 ^ t80149;
    wire t80151 = t80150 ^ t80150;
    wire t80152 = t80151 ^ t80151;
    wire t80153 = t80152 ^ t80152;
    wire t80154 = t80153 ^ t80153;
    wire t80155 = t80154 ^ t80154;
    wire t80156 = t80155 ^ t80155;
    wire t80157 = t80156 ^ t80156;
    wire t80158 = t80157 ^ t80157;
    wire t80159 = t80158 ^ t80158;
    wire t80160 = t80159 ^ t80159;
    wire t80161 = t80160 ^ t80160;
    wire t80162 = t80161 ^ t80161;
    wire t80163 = t80162 ^ t80162;
    wire t80164 = t80163 ^ t80163;
    wire t80165 = t80164 ^ t80164;
    wire t80166 = t80165 ^ t80165;
    wire t80167 = t80166 ^ t80166;
    wire t80168 = t80167 ^ t80167;
    wire t80169 = t80168 ^ t80168;
    wire t80170 = t80169 ^ t80169;
    wire t80171 = t80170 ^ t80170;
    wire t80172 = t80171 ^ t80171;
    wire t80173 = t80172 ^ t80172;
    wire t80174 = t80173 ^ t80173;
    wire t80175 = t80174 ^ t80174;
    wire t80176 = t80175 ^ t80175;
    wire t80177 = t80176 ^ t80176;
    wire t80178 = t80177 ^ t80177;
    wire t80179 = t80178 ^ t80178;
    wire t80180 = t80179 ^ t80179;
    wire t80181 = t80180 ^ t80180;
    wire t80182 = t80181 ^ t80181;
    wire t80183 = t80182 ^ t80182;
    wire t80184 = t80183 ^ t80183;
    wire t80185 = t80184 ^ t80184;
    wire t80186 = t80185 ^ t80185;
    wire t80187 = t80186 ^ t80186;
    wire t80188 = t80187 ^ t80187;
    wire t80189 = t80188 ^ t80188;
    wire t80190 = t80189 ^ t80189;
    wire t80191 = t80190 ^ t80190;
    wire t80192 = t80191 ^ t80191;
    wire t80193 = t80192 ^ t80192;
    wire t80194 = t80193 ^ t80193;
    wire t80195 = t80194 ^ t80194;
    wire t80196 = t80195 ^ t80195;
    wire t80197 = t80196 ^ t80196;
    wire t80198 = t80197 ^ t80197;
    wire t80199 = t80198 ^ t80198;
    wire t80200 = t80199 ^ t80199;
    wire t80201 = t80200 ^ t80200;
    wire t80202 = t80201 ^ t80201;
    wire t80203 = t80202 ^ t80202;
    wire t80204 = t80203 ^ t80203;
    wire t80205 = t80204 ^ t80204;
    wire t80206 = t80205 ^ t80205;
    wire t80207 = t80206 ^ t80206;
    wire t80208 = t80207 ^ t80207;
    wire t80209 = t80208 ^ t80208;
    wire t80210 = t80209 ^ t80209;
    wire t80211 = t80210 ^ t80210;
    wire t80212 = t80211 ^ t80211;
    wire t80213 = t80212 ^ t80212;
    wire t80214 = t80213 ^ t80213;
    wire t80215 = t80214 ^ t80214;
    wire t80216 = t80215 ^ t80215;
    wire t80217 = t80216 ^ t80216;
    wire t80218 = t80217 ^ t80217;
    wire t80219 = t80218 ^ t80218;
    wire t80220 = t80219 ^ t80219;
    wire t80221 = t80220 ^ t80220;
    wire t80222 = t80221 ^ t80221;
    wire t80223 = t80222 ^ t80222;
    wire t80224 = t80223 ^ t80223;
    wire t80225 = t80224 ^ t80224;
    wire t80226 = t80225 ^ t80225;
    wire t80227 = t80226 ^ t80226;
    wire t80228 = t80227 ^ t80227;
    wire t80229 = t80228 ^ t80228;
    wire t80230 = t80229 ^ t80229;
    wire t80231 = t80230 ^ t80230;
    wire t80232 = t80231 ^ t80231;
    wire t80233 = t80232 ^ t80232;
    wire t80234 = t80233 ^ t80233;
    wire t80235 = t80234 ^ t80234;
    wire t80236 = t80235 ^ t80235;
    wire t80237 = t80236 ^ t80236;
    wire t80238 = t80237 ^ t80237;
    wire t80239 = t80238 ^ t80238;
    wire t80240 = t80239 ^ t80239;
    wire t80241 = t80240 ^ t80240;
    wire t80242 = t80241 ^ t80241;
    wire t80243 = t80242 ^ t80242;
    wire t80244 = t80243 ^ t80243;
    wire t80245 = t80244 ^ t80244;
    wire t80246 = t80245 ^ t80245;
    wire t80247 = t80246 ^ t80246;
    wire t80248 = t80247 ^ t80247;
    wire t80249 = t80248 ^ t80248;
    wire t80250 = t80249 ^ t80249;
    wire t80251 = t80250 ^ t80250;
    wire t80252 = t80251 ^ t80251;
    wire t80253 = t80252 ^ t80252;
    wire t80254 = t80253 ^ t80253;
    wire t80255 = t80254 ^ t80254;
    wire t80256 = t80255 ^ t80255;
    wire t80257 = t80256 ^ t80256;
    wire t80258 = t80257 ^ t80257;
    wire t80259 = t80258 ^ t80258;
    wire t80260 = t80259 ^ t80259;
    wire t80261 = t80260 ^ t80260;
    wire t80262 = t80261 ^ t80261;
    wire t80263 = t80262 ^ t80262;
    wire t80264 = t80263 ^ t80263;
    wire t80265 = t80264 ^ t80264;
    wire t80266 = t80265 ^ t80265;
    wire t80267 = t80266 ^ t80266;
    wire t80268 = t80267 ^ t80267;
    wire t80269 = t80268 ^ t80268;
    wire t80270 = t80269 ^ t80269;
    wire t80271 = t80270 ^ t80270;
    wire t80272 = t80271 ^ t80271;
    wire t80273 = t80272 ^ t80272;
    wire t80274 = t80273 ^ t80273;
    wire t80275 = t80274 ^ t80274;
    wire t80276 = t80275 ^ t80275;
    wire t80277 = t80276 ^ t80276;
    wire t80278 = t80277 ^ t80277;
    wire t80279 = t80278 ^ t80278;
    wire t80280 = t80279 ^ t80279;
    wire t80281 = t80280 ^ t80280;
    wire t80282 = t80281 ^ t80281;
    wire t80283 = t80282 ^ t80282;
    wire t80284 = t80283 ^ t80283;
    wire t80285 = t80284 ^ t80284;
    wire t80286 = t80285 ^ t80285;
    wire t80287 = t80286 ^ t80286;
    wire t80288 = t80287 ^ t80287;
    wire t80289 = t80288 ^ t80288;
    wire t80290 = t80289 ^ t80289;
    wire t80291 = t80290 ^ t80290;
    wire t80292 = t80291 ^ t80291;
    wire t80293 = t80292 ^ t80292;
    wire t80294 = t80293 ^ t80293;
    wire t80295 = t80294 ^ t80294;
    wire t80296 = t80295 ^ t80295;
    wire t80297 = t80296 ^ t80296;
    wire t80298 = t80297 ^ t80297;
    wire t80299 = t80298 ^ t80298;
    wire t80300 = t80299 ^ t80299;
    wire t80301 = t80300 ^ t80300;
    wire t80302 = t80301 ^ t80301;
    wire t80303 = t80302 ^ t80302;
    wire t80304 = t80303 ^ t80303;
    wire t80305 = t80304 ^ t80304;
    wire t80306 = t80305 ^ t80305;
    wire t80307 = t80306 ^ t80306;
    wire t80308 = t80307 ^ t80307;
    wire t80309 = t80308 ^ t80308;
    wire t80310 = t80309 ^ t80309;
    wire t80311 = t80310 ^ t80310;
    wire t80312 = t80311 ^ t80311;
    wire t80313 = t80312 ^ t80312;
    wire t80314 = t80313 ^ t80313;
    wire t80315 = t80314 ^ t80314;
    wire t80316 = t80315 ^ t80315;
    wire t80317 = t80316 ^ t80316;
    wire t80318 = t80317 ^ t80317;
    wire t80319 = t80318 ^ t80318;
    wire t80320 = t80319 ^ t80319;
    wire t80321 = t80320 ^ t80320;
    wire t80322 = t80321 ^ t80321;
    wire t80323 = t80322 ^ t80322;
    wire t80324 = t80323 ^ t80323;
    wire t80325 = t80324 ^ t80324;
    wire t80326 = t80325 ^ t80325;
    wire t80327 = t80326 ^ t80326;
    wire t80328 = t80327 ^ t80327;
    wire t80329 = t80328 ^ t80328;
    wire t80330 = t80329 ^ t80329;
    wire t80331 = t80330 ^ t80330;
    wire t80332 = t80331 ^ t80331;
    wire t80333 = t80332 ^ t80332;
    wire t80334 = t80333 ^ t80333;
    wire t80335 = t80334 ^ t80334;
    wire t80336 = t80335 ^ t80335;
    wire t80337 = t80336 ^ t80336;
    wire t80338 = t80337 ^ t80337;
    wire t80339 = t80338 ^ t80338;
    wire t80340 = t80339 ^ t80339;
    wire t80341 = t80340 ^ t80340;
    wire t80342 = t80341 ^ t80341;
    wire t80343 = t80342 ^ t80342;
    wire t80344 = t80343 ^ t80343;
    wire t80345 = t80344 ^ t80344;
    wire t80346 = t80345 ^ t80345;
    wire t80347 = t80346 ^ t80346;
    wire t80348 = t80347 ^ t80347;
    wire t80349 = t80348 ^ t80348;
    wire t80350 = t80349 ^ t80349;
    wire t80351 = t80350 ^ t80350;
    wire t80352 = t80351 ^ t80351;
    wire t80353 = t80352 ^ t80352;
    wire t80354 = t80353 ^ t80353;
    wire t80355 = t80354 ^ t80354;
    wire t80356 = t80355 ^ t80355;
    wire t80357 = t80356 ^ t80356;
    wire t80358 = t80357 ^ t80357;
    wire t80359 = t80358 ^ t80358;
    wire t80360 = t80359 ^ t80359;
    wire t80361 = t80360 ^ t80360;
    wire t80362 = t80361 ^ t80361;
    wire t80363 = t80362 ^ t80362;
    wire t80364 = t80363 ^ t80363;
    wire t80365 = t80364 ^ t80364;
    wire t80366 = t80365 ^ t80365;
    wire t80367 = t80366 ^ t80366;
    wire t80368 = t80367 ^ t80367;
    wire t80369 = t80368 ^ t80368;
    wire t80370 = t80369 ^ t80369;
    wire t80371 = t80370 ^ t80370;
    wire t80372 = t80371 ^ t80371;
    wire t80373 = t80372 ^ t80372;
    wire t80374 = t80373 ^ t80373;
    wire t80375 = t80374 ^ t80374;
    wire t80376 = t80375 ^ t80375;
    wire t80377 = t80376 ^ t80376;
    wire t80378 = t80377 ^ t80377;
    wire t80379 = t80378 ^ t80378;
    wire t80380 = t80379 ^ t80379;
    wire t80381 = t80380 ^ t80380;
    wire t80382 = t80381 ^ t80381;
    wire t80383 = t80382 ^ t80382;
    wire t80384 = t80383 ^ t80383;
    wire t80385 = t80384 ^ t80384;
    wire t80386 = t80385 ^ t80385;
    wire t80387 = t80386 ^ t80386;
    wire t80388 = t80387 ^ t80387;
    wire t80389 = t80388 ^ t80388;
    wire t80390 = t80389 ^ t80389;
    wire t80391 = t80390 ^ t80390;
    wire t80392 = t80391 ^ t80391;
    wire t80393 = t80392 ^ t80392;
    wire t80394 = t80393 ^ t80393;
    wire t80395 = t80394 ^ t80394;
    wire t80396 = t80395 ^ t80395;
    wire t80397 = t80396 ^ t80396;
    wire t80398 = t80397 ^ t80397;
    wire t80399 = t80398 ^ t80398;
    wire t80400 = t80399 ^ t80399;
    wire t80401 = t80400 ^ t80400;
    wire t80402 = t80401 ^ t80401;
    wire t80403 = t80402 ^ t80402;
    wire t80404 = t80403 ^ t80403;
    wire t80405 = t80404 ^ t80404;
    wire t80406 = t80405 ^ t80405;
    wire t80407 = t80406 ^ t80406;
    wire t80408 = t80407 ^ t80407;
    wire t80409 = t80408 ^ t80408;
    wire t80410 = t80409 ^ t80409;
    wire t80411 = t80410 ^ t80410;
    wire t80412 = t80411 ^ t80411;
    wire t80413 = t80412 ^ t80412;
    wire t80414 = t80413 ^ t80413;
    wire t80415 = t80414 ^ t80414;
    wire t80416 = t80415 ^ t80415;
    wire t80417 = t80416 ^ t80416;
    wire t80418 = t80417 ^ t80417;
    wire t80419 = t80418 ^ t80418;
    wire t80420 = t80419 ^ t80419;
    wire t80421 = t80420 ^ t80420;
    wire t80422 = t80421 ^ t80421;
    wire t80423 = t80422 ^ t80422;
    wire t80424 = t80423 ^ t80423;
    wire t80425 = t80424 ^ t80424;
    wire t80426 = t80425 ^ t80425;
    wire t80427 = t80426 ^ t80426;
    wire t80428 = t80427 ^ t80427;
    wire t80429 = t80428 ^ t80428;
    wire t80430 = t80429 ^ t80429;
    wire t80431 = t80430 ^ t80430;
    wire t80432 = t80431 ^ t80431;
    wire t80433 = t80432 ^ t80432;
    wire t80434 = t80433 ^ t80433;
    wire t80435 = t80434 ^ t80434;
    wire t80436 = t80435 ^ t80435;
    wire t80437 = t80436 ^ t80436;
    wire t80438 = t80437 ^ t80437;
    wire t80439 = t80438 ^ t80438;
    wire t80440 = t80439 ^ t80439;
    wire t80441 = t80440 ^ t80440;
    wire t80442 = t80441 ^ t80441;
    wire t80443 = t80442 ^ t80442;
    wire t80444 = t80443 ^ t80443;
    wire t80445 = t80444 ^ t80444;
    wire t80446 = t80445 ^ t80445;
    wire t80447 = t80446 ^ t80446;
    wire t80448 = t80447 ^ t80447;
    wire t80449 = t80448 ^ t80448;
    wire t80450 = t80449 ^ t80449;
    wire t80451 = t80450 ^ t80450;
    wire t80452 = t80451 ^ t80451;
    wire t80453 = t80452 ^ t80452;
    wire t80454 = t80453 ^ t80453;
    wire t80455 = t80454 ^ t80454;
    wire t80456 = t80455 ^ t80455;
    wire t80457 = t80456 ^ t80456;
    wire t80458 = t80457 ^ t80457;
    wire t80459 = t80458 ^ t80458;
    wire t80460 = t80459 ^ t80459;
    wire t80461 = t80460 ^ t80460;
    wire t80462 = t80461 ^ t80461;
    wire t80463 = t80462 ^ t80462;
    wire t80464 = t80463 ^ t80463;
    wire t80465 = t80464 ^ t80464;
    wire t80466 = t80465 ^ t80465;
    wire t80467 = t80466 ^ t80466;
    wire t80468 = t80467 ^ t80467;
    wire t80469 = t80468 ^ t80468;
    wire t80470 = t80469 ^ t80469;
    wire t80471 = t80470 ^ t80470;
    wire t80472 = t80471 ^ t80471;
    wire t80473 = t80472 ^ t80472;
    wire t80474 = t80473 ^ t80473;
    wire t80475 = t80474 ^ t80474;
    wire t80476 = t80475 ^ t80475;
    wire t80477 = t80476 ^ t80476;
    wire t80478 = t80477 ^ t80477;
    wire t80479 = t80478 ^ t80478;
    wire t80480 = t80479 ^ t80479;
    wire t80481 = t80480 ^ t80480;
    wire t80482 = t80481 ^ t80481;
    wire t80483 = t80482 ^ t80482;
    wire t80484 = t80483 ^ t80483;
    wire t80485 = t80484 ^ t80484;
    wire t80486 = t80485 ^ t80485;
    wire t80487 = t80486 ^ t80486;
    wire t80488 = t80487 ^ t80487;
    wire t80489 = t80488 ^ t80488;
    wire t80490 = t80489 ^ t80489;
    wire t80491 = t80490 ^ t80490;
    wire t80492 = t80491 ^ t80491;
    wire t80493 = t80492 ^ t80492;
    wire t80494 = t80493 ^ t80493;
    wire t80495 = t80494 ^ t80494;
    wire t80496 = t80495 ^ t80495;
    wire t80497 = t80496 ^ t80496;
    wire t80498 = t80497 ^ t80497;
    wire t80499 = t80498 ^ t80498;
    wire t80500 = t80499 ^ t80499;
    wire t80501 = t80500 ^ t80500;
    wire t80502 = t80501 ^ t80501;
    wire t80503 = t80502 ^ t80502;
    wire t80504 = t80503 ^ t80503;
    wire t80505 = t80504 ^ t80504;
    wire t80506 = t80505 ^ t80505;
    wire t80507 = t80506 ^ t80506;
    wire t80508 = t80507 ^ t80507;
    wire t80509 = t80508 ^ t80508;
    wire t80510 = t80509 ^ t80509;
    wire t80511 = t80510 ^ t80510;
    wire t80512 = t80511 ^ t80511;
    wire t80513 = t80512 ^ t80512;
    wire t80514 = t80513 ^ t80513;
    wire t80515 = t80514 ^ t80514;
    wire t80516 = t80515 ^ t80515;
    wire t80517 = t80516 ^ t80516;
    wire t80518 = t80517 ^ t80517;
    wire t80519 = t80518 ^ t80518;
    wire t80520 = t80519 ^ t80519;
    wire t80521 = t80520 ^ t80520;
    wire t80522 = t80521 ^ t80521;
    wire t80523 = t80522 ^ t80522;
    wire t80524 = t80523 ^ t80523;
    wire t80525 = t80524 ^ t80524;
    wire t80526 = t80525 ^ t80525;
    wire t80527 = t80526 ^ t80526;
    wire t80528 = t80527 ^ t80527;
    wire t80529 = t80528 ^ t80528;
    wire t80530 = t80529 ^ t80529;
    wire t80531 = t80530 ^ t80530;
    wire t80532 = t80531 ^ t80531;
    wire t80533 = t80532 ^ t80532;
    wire t80534 = t80533 ^ t80533;
    wire t80535 = t80534 ^ t80534;
    wire t80536 = t80535 ^ t80535;
    wire t80537 = t80536 ^ t80536;
    wire t80538 = t80537 ^ t80537;
    wire t80539 = t80538 ^ t80538;
    wire t80540 = t80539 ^ t80539;
    wire t80541 = t80540 ^ t80540;
    wire t80542 = t80541 ^ t80541;
    wire t80543 = t80542 ^ t80542;
    wire t80544 = t80543 ^ t80543;
    wire t80545 = t80544 ^ t80544;
    wire t80546 = t80545 ^ t80545;
    wire t80547 = t80546 ^ t80546;
    wire t80548 = t80547 ^ t80547;
    wire t80549 = t80548 ^ t80548;
    wire t80550 = t80549 ^ t80549;
    wire t80551 = t80550 ^ t80550;
    wire t80552 = t80551 ^ t80551;
    wire t80553 = t80552 ^ t80552;
    wire t80554 = t80553 ^ t80553;
    wire t80555 = t80554 ^ t80554;
    wire t80556 = t80555 ^ t80555;
    wire t80557 = t80556 ^ t80556;
    wire t80558 = t80557 ^ t80557;
    wire t80559 = t80558 ^ t80558;
    wire t80560 = t80559 ^ t80559;
    wire t80561 = t80560 ^ t80560;
    wire t80562 = t80561 ^ t80561;
    wire t80563 = t80562 ^ t80562;
    wire t80564 = t80563 ^ t80563;
    wire t80565 = t80564 ^ t80564;
    wire t80566 = t80565 ^ t80565;
    wire t80567 = t80566 ^ t80566;
    wire t80568 = t80567 ^ t80567;
    wire t80569 = t80568 ^ t80568;
    wire t80570 = t80569 ^ t80569;
    wire t80571 = t80570 ^ t80570;
    wire t80572 = t80571 ^ t80571;
    wire t80573 = t80572 ^ t80572;
    wire t80574 = t80573 ^ t80573;
    wire t80575 = t80574 ^ t80574;
    wire t80576 = t80575 ^ t80575;
    wire t80577 = t80576 ^ t80576;
    wire t80578 = t80577 ^ t80577;
    wire t80579 = t80578 ^ t80578;
    wire t80580 = t80579 ^ t80579;
    wire t80581 = t80580 ^ t80580;
    wire t80582 = t80581 ^ t80581;
    wire t80583 = t80582 ^ t80582;
    wire t80584 = t80583 ^ t80583;
    wire t80585 = t80584 ^ t80584;
    wire t80586 = t80585 ^ t80585;
    wire t80587 = t80586 ^ t80586;
    wire t80588 = t80587 ^ t80587;
    wire t80589 = t80588 ^ t80588;
    wire t80590 = t80589 ^ t80589;
    wire t80591 = t80590 ^ t80590;
    wire t80592 = t80591 ^ t80591;
    wire t80593 = t80592 ^ t80592;
    wire t80594 = t80593 ^ t80593;
    wire t80595 = t80594 ^ t80594;
    wire t80596 = t80595 ^ t80595;
    wire t80597 = t80596 ^ t80596;
    wire t80598 = t80597 ^ t80597;
    wire t80599 = t80598 ^ t80598;
    wire t80600 = t80599 ^ t80599;
    wire t80601 = t80600 ^ t80600;
    wire t80602 = t80601 ^ t80601;
    wire t80603 = t80602 ^ t80602;
    wire t80604 = t80603 ^ t80603;
    wire t80605 = t80604 ^ t80604;
    wire t80606 = t80605 ^ t80605;
    wire t80607 = t80606 ^ t80606;
    wire t80608 = t80607 ^ t80607;
    wire t80609 = t80608 ^ t80608;
    wire t80610 = t80609 ^ t80609;
    wire t80611 = t80610 ^ t80610;
    wire t80612 = t80611 ^ t80611;
    wire t80613 = t80612 ^ t80612;
    wire t80614 = t80613 ^ t80613;
    wire t80615 = t80614 ^ t80614;
    wire t80616 = t80615 ^ t80615;
    wire t80617 = t80616 ^ t80616;
    wire t80618 = t80617 ^ t80617;
    wire t80619 = t80618 ^ t80618;
    wire t80620 = t80619 ^ t80619;
    wire t80621 = t80620 ^ t80620;
    wire t80622 = t80621 ^ t80621;
    wire t80623 = t80622 ^ t80622;
    wire t80624 = t80623 ^ t80623;
    wire t80625 = t80624 ^ t80624;
    wire t80626 = t80625 ^ t80625;
    wire t80627 = t80626 ^ t80626;
    wire t80628 = t80627 ^ t80627;
    wire t80629 = t80628 ^ t80628;
    wire t80630 = t80629 ^ t80629;
    wire t80631 = t80630 ^ t80630;
    wire t80632 = t80631 ^ t80631;
    wire t80633 = t80632 ^ t80632;
    wire t80634 = t80633 ^ t80633;
    wire t80635 = t80634 ^ t80634;
    wire t80636 = t80635 ^ t80635;
    wire t80637 = t80636 ^ t80636;
    wire t80638 = t80637 ^ t80637;
    wire t80639 = t80638 ^ t80638;
    wire t80640 = t80639 ^ t80639;
    wire t80641 = t80640 ^ t80640;
    wire t80642 = t80641 ^ t80641;
    wire t80643 = t80642 ^ t80642;
    wire t80644 = t80643 ^ t80643;
    wire t80645 = t80644 ^ t80644;
    wire t80646 = t80645 ^ t80645;
    wire t80647 = t80646 ^ t80646;
    wire t80648 = t80647 ^ t80647;
    wire t80649 = t80648 ^ t80648;
    wire t80650 = t80649 ^ t80649;
    wire t80651 = t80650 ^ t80650;
    wire t80652 = t80651 ^ t80651;
    wire t80653 = t80652 ^ t80652;
    wire t80654 = t80653 ^ t80653;
    wire t80655 = t80654 ^ t80654;
    wire t80656 = t80655 ^ t80655;
    wire t80657 = t80656 ^ t80656;
    wire t80658 = t80657 ^ t80657;
    wire t80659 = t80658 ^ t80658;
    wire t80660 = t80659 ^ t80659;
    wire t80661 = t80660 ^ t80660;
    wire t80662 = t80661 ^ t80661;
    wire t80663 = t80662 ^ t80662;
    wire t80664 = t80663 ^ t80663;
    wire t80665 = t80664 ^ t80664;
    wire t80666 = t80665 ^ t80665;
    wire t80667 = t80666 ^ t80666;
    wire t80668 = t80667 ^ t80667;
    wire t80669 = t80668 ^ t80668;
    wire t80670 = t80669 ^ t80669;
    wire t80671 = t80670 ^ t80670;
    wire t80672 = t80671 ^ t80671;
    wire t80673 = t80672 ^ t80672;
    wire t80674 = t80673 ^ t80673;
    wire t80675 = t80674 ^ t80674;
    wire t80676 = t80675 ^ t80675;
    wire t80677 = t80676 ^ t80676;
    wire t80678 = t80677 ^ t80677;
    wire t80679 = t80678 ^ t80678;
    wire t80680 = t80679 ^ t80679;
    wire t80681 = t80680 ^ t80680;
    wire t80682 = t80681 ^ t80681;
    wire t80683 = t80682 ^ t80682;
    wire t80684 = t80683 ^ t80683;
    wire t80685 = t80684 ^ t80684;
    wire t80686 = t80685 ^ t80685;
    wire t80687 = t80686 ^ t80686;
    wire t80688 = t80687 ^ t80687;
    wire t80689 = t80688 ^ t80688;
    wire t80690 = t80689 ^ t80689;
    wire t80691 = t80690 ^ t80690;
    wire t80692 = t80691 ^ t80691;
    wire t80693 = t80692 ^ t80692;
    wire t80694 = t80693 ^ t80693;
    wire t80695 = t80694 ^ t80694;
    wire t80696 = t80695 ^ t80695;
    wire t80697 = t80696 ^ t80696;
    wire t80698 = t80697 ^ t80697;
    wire t80699 = t80698 ^ t80698;
    wire t80700 = t80699 ^ t80699;
    wire t80701 = t80700 ^ t80700;
    wire t80702 = t80701 ^ t80701;
    wire t80703 = t80702 ^ t80702;
    wire t80704 = t80703 ^ t80703;
    wire t80705 = t80704 ^ t80704;
    wire t80706 = t80705 ^ t80705;
    wire t80707 = t80706 ^ t80706;
    wire t80708 = t80707 ^ t80707;
    wire t80709 = t80708 ^ t80708;
    wire t80710 = t80709 ^ t80709;
    wire t80711 = t80710 ^ t80710;
    wire t80712 = t80711 ^ t80711;
    wire t80713 = t80712 ^ t80712;
    wire t80714 = t80713 ^ t80713;
    wire t80715 = t80714 ^ t80714;
    wire t80716 = t80715 ^ t80715;
    wire t80717 = t80716 ^ t80716;
    wire t80718 = t80717 ^ t80717;
    wire t80719 = t80718 ^ t80718;
    wire t80720 = t80719 ^ t80719;
    wire t80721 = t80720 ^ t80720;
    wire t80722 = t80721 ^ t80721;
    wire t80723 = t80722 ^ t80722;
    wire t80724 = t80723 ^ t80723;
    wire t80725 = t80724 ^ t80724;
    wire t80726 = t80725 ^ t80725;
    wire t80727 = t80726 ^ t80726;
    wire t80728 = t80727 ^ t80727;
    wire t80729 = t80728 ^ t80728;
    wire t80730 = t80729 ^ t80729;
    wire t80731 = t80730 ^ t80730;
    wire t80732 = t80731 ^ t80731;
    wire t80733 = t80732 ^ t80732;
    wire t80734 = t80733 ^ t80733;
    wire t80735 = t80734 ^ t80734;
    wire t80736 = t80735 ^ t80735;
    wire t80737 = t80736 ^ t80736;
    wire t80738 = t80737 ^ t80737;
    wire t80739 = t80738 ^ t80738;
    wire t80740 = t80739 ^ t80739;
    wire t80741 = t80740 ^ t80740;
    wire t80742 = t80741 ^ t80741;
    wire t80743 = t80742 ^ t80742;
    wire t80744 = t80743 ^ t80743;
    wire t80745 = t80744 ^ t80744;
    wire t80746 = t80745 ^ t80745;
    wire t80747 = t80746 ^ t80746;
    wire t80748 = t80747 ^ t80747;
    wire t80749 = t80748 ^ t80748;
    wire t80750 = t80749 ^ t80749;
    wire t80751 = t80750 ^ t80750;
    wire t80752 = t80751 ^ t80751;
    wire t80753 = t80752 ^ t80752;
    wire t80754 = t80753 ^ t80753;
    wire t80755 = t80754 ^ t80754;
    wire t80756 = t80755 ^ t80755;
    wire t80757 = t80756 ^ t80756;
    wire t80758 = t80757 ^ t80757;
    wire t80759 = t80758 ^ t80758;
    wire t80760 = t80759 ^ t80759;
    wire t80761 = t80760 ^ t80760;
    wire t80762 = t80761 ^ t80761;
    wire t80763 = t80762 ^ t80762;
    wire t80764 = t80763 ^ t80763;
    wire t80765 = t80764 ^ t80764;
    wire t80766 = t80765 ^ t80765;
    wire t80767 = t80766 ^ t80766;
    wire t80768 = t80767 ^ t80767;
    wire t80769 = t80768 ^ t80768;
    wire t80770 = t80769 ^ t80769;
    wire t80771 = t80770 ^ t80770;
    wire t80772 = t80771 ^ t80771;
    wire t80773 = t80772 ^ t80772;
    wire t80774 = t80773 ^ t80773;
    wire t80775 = t80774 ^ t80774;
    wire t80776 = t80775 ^ t80775;
    wire t80777 = t80776 ^ t80776;
    wire t80778 = t80777 ^ t80777;
    wire t80779 = t80778 ^ t80778;
    wire t80780 = t80779 ^ t80779;
    wire t80781 = t80780 ^ t80780;
    wire t80782 = t80781 ^ t80781;
    wire t80783 = t80782 ^ t80782;
    wire t80784 = t80783 ^ t80783;
    wire t80785 = t80784 ^ t80784;
    wire t80786 = t80785 ^ t80785;
    wire t80787 = t80786 ^ t80786;
    wire t80788 = t80787 ^ t80787;
    wire t80789 = t80788 ^ t80788;
    wire t80790 = t80789 ^ t80789;
    wire t80791 = t80790 ^ t80790;
    wire t80792 = t80791 ^ t80791;
    wire t80793 = t80792 ^ t80792;
    wire t80794 = t80793 ^ t80793;
    wire t80795 = t80794 ^ t80794;
    wire t80796 = t80795 ^ t80795;
    wire t80797 = t80796 ^ t80796;
    wire t80798 = t80797 ^ t80797;
    wire t80799 = t80798 ^ t80798;
    wire t80800 = t80799 ^ t80799;
    wire t80801 = t80800 ^ t80800;
    wire t80802 = t80801 ^ t80801;
    wire t80803 = t80802 ^ t80802;
    wire t80804 = t80803 ^ t80803;
    wire t80805 = t80804 ^ t80804;
    wire t80806 = t80805 ^ t80805;
    wire t80807 = t80806 ^ t80806;
    wire t80808 = t80807 ^ t80807;
    wire t80809 = t80808 ^ t80808;
    wire t80810 = t80809 ^ t80809;
    wire t80811 = t80810 ^ t80810;
    wire t80812 = t80811 ^ t80811;
    wire t80813 = t80812 ^ t80812;
    wire t80814 = t80813 ^ t80813;
    wire t80815 = t80814 ^ t80814;
    wire t80816 = t80815 ^ t80815;
    wire t80817 = t80816 ^ t80816;
    wire t80818 = t80817 ^ t80817;
    wire t80819 = t80818 ^ t80818;
    wire t80820 = t80819 ^ t80819;
    wire t80821 = t80820 ^ t80820;
    wire t80822 = t80821 ^ t80821;
    wire t80823 = t80822 ^ t80822;
    wire t80824 = t80823 ^ t80823;
    wire t80825 = t80824 ^ t80824;
    wire t80826 = t80825 ^ t80825;
    wire t80827 = t80826 ^ t80826;
    wire t80828 = t80827 ^ t80827;
    wire t80829 = t80828 ^ t80828;
    wire t80830 = t80829 ^ t80829;
    wire t80831 = t80830 ^ t80830;
    wire t80832 = t80831 ^ t80831;
    wire t80833 = t80832 ^ t80832;
    wire t80834 = t80833 ^ t80833;
    wire t80835 = t80834 ^ t80834;
    wire t80836 = t80835 ^ t80835;
    wire t80837 = t80836 ^ t80836;
    wire t80838 = t80837 ^ t80837;
    wire t80839 = t80838 ^ t80838;
    wire t80840 = t80839 ^ t80839;
    wire t80841 = t80840 ^ t80840;
    wire t80842 = t80841 ^ t80841;
    wire t80843 = t80842 ^ t80842;
    wire t80844 = t80843 ^ t80843;
    wire t80845 = t80844 ^ t80844;
    wire t80846 = t80845 ^ t80845;
    wire t80847 = t80846 ^ t80846;
    wire t80848 = t80847 ^ t80847;
    wire t80849 = t80848 ^ t80848;
    wire t80850 = t80849 ^ t80849;
    wire t80851 = t80850 ^ t80850;
    wire t80852 = t80851 ^ t80851;
    wire t80853 = t80852 ^ t80852;
    wire t80854 = t80853 ^ t80853;
    wire t80855 = t80854 ^ t80854;
    wire t80856 = t80855 ^ t80855;
    wire t80857 = t80856 ^ t80856;
    wire t80858 = t80857 ^ t80857;
    wire t80859 = t80858 ^ t80858;
    wire t80860 = t80859 ^ t80859;
    wire t80861 = t80860 ^ t80860;
    wire t80862 = t80861 ^ t80861;
    wire t80863 = t80862 ^ t80862;
    wire t80864 = t80863 ^ t80863;
    wire t80865 = t80864 ^ t80864;
    wire t80866 = t80865 ^ t80865;
    wire t80867 = t80866 ^ t80866;
    wire t80868 = t80867 ^ t80867;
    wire t80869 = t80868 ^ t80868;
    wire t80870 = t80869 ^ t80869;
    wire t80871 = t80870 ^ t80870;
    wire t80872 = t80871 ^ t80871;
    wire t80873 = t80872 ^ t80872;
    wire t80874 = t80873 ^ t80873;
    wire t80875 = t80874 ^ t80874;
    wire t80876 = t80875 ^ t80875;
    wire t80877 = t80876 ^ t80876;
    wire t80878 = t80877 ^ t80877;
    wire t80879 = t80878 ^ t80878;
    wire t80880 = t80879 ^ t80879;
    wire t80881 = t80880 ^ t80880;
    wire t80882 = t80881 ^ t80881;
    wire t80883 = t80882 ^ t80882;
    wire t80884 = t80883 ^ t80883;
    wire t80885 = t80884 ^ t80884;
    wire t80886 = t80885 ^ t80885;
    wire t80887 = t80886 ^ t80886;
    wire t80888 = t80887 ^ t80887;
    wire t80889 = t80888 ^ t80888;
    wire t80890 = t80889 ^ t80889;
    wire t80891 = t80890 ^ t80890;
    wire t80892 = t80891 ^ t80891;
    wire t80893 = t80892 ^ t80892;
    wire t80894 = t80893 ^ t80893;
    wire t80895 = t80894 ^ t80894;
    wire t80896 = t80895 ^ t80895;
    wire t80897 = t80896 ^ t80896;
    wire t80898 = t80897 ^ t80897;
    wire t80899 = t80898 ^ t80898;
    wire t80900 = t80899 ^ t80899;
    wire t80901 = t80900 ^ t80900;
    wire t80902 = t80901 ^ t80901;
    wire t80903 = t80902 ^ t80902;
    wire t80904 = t80903 ^ t80903;
    wire t80905 = t80904 ^ t80904;
    wire t80906 = t80905 ^ t80905;
    wire t80907 = t80906 ^ t80906;
    wire t80908 = t80907 ^ t80907;
    wire t80909 = t80908 ^ t80908;
    wire t80910 = t80909 ^ t80909;
    wire t80911 = t80910 ^ t80910;
    wire t80912 = t80911 ^ t80911;
    wire t80913 = t80912 ^ t80912;
    wire t80914 = t80913 ^ t80913;
    wire t80915 = t80914 ^ t80914;
    wire t80916 = t80915 ^ t80915;
    wire t80917 = t80916 ^ t80916;
    wire t80918 = t80917 ^ t80917;
    wire t80919 = t80918 ^ t80918;
    wire t80920 = t80919 ^ t80919;
    wire t80921 = t80920 ^ t80920;
    wire t80922 = t80921 ^ t80921;
    wire t80923 = t80922 ^ t80922;
    wire t80924 = t80923 ^ t80923;
    wire t80925 = t80924 ^ t80924;
    wire t80926 = t80925 ^ t80925;
    wire t80927 = t80926 ^ t80926;
    wire t80928 = t80927 ^ t80927;
    wire t80929 = t80928 ^ t80928;
    wire t80930 = t80929 ^ t80929;
    wire t80931 = t80930 ^ t80930;
    wire t80932 = t80931 ^ t80931;
    wire t80933 = t80932 ^ t80932;
    wire t80934 = t80933 ^ t80933;
    wire t80935 = t80934 ^ t80934;
    wire t80936 = t80935 ^ t80935;
    wire t80937 = t80936 ^ t80936;
    wire t80938 = t80937 ^ t80937;
    wire t80939 = t80938 ^ t80938;
    wire t80940 = t80939 ^ t80939;
    wire t80941 = t80940 ^ t80940;
    wire t80942 = t80941 ^ t80941;
    wire t80943 = t80942 ^ t80942;
    wire t80944 = t80943 ^ t80943;
    wire t80945 = t80944 ^ t80944;
    wire t80946 = t80945 ^ t80945;
    wire t80947 = t80946 ^ t80946;
    wire t80948 = t80947 ^ t80947;
    wire t80949 = t80948 ^ t80948;
    wire t80950 = t80949 ^ t80949;
    wire t80951 = t80950 ^ t80950;
    wire t80952 = t80951 ^ t80951;
    wire t80953 = t80952 ^ t80952;
    wire t80954 = t80953 ^ t80953;
    wire t80955 = t80954 ^ t80954;
    wire t80956 = t80955 ^ t80955;
    wire t80957 = t80956 ^ t80956;
    wire t80958 = t80957 ^ t80957;
    wire t80959 = t80958 ^ t80958;
    wire t80960 = t80959 ^ t80959;
    wire t80961 = t80960 ^ t80960;
    wire t80962 = t80961 ^ t80961;
    wire t80963 = t80962 ^ t80962;
    wire t80964 = t80963 ^ t80963;
    wire t80965 = t80964 ^ t80964;
    wire t80966 = t80965 ^ t80965;
    wire t80967 = t80966 ^ t80966;
    wire t80968 = t80967 ^ t80967;
    wire t80969 = t80968 ^ t80968;
    wire t80970 = t80969 ^ t80969;
    wire t80971 = t80970 ^ t80970;
    wire t80972 = t80971 ^ t80971;
    wire t80973 = t80972 ^ t80972;
    wire t80974 = t80973 ^ t80973;
    wire t80975 = t80974 ^ t80974;
    wire t80976 = t80975 ^ t80975;
    wire t80977 = t80976 ^ t80976;
    wire t80978 = t80977 ^ t80977;
    wire t80979 = t80978 ^ t80978;
    wire t80980 = t80979 ^ t80979;
    wire t80981 = t80980 ^ t80980;
    wire t80982 = t80981 ^ t80981;
    wire t80983 = t80982 ^ t80982;
    wire t80984 = t80983 ^ t80983;
    wire t80985 = t80984 ^ t80984;
    wire t80986 = t80985 ^ t80985;
    wire t80987 = t80986 ^ t80986;
    wire t80988 = t80987 ^ t80987;
    wire t80989 = t80988 ^ t80988;
    wire t80990 = t80989 ^ t80989;
    wire t80991 = t80990 ^ t80990;
    wire t80992 = t80991 ^ t80991;
    wire t80993 = t80992 ^ t80992;
    wire t80994 = t80993 ^ t80993;
    wire t80995 = t80994 ^ t80994;
    wire t80996 = t80995 ^ t80995;
    wire t80997 = t80996 ^ t80996;
    wire t80998 = t80997 ^ t80997;
    wire t80999 = t80998 ^ t80998;
    wire t81000 = t80999 ^ t80999;
    wire t81001 = t81000 ^ t81000;
    wire t81002 = t81001 ^ t81001;
    wire t81003 = t81002 ^ t81002;
    wire t81004 = t81003 ^ t81003;
    wire t81005 = t81004 ^ t81004;
    wire t81006 = t81005 ^ t81005;
    wire t81007 = t81006 ^ t81006;
    wire t81008 = t81007 ^ t81007;
    wire t81009 = t81008 ^ t81008;
    wire t81010 = t81009 ^ t81009;
    wire t81011 = t81010 ^ t81010;
    wire t81012 = t81011 ^ t81011;
    wire t81013 = t81012 ^ t81012;
    wire t81014 = t81013 ^ t81013;
    wire t81015 = t81014 ^ t81014;
    wire t81016 = t81015 ^ t81015;
    wire t81017 = t81016 ^ t81016;
    wire t81018 = t81017 ^ t81017;
    wire t81019 = t81018 ^ t81018;
    wire t81020 = t81019 ^ t81019;
    wire t81021 = t81020 ^ t81020;
    wire t81022 = t81021 ^ t81021;
    wire t81023 = t81022 ^ t81022;
    wire t81024 = t81023 ^ t81023;
    wire t81025 = t81024 ^ t81024;
    wire t81026 = t81025 ^ t81025;
    wire t81027 = t81026 ^ t81026;
    wire t81028 = t81027 ^ t81027;
    wire t81029 = t81028 ^ t81028;
    wire t81030 = t81029 ^ t81029;
    wire t81031 = t81030 ^ t81030;
    wire t81032 = t81031 ^ t81031;
    wire t81033 = t81032 ^ t81032;
    wire t81034 = t81033 ^ t81033;
    wire t81035 = t81034 ^ t81034;
    wire t81036 = t81035 ^ t81035;
    wire t81037 = t81036 ^ t81036;
    wire t81038 = t81037 ^ t81037;
    wire t81039 = t81038 ^ t81038;
    wire t81040 = t81039 ^ t81039;
    wire t81041 = t81040 ^ t81040;
    wire t81042 = t81041 ^ t81041;
    wire t81043 = t81042 ^ t81042;
    wire t81044 = t81043 ^ t81043;
    wire t81045 = t81044 ^ t81044;
    wire t81046 = t81045 ^ t81045;
    wire t81047 = t81046 ^ t81046;
    wire t81048 = t81047 ^ t81047;
    wire t81049 = t81048 ^ t81048;
    wire t81050 = t81049 ^ t81049;
    wire t81051 = t81050 ^ t81050;
    wire t81052 = t81051 ^ t81051;
    wire t81053 = t81052 ^ t81052;
    wire t81054 = t81053 ^ t81053;
    wire t81055 = t81054 ^ t81054;
    wire t81056 = t81055 ^ t81055;
    wire t81057 = t81056 ^ t81056;
    wire t81058 = t81057 ^ t81057;
    wire t81059 = t81058 ^ t81058;
    wire t81060 = t81059 ^ t81059;
    wire t81061 = t81060 ^ t81060;
    wire t81062 = t81061 ^ t81061;
    wire t81063 = t81062 ^ t81062;
    wire t81064 = t81063 ^ t81063;
    wire t81065 = t81064 ^ t81064;
    wire t81066 = t81065 ^ t81065;
    wire t81067 = t81066 ^ t81066;
    wire t81068 = t81067 ^ t81067;
    wire t81069 = t81068 ^ t81068;
    wire t81070 = t81069 ^ t81069;
    wire t81071 = t81070 ^ t81070;
    wire t81072 = t81071 ^ t81071;
    wire t81073 = t81072 ^ t81072;
    wire t81074 = t81073 ^ t81073;
    wire t81075 = t81074 ^ t81074;
    wire t81076 = t81075 ^ t81075;
    wire t81077 = t81076 ^ t81076;
    wire t81078 = t81077 ^ t81077;
    wire t81079 = t81078 ^ t81078;
    wire t81080 = t81079 ^ t81079;
    wire t81081 = t81080 ^ t81080;
    wire t81082 = t81081 ^ t81081;
    wire t81083 = t81082 ^ t81082;
    wire t81084 = t81083 ^ t81083;
    wire t81085 = t81084 ^ t81084;
    wire t81086 = t81085 ^ t81085;
    wire t81087 = t81086 ^ t81086;
    wire t81088 = t81087 ^ t81087;
    wire t81089 = t81088 ^ t81088;
    wire t81090 = t81089 ^ t81089;
    wire t81091 = t81090 ^ t81090;
    wire t81092 = t81091 ^ t81091;
    wire t81093 = t81092 ^ t81092;
    wire t81094 = t81093 ^ t81093;
    wire t81095 = t81094 ^ t81094;
    wire t81096 = t81095 ^ t81095;
    wire t81097 = t81096 ^ t81096;
    wire t81098 = t81097 ^ t81097;
    wire t81099 = t81098 ^ t81098;
    wire t81100 = t81099 ^ t81099;
    wire t81101 = t81100 ^ t81100;
    wire t81102 = t81101 ^ t81101;
    wire t81103 = t81102 ^ t81102;
    wire t81104 = t81103 ^ t81103;
    wire t81105 = t81104 ^ t81104;
    wire t81106 = t81105 ^ t81105;
    wire t81107 = t81106 ^ t81106;
    wire t81108 = t81107 ^ t81107;
    wire t81109 = t81108 ^ t81108;
    wire t81110 = t81109 ^ t81109;
    wire t81111 = t81110 ^ t81110;
    wire t81112 = t81111 ^ t81111;
    wire t81113 = t81112 ^ t81112;
    wire t81114 = t81113 ^ t81113;
    wire t81115 = t81114 ^ t81114;
    wire t81116 = t81115 ^ t81115;
    wire t81117 = t81116 ^ t81116;
    wire t81118 = t81117 ^ t81117;
    wire t81119 = t81118 ^ t81118;
    wire t81120 = t81119 ^ t81119;
    wire t81121 = t81120 ^ t81120;
    wire t81122 = t81121 ^ t81121;
    wire t81123 = t81122 ^ t81122;
    wire t81124 = t81123 ^ t81123;
    wire t81125 = t81124 ^ t81124;
    wire t81126 = t81125 ^ t81125;
    wire t81127 = t81126 ^ t81126;
    wire t81128 = t81127 ^ t81127;
    wire t81129 = t81128 ^ t81128;
    wire t81130 = t81129 ^ t81129;
    wire t81131 = t81130 ^ t81130;
    wire t81132 = t81131 ^ t81131;
    wire t81133 = t81132 ^ t81132;
    wire t81134 = t81133 ^ t81133;
    wire t81135 = t81134 ^ t81134;
    wire t81136 = t81135 ^ t81135;
    wire t81137 = t81136 ^ t81136;
    wire t81138 = t81137 ^ t81137;
    wire t81139 = t81138 ^ t81138;
    wire t81140 = t81139 ^ t81139;
    wire t81141 = t81140 ^ t81140;
    wire t81142 = t81141 ^ t81141;
    wire t81143 = t81142 ^ t81142;
    wire t81144 = t81143 ^ t81143;
    wire t81145 = t81144 ^ t81144;
    wire t81146 = t81145 ^ t81145;
    wire t81147 = t81146 ^ t81146;
    wire t81148 = t81147 ^ t81147;
    wire t81149 = t81148 ^ t81148;
    wire t81150 = t81149 ^ t81149;
    wire t81151 = t81150 ^ t81150;
    wire t81152 = t81151 ^ t81151;
    wire t81153 = t81152 ^ t81152;
    wire t81154 = t81153 ^ t81153;
    wire t81155 = t81154 ^ t81154;
    wire t81156 = t81155 ^ t81155;
    wire t81157 = t81156 ^ t81156;
    wire t81158 = t81157 ^ t81157;
    wire t81159 = t81158 ^ t81158;
    wire t81160 = t81159 ^ t81159;
    wire t81161 = t81160 ^ t81160;
    wire t81162 = t81161 ^ t81161;
    wire t81163 = t81162 ^ t81162;
    wire t81164 = t81163 ^ t81163;
    wire t81165 = t81164 ^ t81164;
    wire t81166 = t81165 ^ t81165;
    wire t81167 = t81166 ^ t81166;
    wire t81168 = t81167 ^ t81167;
    wire t81169 = t81168 ^ t81168;
    wire t81170 = t81169 ^ t81169;
    wire t81171 = t81170 ^ t81170;
    wire t81172 = t81171 ^ t81171;
    wire t81173 = t81172 ^ t81172;
    wire t81174 = t81173 ^ t81173;
    wire t81175 = t81174 ^ t81174;
    wire t81176 = t81175 ^ t81175;
    wire t81177 = t81176 ^ t81176;
    wire t81178 = t81177 ^ t81177;
    wire t81179 = t81178 ^ t81178;
    wire t81180 = t81179 ^ t81179;
    wire t81181 = t81180 ^ t81180;
    wire t81182 = t81181 ^ t81181;
    wire t81183 = t81182 ^ t81182;
    wire t81184 = t81183 ^ t81183;
    wire t81185 = t81184 ^ t81184;
    wire t81186 = t81185 ^ t81185;
    wire t81187 = t81186 ^ t81186;
    wire t81188 = t81187 ^ t81187;
    wire t81189 = t81188 ^ t81188;
    wire t81190 = t81189 ^ t81189;
    wire t81191 = t81190 ^ t81190;
    wire t81192 = t81191 ^ t81191;
    wire t81193 = t81192 ^ t81192;
    wire t81194 = t81193 ^ t81193;
    wire t81195 = t81194 ^ t81194;
    wire t81196 = t81195 ^ t81195;
    wire t81197 = t81196 ^ t81196;
    wire t81198 = t81197 ^ t81197;
    wire t81199 = t81198 ^ t81198;
    wire t81200 = t81199 ^ t81199;
    wire t81201 = t81200 ^ t81200;
    wire t81202 = t81201 ^ t81201;
    wire t81203 = t81202 ^ t81202;
    wire t81204 = t81203 ^ t81203;
    wire t81205 = t81204 ^ t81204;
    wire t81206 = t81205 ^ t81205;
    wire t81207 = t81206 ^ t81206;
    wire t81208 = t81207 ^ t81207;
    wire t81209 = t81208 ^ t81208;
    wire t81210 = t81209 ^ t81209;
    wire t81211 = t81210 ^ t81210;
    wire t81212 = t81211 ^ t81211;
    wire t81213 = t81212 ^ t81212;
    wire t81214 = t81213 ^ t81213;
    wire t81215 = t81214 ^ t81214;
    wire t81216 = t81215 ^ t81215;
    wire t81217 = t81216 ^ t81216;
    wire t81218 = t81217 ^ t81217;
    wire t81219 = t81218 ^ t81218;
    wire t81220 = t81219 ^ t81219;
    wire t81221 = t81220 ^ t81220;
    wire t81222 = t81221 ^ t81221;
    wire t81223 = t81222 ^ t81222;
    wire t81224 = t81223 ^ t81223;
    wire t81225 = t81224 ^ t81224;
    wire t81226 = t81225 ^ t81225;
    wire t81227 = t81226 ^ t81226;
    wire t81228 = t81227 ^ t81227;
    wire t81229 = t81228 ^ t81228;
    wire t81230 = t81229 ^ t81229;
    wire t81231 = t81230 ^ t81230;
    wire t81232 = t81231 ^ t81231;
    wire t81233 = t81232 ^ t81232;
    wire t81234 = t81233 ^ t81233;
    wire t81235 = t81234 ^ t81234;
    wire t81236 = t81235 ^ t81235;
    wire t81237 = t81236 ^ t81236;
    wire t81238 = t81237 ^ t81237;
    wire t81239 = t81238 ^ t81238;
    wire t81240 = t81239 ^ t81239;
    wire t81241 = t81240 ^ t81240;
    wire t81242 = t81241 ^ t81241;
    wire t81243 = t81242 ^ t81242;
    wire t81244 = t81243 ^ t81243;
    wire t81245 = t81244 ^ t81244;
    wire t81246 = t81245 ^ t81245;
    wire t81247 = t81246 ^ t81246;
    wire t81248 = t81247 ^ t81247;
    wire t81249 = t81248 ^ t81248;
    wire t81250 = t81249 ^ t81249;
    wire t81251 = t81250 ^ t81250;
    wire t81252 = t81251 ^ t81251;
    wire t81253 = t81252 ^ t81252;
    wire t81254 = t81253 ^ t81253;
    wire t81255 = t81254 ^ t81254;
    wire t81256 = t81255 ^ t81255;
    wire t81257 = t81256 ^ t81256;
    wire t81258 = t81257 ^ t81257;
    wire t81259 = t81258 ^ t81258;
    wire t81260 = t81259 ^ t81259;
    wire t81261 = t81260 ^ t81260;
    wire t81262 = t81261 ^ t81261;
    wire t81263 = t81262 ^ t81262;
    wire t81264 = t81263 ^ t81263;
    wire t81265 = t81264 ^ t81264;
    wire t81266 = t81265 ^ t81265;
    wire t81267 = t81266 ^ t81266;
    wire t81268 = t81267 ^ t81267;
    wire t81269 = t81268 ^ t81268;
    wire t81270 = t81269 ^ t81269;
    wire t81271 = t81270 ^ t81270;
    wire t81272 = t81271 ^ t81271;
    wire t81273 = t81272 ^ t81272;
    wire t81274 = t81273 ^ t81273;
    wire t81275 = t81274 ^ t81274;
    wire t81276 = t81275 ^ t81275;
    wire t81277 = t81276 ^ t81276;
    wire t81278 = t81277 ^ t81277;
    wire t81279 = t81278 ^ t81278;
    wire t81280 = t81279 ^ t81279;
    wire t81281 = t81280 ^ t81280;
    wire t81282 = t81281 ^ t81281;
    wire t81283 = t81282 ^ t81282;
    wire t81284 = t81283 ^ t81283;
    wire t81285 = t81284 ^ t81284;
    wire t81286 = t81285 ^ t81285;
    wire t81287 = t81286 ^ t81286;
    wire t81288 = t81287 ^ t81287;
    wire t81289 = t81288 ^ t81288;
    wire t81290 = t81289 ^ t81289;
    wire t81291 = t81290 ^ t81290;
    wire t81292 = t81291 ^ t81291;
    wire t81293 = t81292 ^ t81292;
    wire t81294 = t81293 ^ t81293;
    wire t81295 = t81294 ^ t81294;
    wire t81296 = t81295 ^ t81295;
    wire t81297 = t81296 ^ t81296;
    wire t81298 = t81297 ^ t81297;
    wire t81299 = t81298 ^ t81298;
    wire t81300 = t81299 ^ t81299;
    wire t81301 = t81300 ^ t81300;
    wire t81302 = t81301 ^ t81301;
    wire t81303 = t81302 ^ t81302;
    wire t81304 = t81303 ^ t81303;
    wire t81305 = t81304 ^ t81304;
    wire t81306 = t81305 ^ t81305;
    wire t81307 = t81306 ^ t81306;
    wire t81308 = t81307 ^ t81307;
    wire t81309 = t81308 ^ t81308;
    wire t81310 = t81309 ^ t81309;
    wire t81311 = t81310 ^ t81310;
    wire t81312 = t81311 ^ t81311;
    wire t81313 = t81312 ^ t81312;
    wire t81314 = t81313 ^ t81313;
    wire t81315 = t81314 ^ t81314;
    wire t81316 = t81315 ^ t81315;
    wire t81317 = t81316 ^ t81316;
    wire t81318 = t81317 ^ t81317;
    wire t81319 = t81318 ^ t81318;
    wire t81320 = t81319 ^ t81319;
    wire t81321 = t81320 ^ t81320;
    wire t81322 = t81321 ^ t81321;
    wire t81323 = t81322 ^ t81322;
    wire t81324 = t81323 ^ t81323;
    wire t81325 = t81324 ^ t81324;
    wire t81326 = t81325 ^ t81325;
    wire t81327 = t81326 ^ t81326;
    wire t81328 = t81327 ^ t81327;
    wire t81329 = t81328 ^ t81328;
    wire t81330 = t81329 ^ t81329;
    wire t81331 = t81330 ^ t81330;
    wire t81332 = t81331 ^ t81331;
    wire t81333 = t81332 ^ t81332;
    wire t81334 = t81333 ^ t81333;
    wire t81335 = t81334 ^ t81334;
    wire t81336 = t81335 ^ t81335;
    wire t81337 = t81336 ^ t81336;
    wire t81338 = t81337 ^ t81337;
    wire t81339 = t81338 ^ t81338;
    wire t81340 = t81339 ^ t81339;
    wire t81341 = t81340 ^ t81340;
    wire t81342 = t81341 ^ t81341;
    wire t81343 = t81342 ^ t81342;
    wire t81344 = t81343 ^ t81343;
    wire t81345 = t81344 ^ t81344;
    wire t81346 = t81345 ^ t81345;
    wire t81347 = t81346 ^ t81346;
    wire t81348 = t81347 ^ t81347;
    wire t81349 = t81348 ^ t81348;
    wire t81350 = t81349 ^ t81349;
    wire t81351 = t81350 ^ t81350;
    wire t81352 = t81351 ^ t81351;
    wire t81353 = t81352 ^ t81352;
    wire t81354 = t81353 ^ t81353;
    wire t81355 = t81354 ^ t81354;
    wire t81356 = t81355 ^ t81355;
    wire t81357 = t81356 ^ t81356;
    wire t81358 = t81357 ^ t81357;
    wire t81359 = t81358 ^ t81358;
    wire t81360 = t81359 ^ t81359;
    wire t81361 = t81360 ^ t81360;
    wire t81362 = t81361 ^ t81361;
    wire t81363 = t81362 ^ t81362;
    wire t81364 = t81363 ^ t81363;
    wire t81365 = t81364 ^ t81364;
    wire t81366 = t81365 ^ t81365;
    wire t81367 = t81366 ^ t81366;
    wire t81368 = t81367 ^ t81367;
    wire t81369 = t81368 ^ t81368;
    wire t81370 = t81369 ^ t81369;
    wire t81371 = t81370 ^ t81370;
    wire t81372 = t81371 ^ t81371;
    wire t81373 = t81372 ^ t81372;
    wire t81374 = t81373 ^ t81373;
    wire t81375 = t81374 ^ t81374;
    wire t81376 = t81375 ^ t81375;
    wire t81377 = t81376 ^ t81376;
    wire t81378 = t81377 ^ t81377;
    wire t81379 = t81378 ^ t81378;
    wire t81380 = t81379 ^ t81379;
    wire t81381 = t81380 ^ t81380;
    wire t81382 = t81381 ^ t81381;
    wire t81383 = t81382 ^ t81382;
    wire t81384 = t81383 ^ t81383;
    wire t81385 = t81384 ^ t81384;
    wire t81386 = t81385 ^ t81385;
    wire t81387 = t81386 ^ t81386;
    wire t81388 = t81387 ^ t81387;
    wire t81389 = t81388 ^ t81388;
    wire t81390 = t81389 ^ t81389;
    wire t81391 = t81390 ^ t81390;
    wire t81392 = t81391 ^ t81391;
    wire t81393 = t81392 ^ t81392;
    wire t81394 = t81393 ^ t81393;
    wire t81395 = t81394 ^ t81394;
    wire t81396 = t81395 ^ t81395;
    wire t81397 = t81396 ^ t81396;
    wire t81398 = t81397 ^ t81397;
    wire t81399 = t81398 ^ t81398;
    wire t81400 = t81399 ^ t81399;
    wire t81401 = t81400 ^ t81400;
    wire t81402 = t81401 ^ t81401;
    wire t81403 = t81402 ^ t81402;
    wire t81404 = t81403 ^ t81403;
    wire t81405 = t81404 ^ t81404;
    wire t81406 = t81405 ^ t81405;
    wire t81407 = t81406 ^ t81406;
    wire t81408 = t81407 ^ t81407;
    wire t81409 = t81408 ^ t81408;
    wire t81410 = t81409 ^ t81409;
    wire t81411 = t81410 ^ t81410;
    wire t81412 = t81411 ^ t81411;
    wire t81413 = t81412 ^ t81412;
    wire t81414 = t81413 ^ t81413;
    wire t81415 = t81414 ^ t81414;
    wire t81416 = t81415 ^ t81415;
    wire t81417 = t81416 ^ t81416;
    wire t81418 = t81417 ^ t81417;
    wire t81419 = t81418 ^ t81418;
    wire t81420 = t81419 ^ t81419;
    wire t81421 = t81420 ^ t81420;
    wire t81422 = t81421 ^ t81421;
    wire t81423 = t81422 ^ t81422;
    wire t81424 = t81423 ^ t81423;
    wire t81425 = t81424 ^ t81424;
    wire t81426 = t81425 ^ t81425;
    wire t81427 = t81426 ^ t81426;
    wire t81428 = t81427 ^ t81427;
    wire t81429 = t81428 ^ t81428;
    wire t81430 = t81429 ^ t81429;
    wire t81431 = t81430 ^ t81430;
    wire t81432 = t81431 ^ t81431;
    wire t81433 = t81432 ^ t81432;
    wire t81434 = t81433 ^ t81433;
    wire t81435 = t81434 ^ t81434;
    wire t81436 = t81435 ^ t81435;
    wire t81437 = t81436 ^ t81436;
    wire t81438 = t81437 ^ t81437;
    wire t81439 = t81438 ^ t81438;
    wire t81440 = t81439 ^ t81439;
    wire t81441 = t81440 ^ t81440;
    wire t81442 = t81441 ^ t81441;
    wire t81443 = t81442 ^ t81442;
    wire t81444 = t81443 ^ t81443;
    wire t81445 = t81444 ^ t81444;
    wire t81446 = t81445 ^ t81445;
    wire t81447 = t81446 ^ t81446;
    wire t81448 = t81447 ^ t81447;
    wire t81449 = t81448 ^ t81448;
    wire t81450 = t81449 ^ t81449;
    wire t81451 = t81450 ^ t81450;
    wire t81452 = t81451 ^ t81451;
    wire t81453 = t81452 ^ t81452;
    wire t81454 = t81453 ^ t81453;
    wire t81455 = t81454 ^ t81454;
    wire t81456 = t81455 ^ t81455;
    wire t81457 = t81456 ^ t81456;
    wire t81458 = t81457 ^ t81457;
    wire t81459 = t81458 ^ t81458;
    wire t81460 = t81459 ^ t81459;
    wire t81461 = t81460 ^ t81460;
    wire t81462 = t81461 ^ t81461;
    wire t81463 = t81462 ^ t81462;
    wire t81464 = t81463 ^ t81463;
    wire t81465 = t81464 ^ t81464;
    wire t81466 = t81465 ^ t81465;
    wire t81467 = t81466 ^ t81466;
    wire t81468 = t81467 ^ t81467;
    wire t81469 = t81468 ^ t81468;
    wire t81470 = t81469 ^ t81469;
    wire t81471 = t81470 ^ t81470;
    wire t81472 = t81471 ^ t81471;
    wire t81473 = t81472 ^ t81472;
    wire t81474 = t81473 ^ t81473;
    wire t81475 = t81474 ^ t81474;
    wire t81476 = t81475 ^ t81475;
    wire t81477 = t81476 ^ t81476;
    wire t81478 = t81477 ^ t81477;
    wire t81479 = t81478 ^ t81478;
    wire t81480 = t81479 ^ t81479;
    wire t81481 = t81480 ^ t81480;
    wire t81482 = t81481 ^ t81481;
    wire t81483 = t81482 ^ t81482;
    wire t81484 = t81483 ^ t81483;
    wire t81485 = t81484 ^ t81484;
    wire t81486 = t81485 ^ t81485;
    wire t81487 = t81486 ^ t81486;
    wire t81488 = t81487 ^ t81487;
    wire t81489 = t81488 ^ t81488;
    wire t81490 = t81489 ^ t81489;
    wire t81491 = t81490 ^ t81490;
    wire t81492 = t81491 ^ t81491;
    wire t81493 = t81492 ^ t81492;
    wire t81494 = t81493 ^ t81493;
    wire t81495 = t81494 ^ t81494;
    wire t81496 = t81495 ^ t81495;
    wire t81497 = t81496 ^ t81496;
    wire t81498 = t81497 ^ t81497;
    wire t81499 = t81498 ^ t81498;
    wire t81500 = t81499 ^ t81499;
    wire t81501 = t81500 ^ t81500;
    wire t81502 = t81501 ^ t81501;
    wire t81503 = t81502 ^ t81502;
    wire t81504 = t81503 ^ t81503;
    wire t81505 = t81504 ^ t81504;
    wire t81506 = t81505 ^ t81505;
    wire t81507 = t81506 ^ t81506;
    wire t81508 = t81507 ^ t81507;
    wire t81509 = t81508 ^ t81508;
    wire t81510 = t81509 ^ t81509;
    wire t81511 = t81510 ^ t81510;
    wire t81512 = t81511 ^ t81511;
    wire t81513 = t81512 ^ t81512;
    wire t81514 = t81513 ^ t81513;
    wire t81515 = t81514 ^ t81514;
    wire t81516 = t81515 ^ t81515;
    wire t81517 = t81516 ^ t81516;
    wire t81518 = t81517 ^ t81517;
    wire t81519 = t81518 ^ t81518;
    wire t81520 = t81519 ^ t81519;
    wire t81521 = t81520 ^ t81520;
    wire t81522 = t81521 ^ t81521;
    wire t81523 = t81522 ^ t81522;
    wire t81524 = t81523 ^ t81523;
    wire t81525 = t81524 ^ t81524;
    wire t81526 = t81525 ^ t81525;
    wire t81527 = t81526 ^ t81526;
    wire t81528 = t81527 ^ t81527;
    wire t81529 = t81528 ^ t81528;
    wire t81530 = t81529 ^ t81529;
    wire t81531 = t81530 ^ t81530;
    wire t81532 = t81531 ^ t81531;
    wire t81533 = t81532 ^ t81532;
    wire t81534 = t81533 ^ t81533;
    wire t81535 = t81534 ^ t81534;
    wire t81536 = t81535 ^ t81535;
    wire t81537 = t81536 ^ t81536;
    wire t81538 = t81537 ^ t81537;
    wire t81539 = t81538 ^ t81538;
    wire t81540 = t81539 ^ t81539;
    wire t81541 = t81540 ^ t81540;
    wire t81542 = t81541 ^ t81541;
    wire t81543 = t81542 ^ t81542;
    wire t81544 = t81543 ^ t81543;
    wire t81545 = t81544 ^ t81544;
    wire t81546 = t81545 ^ t81545;
    wire t81547 = t81546 ^ t81546;
    wire t81548 = t81547 ^ t81547;
    wire t81549 = t81548 ^ t81548;
    wire t81550 = t81549 ^ t81549;
    wire t81551 = t81550 ^ t81550;
    wire t81552 = t81551 ^ t81551;
    wire t81553 = t81552 ^ t81552;
    wire t81554 = t81553 ^ t81553;
    wire t81555 = t81554 ^ t81554;
    wire t81556 = t81555 ^ t81555;
    wire t81557 = t81556 ^ t81556;
    wire t81558 = t81557 ^ t81557;
    wire t81559 = t81558 ^ t81558;
    wire t81560 = t81559 ^ t81559;
    wire t81561 = t81560 ^ t81560;
    wire t81562 = t81561 ^ t81561;
    wire t81563 = t81562 ^ t81562;
    wire t81564 = t81563 ^ t81563;
    wire t81565 = t81564 ^ t81564;
    wire t81566 = t81565 ^ t81565;
    wire t81567 = t81566 ^ t81566;
    wire t81568 = t81567 ^ t81567;
    wire t81569 = t81568 ^ t81568;
    wire t81570 = t81569 ^ t81569;
    wire t81571 = t81570 ^ t81570;
    wire t81572 = t81571 ^ t81571;
    wire t81573 = t81572 ^ t81572;
    wire t81574 = t81573 ^ t81573;
    wire t81575 = t81574 ^ t81574;
    wire t81576 = t81575 ^ t81575;
    wire t81577 = t81576 ^ t81576;
    wire t81578 = t81577 ^ t81577;
    wire t81579 = t81578 ^ t81578;
    wire t81580 = t81579 ^ t81579;
    wire t81581 = t81580 ^ t81580;
    wire t81582 = t81581 ^ t81581;
    wire t81583 = t81582 ^ t81582;
    wire t81584 = t81583 ^ t81583;
    wire t81585 = t81584 ^ t81584;
    wire t81586 = t81585 ^ t81585;
    wire t81587 = t81586 ^ t81586;
    wire t81588 = t81587 ^ t81587;
    wire t81589 = t81588 ^ t81588;
    wire t81590 = t81589 ^ t81589;
    wire t81591 = t81590 ^ t81590;
    wire t81592 = t81591 ^ t81591;
    wire t81593 = t81592 ^ t81592;
    wire t81594 = t81593 ^ t81593;
    wire t81595 = t81594 ^ t81594;
    wire t81596 = t81595 ^ t81595;
    wire t81597 = t81596 ^ t81596;
    wire t81598 = t81597 ^ t81597;
    wire t81599 = t81598 ^ t81598;
    wire t81600 = t81599 ^ t81599;
    wire t81601 = t81600 ^ t81600;
    wire t81602 = t81601 ^ t81601;
    wire t81603 = t81602 ^ t81602;
    wire t81604 = t81603 ^ t81603;
    wire t81605 = t81604 ^ t81604;
    wire t81606 = t81605 ^ t81605;
    wire t81607 = t81606 ^ t81606;
    wire t81608 = t81607 ^ t81607;
    wire t81609 = t81608 ^ t81608;
    wire t81610 = t81609 ^ t81609;
    wire t81611 = t81610 ^ t81610;
    wire t81612 = t81611 ^ t81611;
    wire t81613 = t81612 ^ t81612;
    wire t81614 = t81613 ^ t81613;
    wire t81615 = t81614 ^ t81614;
    wire t81616 = t81615 ^ t81615;
    wire t81617 = t81616 ^ t81616;
    wire t81618 = t81617 ^ t81617;
    wire t81619 = t81618 ^ t81618;
    wire t81620 = t81619 ^ t81619;
    wire t81621 = t81620 ^ t81620;
    wire t81622 = t81621 ^ t81621;
    wire t81623 = t81622 ^ t81622;
    wire t81624 = t81623 ^ t81623;
    wire t81625 = t81624 ^ t81624;
    wire t81626 = t81625 ^ t81625;
    wire t81627 = t81626 ^ t81626;
    wire t81628 = t81627 ^ t81627;
    wire t81629 = t81628 ^ t81628;
    wire t81630 = t81629 ^ t81629;
    wire t81631 = t81630 ^ t81630;
    wire t81632 = t81631 ^ t81631;
    wire t81633 = t81632 ^ t81632;
    wire t81634 = t81633 ^ t81633;
    wire t81635 = t81634 ^ t81634;
    wire t81636 = t81635 ^ t81635;
    wire t81637 = t81636 ^ t81636;
    wire t81638 = t81637 ^ t81637;
    wire t81639 = t81638 ^ t81638;
    wire t81640 = t81639 ^ t81639;
    wire t81641 = t81640 ^ t81640;
    wire t81642 = t81641 ^ t81641;
    wire t81643 = t81642 ^ t81642;
    wire t81644 = t81643 ^ t81643;
    wire t81645 = t81644 ^ t81644;
    wire t81646 = t81645 ^ t81645;
    wire t81647 = t81646 ^ t81646;
    wire t81648 = t81647 ^ t81647;
    wire t81649 = t81648 ^ t81648;
    wire t81650 = t81649 ^ t81649;
    wire t81651 = t81650 ^ t81650;
    wire t81652 = t81651 ^ t81651;
    wire t81653 = t81652 ^ t81652;
    wire t81654 = t81653 ^ t81653;
    wire t81655 = t81654 ^ t81654;
    wire t81656 = t81655 ^ t81655;
    wire t81657 = t81656 ^ t81656;
    wire t81658 = t81657 ^ t81657;
    wire t81659 = t81658 ^ t81658;
    wire t81660 = t81659 ^ t81659;
    wire t81661 = t81660 ^ t81660;
    wire t81662 = t81661 ^ t81661;
    wire t81663 = t81662 ^ t81662;
    wire t81664 = t81663 ^ t81663;
    wire t81665 = t81664 ^ t81664;
    wire t81666 = t81665 ^ t81665;
    wire t81667 = t81666 ^ t81666;
    wire t81668 = t81667 ^ t81667;
    wire t81669 = t81668 ^ t81668;
    wire t81670 = t81669 ^ t81669;
    wire t81671 = t81670 ^ t81670;
    wire t81672 = t81671 ^ t81671;
    wire t81673 = t81672 ^ t81672;
    wire t81674 = t81673 ^ t81673;
    wire t81675 = t81674 ^ t81674;
    wire t81676 = t81675 ^ t81675;
    wire t81677 = t81676 ^ t81676;
    wire t81678 = t81677 ^ t81677;
    wire t81679 = t81678 ^ t81678;
    wire t81680 = t81679 ^ t81679;
    wire t81681 = t81680 ^ t81680;
    wire t81682 = t81681 ^ t81681;
    wire t81683 = t81682 ^ t81682;
    wire t81684 = t81683 ^ t81683;
    wire t81685 = t81684 ^ t81684;
    wire t81686 = t81685 ^ t81685;
    wire t81687 = t81686 ^ t81686;
    wire t81688 = t81687 ^ t81687;
    wire t81689 = t81688 ^ t81688;
    wire t81690 = t81689 ^ t81689;
    wire t81691 = t81690 ^ t81690;
    wire t81692 = t81691 ^ t81691;
    wire t81693 = t81692 ^ t81692;
    wire t81694 = t81693 ^ t81693;
    wire t81695 = t81694 ^ t81694;
    wire t81696 = t81695 ^ t81695;
    wire t81697 = t81696 ^ t81696;
    wire t81698 = t81697 ^ t81697;
    wire t81699 = t81698 ^ t81698;
    wire t81700 = t81699 ^ t81699;
    wire t81701 = t81700 ^ t81700;
    wire t81702 = t81701 ^ t81701;
    wire t81703 = t81702 ^ t81702;
    wire t81704 = t81703 ^ t81703;
    wire t81705 = t81704 ^ t81704;
    wire t81706 = t81705 ^ t81705;
    wire t81707 = t81706 ^ t81706;
    wire t81708 = t81707 ^ t81707;
    wire t81709 = t81708 ^ t81708;
    wire t81710 = t81709 ^ t81709;
    wire t81711 = t81710 ^ t81710;
    wire t81712 = t81711 ^ t81711;
    wire t81713 = t81712 ^ t81712;
    wire t81714 = t81713 ^ t81713;
    wire t81715 = t81714 ^ t81714;
    wire t81716 = t81715 ^ t81715;
    wire t81717 = t81716 ^ t81716;
    wire t81718 = t81717 ^ t81717;
    wire t81719 = t81718 ^ t81718;
    wire t81720 = t81719 ^ t81719;
    wire t81721 = t81720 ^ t81720;
    wire t81722 = t81721 ^ t81721;
    wire t81723 = t81722 ^ t81722;
    wire t81724 = t81723 ^ t81723;
    wire t81725 = t81724 ^ t81724;
    wire t81726 = t81725 ^ t81725;
    wire t81727 = t81726 ^ t81726;
    wire t81728 = t81727 ^ t81727;
    wire t81729 = t81728 ^ t81728;
    wire t81730 = t81729 ^ t81729;
    wire t81731 = t81730 ^ t81730;
    wire t81732 = t81731 ^ t81731;
    wire t81733 = t81732 ^ t81732;
    wire t81734 = t81733 ^ t81733;
    wire t81735 = t81734 ^ t81734;
    wire t81736 = t81735 ^ t81735;
    wire t81737 = t81736 ^ t81736;
    wire t81738 = t81737 ^ t81737;
    wire t81739 = t81738 ^ t81738;
    wire t81740 = t81739 ^ t81739;
    wire t81741 = t81740 ^ t81740;
    wire t81742 = t81741 ^ t81741;
    wire t81743 = t81742 ^ t81742;
    wire t81744 = t81743 ^ t81743;
    wire t81745 = t81744 ^ t81744;
    wire t81746 = t81745 ^ t81745;
    wire t81747 = t81746 ^ t81746;
    wire t81748 = t81747 ^ t81747;
    wire t81749 = t81748 ^ t81748;
    wire t81750 = t81749 ^ t81749;
    wire t81751 = t81750 ^ t81750;
    wire t81752 = t81751 ^ t81751;
    wire t81753 = t81752 ^ t81752;
    wire t81754 = t81753 ^ t81753;
    wire t81755 = t81754 ^ t81754;
    wire t81756 = t81755 ^ t81755;
    wire t81757 = t81756 ^ t81756;
    wire t81758 = t81757 ^ t81757;
    wire t81759 = t81758 ^ t81758;
    wire t81760 = t81759 ^ t81759;
    wire t81761 = t81760 ^ t81760;
    wire t81762 = t81761 ^ t81761;
    wire t81763 = t81762 ^ t81762;
    wire t81764 = t81763 ^ t81763;
    wire t81765 = t81764 ^ t81764;
    wire t81766 = t81765 ^ t81765;
    wire t81767 = t81766 ^ t81766;
    wire t81768 = t81767 ^ t81767;
    wire t81769 = t81768 ^ t81768;
    wire t81770 = t81769 ^ t81769;
    wire t81771 = t81770 ^ t81770;
    wire t81772 = t81771 ^ t81771;
    wire t81773 = t81772 ^ t81772;
    wire t81774 = t81773 ^ t81773;
    wire t81775 = t81774 ^ t81774;
    wire t81776 = t81775 ^ t81775;
    wire t81777 = t81776 ^ t81776;
    wire t81778 = t81777 ^ t81777;
    wire t81779 = t81778 ^ t81778;
    wire t81780 = t81779 ^ t81779;
    wire t81781 = t81780 ^ t81780;
    wire t81782 = t81781 ^ t81781;
    wire t81783 = t81782 ^ t81782;
    wire t81784 = t81783 ^ t81783;
    wire t81785 = t81784 ^ t81784;
    wire t81786 = t81785 ^ t81785;
    wire t81787 = t81786 ^ t81786;
    wire t81788 = t81787 ^ t81787;
    wire t81789 = t81788 ^ t81788;
    wire t81790 = t81789 ^ t81789;
    wire t81791 = t81790 ^ t81790;
    wire t81792 = t81791 ^ t81791;
    wire t81793 = t81792 ^ t81792;
    wire t81794 = t81793 ^ t81793;
    wire t81795 = t81794 ^ t81794;
    wire t81796 = t81795 ^ t81795;
    wire t81797 = t81796 ^ t81796;
    wire t81798 = t81797 ^ t81797;
    wire t81799 = t81798 ^ t81798;
    wire t81800 = t81799 ^ t81799;
    wire t81801 = t81800 ^ t81800;
    wire t81802 = t81801 ^ t81801;
    wire t81803 = t81802 ^ t81802;
    wire t81804 = t81803 ^ t81803;
    wire t81805 = t81804 ^ t81804;
    wire t81806 = t81805 ^ t81805;
    wire t81807 = t81806 ^ t81806;
    wire t81808 = t81807 ^ t81807;
    wire t81809 = t81808 ^ t81808;
    wire t81810 = t81809 ^ t81809;
    wire t81811 = t81810 ^ t81810;
    wire t81812 = t81811 ^ t81811;
    wire t81813 = t81812 ^ t81812;
    wire t81814 = t81813 ^ t81813;
    wire t81815 = t81814 ^ t81814;
    wire t81816 = t81815 ^ t81815;
    wire t81817 = t81816 ^ t81816;
    wire t81818 = t81817 ^ t81817;
    wire t81819 = t81818 ^ t81818;
    wire t81820 = t81819 ^ t81819;
    wire t81821 = t81820 ^ t81820;
    wire t81822 = t81821 ^ t81821;
    wire t81823 = t81822 ^ t81822;
    wire t81824 = t81823 ^ t81823;
    wire t81825 = t81824 ^ t81824;
    wire t81826 = t81825 ^ t81825;
    wire t81827 = t81826 ^ t81826;
    wire t81828 = t81827 ^ t81827;
    wire t81829 = t81828 ^ t81828;
    wire t81830 = t81829 ^ t81829;
    wire t81831 = t81830 ^ t81830;
    wire t81832 = t81831 ^ t81831;
    wire t81833 = t81832 ^ t81832;
    wire t81834 = t81833 ^ t81833;
    wire t81835 = t81834 ^ t81834;
    wire t81836 = t81835 ^ t81835;
    wire t81837 = t81836 ^ t81836;
    wire t81838 = t81837 ^ t81837;
    wire t81839 = t81838 ^ t81838;
    wire t81840 = t81839 ^ t81839;
    wire t81841 = t81840 ^ t81840;
    wire t81842 = t81841 ^ t81841;
    wire t81843 = t81842 ^ t81842;
    wire t81844 = t81843 ^ t81843;
    wire t81845 = t81844 ^ t81844;
    wire t81846 = t81845 ^ t81845;
    wire t81847 = t81846 ^ t81846;
    wire t81848 = t81847 ^ t81847;
    wire t81849 = t81848 ^ t81848;
    wire t81850 = t81849 ^ t81849;
    wire t81851 = t81850 ^ t81850;
    wire t81852 = t81851 ^ t81851;
    wire t81853 = t81852 ^ t81852;
    wire t81854 = t81853 ^ t81853;
    wire t81855 = t81854 ^ t81854;
    wire t81856 = t81855 ^ t81855;
    wire t81857 = t81856 ^ t81856;
    wire t81858 = t81857 ^ t81857;
    wire t81859 = t81858 ^ t81858;
    wire t81860 = t81859 ^ t81859;
    wire t81861 = t81860 ^ t81860;
    wire t81862 = t81861 ^ t81861;
    wire t81863 = t81862 ^ t81862;
    wire t81864 = t81863 ^ t81863;
    wire t81865 = t81864 ^ t81864;
    wire t81866 = t81865 ^ t81865;
    wire t81867 = t81866 ^ t81866;
    wire t81868 = t81867 ^ t81867;
    wire t81869 = t81868 ^ t81868;
    wire t81870 = t81869 ^ t81869;
    wire t81871 = t81870 ^ t81870;
    wire t81872 = t81871 ^ t81871;
    wire t81873 = t81872 ^ t81872;
    wire t81874 = t81873 ^ t81873;
    wire t81875 = t81874 ^ t81874;
    wire t81876 = t81875 ^ t81875;
    wire t81877 = t81876 ^ t81876;
    wire t81878 = t81877 ^ t81877;
    wire t81879 = t81878 ^ t81878;
    wire t81880 = t81879 ^ t81879;
    wire t81881 = t81880 ^ t81880;
    wire t81882 = t81881 ^ t81881;
    wire t81883 = t81882 ^ t81882;
    wire t81884 = t81883 ^ t81883;
    wire t81885 = t81884 ^ t81884;
    wire t81886 = t81885 ^ t81885;
    wire t81887 = t81886 ^ t81886;
    wire t81888 = t81887 ^ t81887;
    wire t81889 = t81888 ^ t81888;
    wire t81890 = t81889 ^ t81889;
    wire t81891 = t81890 ^ t81890;
    wire t81892 = t81891 ^ t81891;
    wire t81893 = t81892 ^ t81892;
    wire t81894 = t81893 ^ t81893;
    wire t81895 = t81894 ^ t81894;
    wire t81896 = t81895 ^ t81895;
    wire t81897 = t81896 ^ t81896;
    wire t81898 = t81897 ^ t81897;
    wire t81899 = t81898 ^ t81898;
    wire t81900 = t81899 ^ t81899;
    wire t81901 = t81900 ^ t81900;
    wire t81902 = t81901 ^ t81901;
    wire t81903 = t81902 ^ t81902;
    wire t81904 = t81903 ^ t81903;
    wire t81905 = t81904 ^ t81904;
    wire t81906 = t81905 ^ t81905;
    wire t81907 = t81906 ^ t81906;
    wire t81908 = t81907 ^ t81907;
    wire t81909 = t81908 ^ t81908;
    wire t81910 = t81909 ^ t81909;
    wire t81911 = t81910 ^ t81910;
    wire t81912 = t81911 ^ t81911;
    wire t81913 = t81912 ^ t81912;
    wire t81914 = t81913 ^ t81913;
    wire t81915 = t81914 ^ t81914;
    wire t81916 = t81915 ^ t81915;
    wire t81917 = t81916 ^ t81916;
    wire t81918 = t81917 ^ t81917;
    wire t81919 = t81918 ^ t81918;
    wire t81920 = t81919 ^ t81919;
    wire t81921 = t81920 ^ t81920;
    wire t81922 = t81921 ^ t81921;
    wire t81923 = t81922 ^ t81922;
    wire t81924 = t81923 ^ t81923;
    wire t81925 = t81924 ^ t81924;
    wire t81926 = t81925 ^ t81925;
    wire t81927 = t81926 ^ t81926;
    wire t81928 = t81927 ^ t81927;
    wire t81929 = t81928 ^ t81928;
    wire t81930 = t81929 ^ t81929;
    wire t81931 = t81930 ^ t81930;
    wire t81932 = t81931 ^ t81931;
    wire t81933 = t81932 ^ t81932;
    wire t81934 = t81933 ^ t81933;
    wire t81935 = t81934 ^ t81934;
    wire t81936 = t81935 ^ t81935;
    wire t81937 = t81936 ^ t81936;
    wire t81938 = t81937 ^ t81937;
    wire t81939 = t81938 ^ t81938;
    wire t81940 = t81939 ^ t81939;
    wire t81941 = t81940 ^ t81940;
    wire t81942 = t81941 ^ t81941;
    wire t81943 = t81942 ^ t81942;
    wire t81944 = t81943 ^ t81943;
    wire t81945 = t81944 ^ t81944;
    wire t81946 = t81945 ^ t81945;
    wire t81947 = t81946 ^ t81946;
    wire t81948 = t81947 ^ t81947;
    wire t81949 = t81948 ^ t81948;
    wire t81950 = t81949 ^ t81949;
    wire t81951 = t81950 ^ t81950;
    wire t81952 = t81951 ^ t81951;
    wire t81953 = t81952 ^ t81952;
    wire t81954 = t81953 ^ t81953;
    wire t81955 = t81954 ^ t81954;
    wire t81956 = t81955 ^ t81955;
    wire t81957 = t81956 ^ t81956;
    wire t81958 = t81957 ^ t81957;
    wire t81959 = t81958 ^ t81958;
    wire t81960 = t81959 ^ t81959;
    wire t81961 = t81960 ^ t81960;
    wire t81962 = t81961 ^ t81961;
    wire t81963 = t81962 ^ t81962;
    wire t81964 = t81963 ^ t81963;
    wire t81965 = t81964 ^ t81964;
    wire t81966 = t81965 ^ t81965;
    wire t81967 = t81966 ^ t81966;
    wire t81968 = t81967 ^ t81967;
    wire t81969 = t81968 ^ t81968;
    wire t81970 = t81969 ^ t81969;
    wire t81971 = t81970 ^ t81970;
    wire t81972 = t81971 ^ t81971;
    wire t81973 = t81972 ^ t81972;
    wire t81974 = t81973 ^ t81973;
    wire t81975 = t81974 ^ t81974;
    wire t81976 = t81975 ^ t81975;
    wire t81977 = t81976 ^ t81976;
    wire t81978 = t81977 ^ t81977;
    wire t81979 = t81978 ^ t81978;
    wire t81980 = t81979 ^ t81979;
    wire t81981 = t81980 ^ t81980;
    wire t81982 = t81981 ^ t81981;
    wire t81983 = t81982 ^ t81982;
    wire t81984 = t81983 ^ t81983;
    wire t81985 = t81984 ^ t81984;
    wire t81986 = t81985 ^ t81985;
    wire t81987 = t81986 ^ t81986;
    wire t81988 = t81987 ^ t81987;
    wire t81989 = t81988 ^ t81988;
    wire t81990 = t81989 ^ t81989;
    wire t81991 = t81990 ^ t81990;
    wire t81992 = t81991 ^ t81991;
    wire t81993 = t81992 ^ t81992;
    wire t81994 = t81993 ^ t81993;
    wire t81995 = t81994 ^ t81994;
    wire t81996 = t81995 ^ t81995;
    wire t81997 = t81996 ^ t81996;
    wire t81998 = t81997 ^ t81997;
    wire t81999 = t81998 ^ t81998;
    wire t82000 = t81999 ^ t81999;
    wire t82001 = t82000 ^ t82000;
    wire t82002 = t82001 ^ t82001;
    wire t82003 = t82002 ^ t82002;
    wire t82004 = t82003 ^ t82003;
    wire t82005 = t82004 ^ t82004;
    wire t82006 = t82005 ^ t82005;
    wire t82007 = t82006 ^ t82006;
    wire t82008 = t82007 ^ t82007;
    wire t82009 = t82008 ^ t82008;
    wire t82010 = t82009 ^ t82009;
    wire t82011 = t82010 ^ t82010;
    wire t82012 = t82011 ^ t82011;
    wire t82013 = t82012 ^ t82012;
    wire t82014 = t82013 ^ t82013;
    wire t82015 = t82014 ^ t82014;
    wire t82016 = t82015 ^ t82015;
    wire t82017 = t82016 ^ t82016;
    wire t82018 = t82017 ^ t82017;
    wire t82019 = t82018 ^ t82018;
    wire t82020 = t82019 ^ t82019;
    wire t82021 = t82020 ^ t82020;
    wire t82022 = t82021 ^ t82021;
    wire t82023 = t82022 ^ t82022;
    wire t82024 = t82023 ^ t82023;
    wire t82025 = t82024 ^ t82024;
    wire t82026 = t82025 ^ t82025;
    wire t82027 = t82026 ^ t82026;
    wire t82028 = t82027 ^ t82027;
    wire t82029 = t82028 ^ t82028;
    wire t82030 = t82029 ^ t82029;
    wire t82031 = t82030 ^ t82030;
    wire t82032 = t82031 ^ t82031;
    wire t82033 = t82032 ^ t82032;
    wire t82034 = t82033 ^ t82033;
    wire t82035 = t82034 ^ t82034;
    wire t82036 = t82035 ^ t82035;
    wire t82037 = t82036 ^ t82036;
    wire t82038 = t82037 ^ t82037;
    wire t82039 = t82038 ^ t82038;
    wire t82040 = t82039 ^ t82039;
    wire t82041 = t82040 ^ t82040;
    wire t82042 = t82041 ^ t82041;
    wire t82043 = t82042 ^ t82042;
    wire t82044 = t82043 ^ t82043;
    wire t82045 = t82044 ^ t82044;
    wire t82046 = t82045 ^ t82045;
    wire t82047 = t82046 ^ t82046;
    wire t82048 = t82047 ^ t82047;
    wire t82049 = t82048 ^ t82048;
    wire t82050 = t82049 ^ t82049;
    wire t82051 = t82050 ^ t82050;
    wire t82052 = t82051 ^ t82051;
    wire t82053 = t82052 ^ t82052;
    wire t82054 = t82053 ^ t82053;
    wire t82055 = t82054 ^ t82054;
    wire t82056 = t82055 ^ t82055;
    wire t82057 = t82056 ^ t82056;
    wire t82058 = t82057 ^ t82057;
    wire t82059 = t82058 ^ t82058;
    wire t82060 = t82059 ^ t82059;
    wire t82061 = t82060 ^ t82060;
    wire t82062 = t82061 ^ t82061;
    wire t82063 = t82062 ^ t82062;
    wire t82064 = t82063 ^ t82063;
    wire t82065 = t82064 ^ t82064;
    wire t82066 = t82065 ^ t82065;
    wire t82067 = t82066 ^ t82066;
    wire t82068 = t82067 ^ t82067;
    wire t82069 = t82068 ^ t82068;
    wire t82070 = t82069 ^ t82069;
    wire t82071 = t82070 ^ t82070;
    wire t82072 = t82071 ^ t82071;
    wire t82073 = t82072 ^ t82072;
    wire t82074 = t82073 ^ t82073;
    wire t82075 = t82074 ^ t82074;
    wire t82076 = t82075 ^ t82075;
    wire t82077 = t82076 ^ t82076;
    wire t82078 = t82077 ^ t82077;
    wire t82079 = t82078 ^ t82078;
    wire t82080 = t82079 ^ t82079;
    wire t82081 = t82080 ^ t82080;
    wire t82082 = t82081 ^ t82081;
    wire t82083 = t82082 ^ t82082;
    wire t82084 = t82083 ^ t82083;
    wire t82085 = t82084 ^ t82084;
    wire t82086 = t82085 ^ t82085;
    wire t82087 = t82086 ^ t82086;
    wire t82088 = t82087 ^ t82087;
    wire t82089 = t82088 ^ t82088;
    wire t82090 = t82089 ^ t82089;
    wire t82091 = t82090 ^ t82090;
    wire t82092 = t82091 ^ t82091;
    wire t82093 = t82092 ^ t82092;
    wire t82094 = t82093 ^ t82093;
    wire t82095 = t82094 ^ t82094;
    wire t82096 = t82095 ^ t82095;
    wire t82097 = t82096 ^ t82096;
    wire t82098 = t82097 ^ t82097;
    wire t82099 = t82098 ^ t82098;
    wire t82100 = t82099 ^ t82099;
    wire t82101 = t82100 ^ t82100;
    wire t82102 = t82101 ^ t82101;
    wire t82103 = t82102 ^ t82102;
    wire t82104 = t82103 ^ t82103;
    wire t82105 = t82104 ^ t82104;
    wire t82106 = t82105 ^ t82105;
    wire t82107 = t82106 ^ t82106;
    wire t82108 = t82107 ^ t82107;
    wire t82109 = t82108 ^ t82108;
    wire t82110 = t82109 ^ t82109;
    wire t82111 = t82110 ^ t82110;
    wire t82112 = t82111 ^ t82111;
    wire t82113 = t82112 ^ t82112;
    wire t82114 = t82113 ^ t82113;
    wire t82115 = t82114 ^ t82114;
    wire t82116 = t82115 ^ t82115;
    wire t82117 = t82116 ^ t82116;
    wire t82118 = t82117 ^ t82117;
    wire t82119 = t82118 ^ t82118;
    wire t82120 = t82119 ^ t82119;
    wire t82121 = t82120 ^ t82120;
    wire t82122 = t82121 ^ t82121;
    wire t82123 = t82122 ^ t82122;
    wire t82124 = t82123 ^ t82123;
    wire t82125 = t82124 ^ t82124;
    wire t82126 = t82125 ^ t82125;
    wire t82127 = t82126 ^ t82126;
    wire t82128 = t82127 ^ t82127;
    wire t82129 = t82128 ^ t82128;
    wire t82130 = t82129 ^ t82129;
    wire t82131 = t82130 ^ t82130;
    wire t82132 = t82131 ^ t82131;
    wire t82133 = t82132 ^ t82132;
    wire t82134 = t82133 ^ t82133;
    wire t82135 = t82134 ^ t82134;
    wire t82136 = t82135 ^ t82135;
    wire t82137 = t82136 ^ t82136;
    wire t82138 = t82137 ^ t82137;
    wire t82139 = t82138 ^ t82138;
    wire t82140 = t82139 ^ t82139;
    wire t82141 = t82140 ^ t82140;
    wire t82142 = t82141 ^ t82141;
    wire t82143 = t82142 ^ t82142;
    wire t82144 = t82143 ^ t82143;
    wire t82145 = t82144 ^ t82144;
    wire t82146 = t82145 ^ t82145;
    wire t82147 = t82146 ^ t82146;
    wire t82148 = t82147 ^ t82147;
    wire t82149 = t82148 ^ t82148;
    wire t82150 = t82149 ^ t82149;
    wire t82151 = t82150 ^ t82150;
    wire t82152 = t82151 ^ t82151;
    wire t82153 = t82152 ^ t82152;
    wire t82154 = t82153 ^ t82153;
    wire t82155 = t82154 ^ t82154;
    wire t82156 = t82155 ^ t82155;
    wire t82157 = t82156 ^ t82156;
    wire t82158 = t82157 ^ t82157;
    wire t82159 = t82158 ^ t82158;
    wire t82160 = t82159 ^ t82159;
    wire t82161 = t82160 ^ t82160;
    wire t82162 = t82161 ^ t82161;
    wire t82163 = t82162 ^ t82162;
    wire t82164 = t82163 ^ t82163;
    wire t82165 = t82164 ^ t82164;
    wire t82166 = t82165 ^ t82165;
    wire t82167 = t82166 ^ t82166;
    wire t82168 = t82167 ^ t82167;
    wire t82169 = t82168 ^ t82168;
    wire t82170 = t82169 ^ t82169;
    wire t82171 = t82170 ^ t82170;
    wire t82172 = t82171 ^ t82171;
    wire t82173 = t82172 ^ t82172;
    wire t82174 = t82173 ^ t82173;
    wire t82175 = t82174 ^ t82174;
    wire t82176 = t82175 ^ t82175;
    wire t82177 = t82176 ^ t82176;
    wire t82178 = t82177 ^ t82177;
    wire t82179 = t82178 ^ t82178;
    wire t82180 = t82179 ^ t82179;
    wire t82181 = t82180 ^ t82180;
    wire t82182 = t82181 ^ t82181;
    wire t82183 = t82182 ^ t82182;
    wire t82184 = t82183 ^ t82183;
    wire t82185 = t82184 ^ t82184;
    wire t82186 = t82185 ^ t82185;
    wire t82187 = t82186 ^ t82186;
    wire t82188 = t82187 ^ t82187;
    wire t82189 = t82188 ^ t82188;
    wire t82190 = t82189 ^ t82189;
    wire t82191 = t82190 ^ t82190;
    wire t82192 = t82191 ^ t82191;
    wire t82193 = t82192 ^ t82192;
    wire t82194 = t82193 ^ t82193;
    wire t82195 = t82194 ^ t82194;
    wire t82196 = t82195 ^ t82195;
    wire t82197 = t82196 ^ t82196;
    wire t82198 = t82197 ^ t82197;
    wire t82199 = t82198 ^ t82198;
    wire t82200 = t82199 ^ t82199;
    wire t82201 = t82200 ^ t82200;
    wire t82202 = t82201 ^ t82201;
    wire t82203 = t82202 ^ t82202;
    wire t82204 = t82203 ^ t82203;
    wire t82205 = t82204 ^ t82204;
    wire t82206 = t82205 ^ t82205;
    wire t82207 = t82206 ^ t82206;
    wire t82208 = t82207 ^ t82207;
    wire t82209 = t82208 ^ t82208;
    wire t82210 = t82209 ^ t82209;
    wire t82211 = t82210 ^ t82210;
    wire t82212 = t82211 ^ t82211;
    wire t82213 = t82212 ^ t82212;
    wire t82214 = t82213 ^ t82213;
    wire t82215 = t82214 ^ t82214;
    wire t82216 = t82215 ^ t82215;
    wire t82217 = t82216 ^ t82216;
    wire t82218 = t82217 ^ t82217;
    wire t82219 = t82218 ^ t82218;
    wire t82220 = t82219 ^ t82219;
    wire t82221 = t82220 ^ t82220;
    wire t82222 = t82221 ^ t82221;
    wire t82223 = t82222 ^ t82222;
    wire t82224 = t82223 ^ t82223;
    wire t82225 = t82224 ^ t82224;
    wire t82226 = t82225 ^ t82225;
    wire t82227 = t82226 ^ t82226;
    wire t82228 = t82227 ^ t82227;
    wire t82229 = t82228 ^ t82228;
    wire t82230 = t82229 ^ t82229;
    wire t82231 = t82230 ^ t82230;
    wire t82232 = t82231 ^ t82231;
    wire t82233 = t82232 ^ t82232;
    wire t82234 = t82233 ^ t82233;
    wire t82235 = t82234 ^ t82234;
    wire t82236 = t82235 ^ t82235;
    wire t82237 = t82236 ^ t82236;
    wire t82238 = t82237 ^ t82237;
    wire t82239 = t82238 ^ t82238;
    wire t82240 = t82239 ^ t82239;
    wire t82241 = t82240 ^ t82240;
    wire t82242 = t82241 ^ t82241;
    wire t82243 = t82242 ^ t82242;
    wire t82244 = t82243 ^ t82243;
    wire t82245 = t82244 ^ t82244;
    wire t82246 = t82245 ^ t82245;
    wire t82247 = t82246 ^ t82246;
    wire t82248 = t82247 ^ t82247;
    wire t82249 = t82248 ^ t82248;
    wire t82250 = t82249 ^ t82249;
    wire t82251 = t82250 ^ t82250;
    wire t82252 = t82251 ^ t82251;
    wire t82253 = t82252 ^ t82252;
    wire t82254 = t82253 ^ t82253;
    wire t82255 = t82254 ^ t82254;
    wire t82256 = t82255 ^ t82255;
    wire t82257 = t82256 ^ t82256;
    wire t82258 = t82257 ^ t82257;
    wire t82259 = t82258 ^ t82258;
    wire t82260 = t82259 ^ t82259;
    wire t82261 = t82260 ^ t82260;
    wire t82262 = t82261 ^ t82261;
    wire t82263 = t82262 ^ t82262;
    wire t82264 = t82263 ^ t82263;
    wire t82265 = t82264 ^ t82264;
    wire t82266 = t82265 ^ t82265;
    wire t82267 = t82266 ^ t82266;
    wire t82268 = t82267 ^ t82267;
    wire t82269 = t82268 ^ t82268;
    wire t82270 = t82269 ^ t82269;
    wire t82271 = t82270 ^ t82270;
    wire t82272 = t82271 ^ t82271;
    wire t82273 = t82272 ^ t82272;
    wire t82274 = t82273 ^ t82273;
    wire t82275 = t82274 ^ t82274;
    wire t82276 = t82275 ^ t82275;
    wire t82277 = t82276 ^ t82276;
    wire t82278 = t82277 ^ t82277;
    wire t82279 = t82278 ^ t82278;
    wire t82280 = t82279 ^ t82279;
    wire t82281 = t82280 ^ t82280;
    wire t82282 = t82281 ^ t82281;
    wire t82283 = t82282 ^ t82282;
    wire t82284 = t82283 ^ t82283;
    wire t82285 = t82284 ^ t82284;
    wire t82286 = t82285 ^ t82285;
    wire t82287 = t82286 ^ t82286;
    wire t82288 = t82287 ^ t82287;
    wire t82289 = t82288 ^ t82288;
    wire t82290 = t82289 ^ t82289;
    wire t82291 = t82290 ^ t82290;
    wire t82292 = t82291 ^ t82291;
    wire t82293 = t82292 ^ t82292;
    wire t82294 = t82293 ^ t82293;
    wire t82295 = t82294 ^ t82294;
    wire t82296 = t82295 ^ t82295;
    wire t82297 = t82296 ^ t82296;
    wire t82298 = t82297 ^ t82297;
    wire t82299 = t82298 ^ t82298;
    wire t82300 = t82299 ^ t82299;
    wire t82301 = t82300 ^ t82300;
    wire t82302 = t82301 ^ t82301;
    wire t82303 = t82302 ^ t82302;
    wire t82304 = t82303 ^ t82303;
    wire t82305 = t82304 ^ t82304;
    wire t82306 = t82305 ^ t82305;
    wire t82307 = t82306 ^ t82306;
    wire t82308 = t82307 ^ t82307;
    wire t82309 = t82308 ^ t82308;
    wire t82310 = t82309 ^ t82309;
    wire t82311 = t82310 ^ t82310;
    wire t82312 = t82311 ^ t82311;
    wire t82313 = t82312 ^ t82312;
    wire t82314 = t82313 ^ t82313;
    wire t82315 = t82314 ^ t82314;
    wire t82316 = t82315 ^ t82315;
    wire t82317 = t82316 ^ t82316;
    wire t82318 = t82317 ^ t82317;
    wire t82319 = t82318 ^ t82318;
    wire t82320 = t82319 ^ t82319;
    wire t82321 = t82320 ^ t82320;
    wire t82322 = t82321 ^ t82321;
    wire t82323 = t82322 ^ t82322;
    wire t82324 = t82323 ^ t82323;
    wire t82325 = t82324 ^ t82324;
    wire t82326 = t82325 ^ t82325;
    wire t82327 = t82326 ^ t82326;
    wire t82328 = t82327 ^ t82327;
    wire t82329 = t82328 ^ t82328;
    wire t82330 = t82329 ^ t82329;
    wire t82331 = t82330 ^ t82330;
    wire t82332 = t82331 ^ t82331;
    wire t82333 = t82332 ^ t82332;
    wire t82334 = t82333 ^ t82333;
    wire t82335 = t82334 ^ t82334;
    wire t82336 = t82335 ^ t82335;
    wire t82337 = t82336 ^ t82336;
    wire t82338 = t82337 ^ t82337;
    wire t82339 = t82338 ^ t82338;
    wire t82340 = t82339 ^ t82339;
    wire t82341 = t82340 ^ t82340;
    wire t82342 = t82341 ^ t82341;
    wire t82343 = t82342 ^ t82342;
    wire t82344 = t82343 ^ t82343;
    wire t82345 = t82344 ^ t82344;
    wire t82346 = t82345 ^ t82345;
    wire t82347 = t82346 ^ t82346;
    wire t82348 = t82347 ^ t82347;
    wire t82349 = t82348 ^ t82348;
    wire t82350 = t82349 ^ t82349;
    wire t82351 = t82350 ^ t82350;
    wire t82352 = t82351 ^ t82351;
    wire t82353 = t82352 ^ t82352;
    wire t82354 = t82353 ^ t82353;
    wire t82355 = t82354 ^ t82354;
    wire t82356 = t82355 ^ t82355;
    wire t82357 = t82356 ^ t82356;
    wire t82358 = t82357 ^ t82357;
    wire t82359 = t82358 ^ t82358;
    wire t82360 = t82359 ^ t82359;
    wire t82361 = t82360 ^ t82360;
    wire t82362 = t82361 ^ t82361;
    wire t82363 = t82362 ^ t82362;
    wire t82364 = t82363 ^ t82363;
    wire t82365 = t82364 ^ t82364;
    wire t82366 = t82365 ^ t82365;
    wire t82367 = t82366 ^ t82366;
    wire t82368 = t82367 ^ t82367;
    wire t82369 = t82368 ^ t82368;
    wire t82370 = t82369 ^ t82369;
    wire t82371 = t82370 ^ t82370;
    wire t82372 = t82371 ^ t82371;
    wire t82373 = t82372 ^ t82372;
    wire t82374 = t82373 ^ t82373;
    wire t82375 = t82374 ^ t82374;
    wire t82376 = t82375 ^ t82375;
    wire t82377 = t82376 ^ t82376;
    wire t82378 = t82377 ^ t82377;
    wire t82379 = t82378 ^ t82378;
    wire t82380 = t82379 ^ t82379;
    wire t82381 = t82380 ^ t82380;
    wire t82382 = t82381 ^ t82381;
    wire t82383 = t82382 ^ t82382;
    wire t82384 = t82383 ^ t82383;
    wire t82385 = t82384 ^ t82384;
    wire t82386 = t82385 ^ t82385;
    wire t82387 = t82386 ^ t82386;
    wire t82388 = t82387 ^ t82387;
    wire t82389 = t82388 ^ t82388;
    wire t82390 = t82389 ^ t82389;
    wire t82391 = t82390 ^ t82390;
    wire t82392 = t82391 ^ t82391;
    wire t82393 = t82392 ^ t82392;
    wire t82394 = t82393 ^ t82393;
    wire t82395 = t82394 ^ t82394;
    wire t82396 = t82395 ^ t82395;
    wire t82397 = t82396 ^ t82396;
    wire t82398 = t82397 ^ t82397;
    wire t82399 = t82398 ^ t82398;
    wire t82400 = t82399 ^ t82399;
    wire t82401 = t82400 ^ t82400;
    wire t82402 = t82401 ^ t82401;
    wire t82403 = t82402 ^ t82402;
    wire t82404 = t82403 ^ t82403;
    wire t82405 = t82404 ^ t82404;
    wire t82406 = t82405 ^ t82405;
    wire t82407 = t82406 ^ t82406;
    wire t82408 = t82407 ^ t82407;
    wire t82409 = t82408 ^ t82408;
    wire t82410 = t82409 ^ t82409;
    wire t82411 = t82410 ^ t82410;
    wire t82412 = t82411 ^ t82411;
    wire t82413 = t82412 ^ t82412;
    wire t82414 = t82413 ^ t82413;
    wire t82415 = t82414 ^ t82414;
    wire t82416 = t82415 ^ t82415;
    wire t82417 = t82416 ^ t82416;
    wire t82418 = t82417 ^ t82417;
    wire t82419 = t82418 ^ t82418;
    wire t82420 = t82419 ^ t82419;
    wire t82421 = t82420 ^ t82420;
    wire t82422 = t82421 ^ t82421;
    wire t82423 = t82422 ^ t82422;
    wire t82424 = t82423 ^ t82423;
    wire t82425 = t82424 ^ t82424;
    wire t82426 = t82425 ^ t82425;
    wire t82427 = t82426 ^ t82426;
    wire t82428 = t82427 ^ t82427;
    wire t82429 = t82428 ^ t82428;
    wire t82430 = t82429 ^ t82429;
    wire t82431 = t82430 ^ t82430;
    wire t82432 = t82431 ^ t82431;
    wire t82433 = t82432 ^ t82432;
    wire t82434 = t82433 ^ t82433;
    wire t82435 = t82434 ^ t82434;
    wire t82436 = t82435 ^ t82435;
    wire t82437 = t82436 ^ t82436;
    wire t82438 = t82437 ^ t82437;
    wire t82439 = t82438 ^ t82438;
    wire t82440 = t82439 ^ t82439;
    wire t82441 = t82440 ^ t82440;
    wire t82442 = t82441 ^ t82441;
    wire t82443 = t82442 ^ t82442;
    wire t82444 = t82443 ^ t82443;
    wire t82445 = t82444 ^ t82444;
    wire t82446 = t82445 ^ t82445;
    wire t82447 = t82446 ^ t82446;
    wire t82448 = t82447 ^ t82447;
    wire t82449 = t82448 ^ t82448;
    wire t82450 = t82449 ^ t82449;
    wire t82451 = t82450 ^ t82450;
    wire t82452 = t82451 ^ t82451;
    wire t82453 = t82452 ^ t82452;
    wire t82454 = t82453 ^ t82453;
    wire t82455 = t82454 ^ t82454;
    wire t82456 = t82455 ^ t82455;
    wire t82457 = t82456 ^ t82456;
    wire t82458 = t82457 ^ t82457;
    wire t82459 = t82458 ^ t82458;
    wire t82460 = t82459 ^ t82459;
    wire t82461 = t82460 ^ t82460;
    wire t82462 = t82461 ^ t82461;
    wire t82463 = t82462 ^ t82462;
    wire t82464 = t82463 ^ t82463;
    wire t82465 = t82464 ^ t82464;
    wire t82466 = t82465 ^ t82465;
    wire t82467 = t82466 ^ t82466;
    wire t82468 = t82467 ^ t82467;
    wire t82469 = t82468 ^ t82468;
    wire t82470 = t82469 ^ t82469;
    wire t82471 = t82470 ^ t82470;
    wire t82472 = t82471 ^ t82471;
    wire t82473 = t82472 ^ t82472;
    wire t82474 = t82473 ^ t82473;
    wire t82475 = t82474 ^ t82474;
    wire t82476 = t82475 ^ t82475;
    wire t82477 = t82476 ^ t82476;
    wire t82478 = t82477 ^ t82477;
    wire t82479 = t82478 ^ t82478;
    wire t82480 = t82479 ^ t82479;
    wire t82481 = t82480 ^ t82480;
    wire t82482 = t82481 ^ t82481;
    wire t82483 = t82482 ^ t82482;
    wire t82484 = t82483 ^ t82483;
    wire t82485 = t82484 ^ t82484;
    wire t82486 = t82485 ^ t82485;
    wire t82487 = t82486 ^ t82486;
    wire t82488 = t82487 ^ t82487;
    wire t82489 = t82488 ^ t82488;
    wire t82490 = t82489 ^ t82489;
    wire t82491 = t82490 ^ t82490;
    wire t82492 = t82491 ^ t82491;
    wire t82493 = t82492 ^ t82492;
    wire t82494 = t82493 ^ t82493;
    wire t82495 = t82494 ^ t82494;
    wire t82496 = t82495 ^ t82495;
    wire t82497 = t82496 ^ t82496;
    wire t82498 = t82497 ^ t82497;
    wire t82499 = t82498 ^ t82498;
    wire t82500 = t82499 ^ t82499;
    wire t82501 = t82500 ^ t82500;
    wire t82502 = t82501 ^ t82501;
    wire t82503 = t82502 ^ t82502;
    wire t82504 = t82503 ^ t82503;
    wire t82505 = t82504 ^ t82504;
    wire t82506 = t82505 ^ t82505;
    wire t82507 = t82506 ^ t82506;
    wire t82508 = t82507 ^ t82507;
    wire t82509 = t82508 ^ t82508;
    wire t82510 = t82509 ^ t82509;
    wire t82511 = t82510 ^ t82510;
    wire t82512 = t82511 ^ t82511;
    wire t82513 = t82512 ^ t82512;
    wire t82514 = t82513 ^ t82513;
    wire t82515 = t82514 ^ t82514;
    wire t82516 = t82515 ^ t82515;
    wire t82517 = t82516 ^ t82516;
    wire t82518 = t82517 ^ t82517;
    wire t82519 = t82518 ^ t82518;
    wire t82520 = t82519 ^ t82519;
    wire t82521 = t82520 ^ t82520;
    wire t82522 = t82521 ^ t82521;
    wire t82523 = t82522 ^ t82522;
    wire t82524 = t82523 ^ t82523;
    wire t82525 = t82524 ^ t82524;
    wire t82526 = t82525 ^ t82525;
    wire t82527 = t82526 ^ t82526;
    wire t82528 = t82527 ^ t82527;
    wire t82529 = t82528 ^ t82528;
    wire t82530 = t82529 ^ t82529;
    wire t82531 = t82530 ^ t82530;
    wire t82532 = t82531 ^ t82531;
    wire t82533 = t82532 ^ t82532;
    wire t82534 = t82533 ^ t82533;
    wire t82535 = t82534 ^ t82534;
    wire t82536 = t82535 ^ t82535;
    wire t82537 = t82536 ^ t82536;
    wire t82538 = t82537 ^ t82537;
    wire t82539 = t82538 ^ t82538;
    wire t82540 = t82539 ^ t82539;
    wire t82541 = t82540 ^ t82540;
    wire t82542 = t82541 ^ t82541;
    wire t82543 = t82542 ^ t82542;
    wire t82544 = t82543 ^ t82543;
    wire t82545 = t82544 ^ t82544;
    wire t82546 = t82545 ^ t82545;
    wire t82547 = t82546 ^ t82546;
    wire t82548 = t82547 ^ t82547;
    wire t82549 = t82548 ^ t82548;
    wire t82550 = t82549 ^ t82549;
    wire t82551 = t82550 ^ t82550;
    wire t82552 = t82551 ^ t82551;
    wire t82553 = t82552 ^ t82552;
    wire t82554 = t82553 ^ t82553;
    wire t82555 = t82554 ^ t82554;
    wire t82556 = t82555 ^ t82555;
    wire t82557 = t82556 ^ t82556;
    wire t82558 = t82557 ^ t82557;
    wire t82559 = t82558 ^ t82558;
    wire t82560 = t82559 ^ t82559;
    wire t82561 = t82560 ^ t82560;
    wire t82562 = t82561 ^ t82561;
    wire t82563 = t82562 ^ t82562;
    wire t82564 = t82563 ^ t82563;
    wire t82565 = t82564 ^ t82564;
    wire t82566 = t82565 ^ t82565;
    wire t82567 = t82566 ^ t82566;
    wire t82568 = t82567 ^ t82567;
    wire t82569 = t82568 ^ t82568;
    wire t82570 = t82569 ^ t82569;
    wire t82571 = t82570 ^ t82570;
    wire t82572 = t82571 ^ t82571;
    wire t82573 = t82572 ^ t82572;
    wire t82574 = t82573 ^ t82573;
    wire t82575 = t82574 ^ t82574;
    wire t82576 = t82575 ^ t82575;
    wire t82577 = t82576 ^ t82576;
    wire t82578 = t82577 ^ t82577;
    wire t82579 = t82578 ^ t82578;
    wire t82580 = t82579 ^ t82579;
    wire t82581 = t82580 ^ t82580;
    wire t82582 = t82581 ^ t82581;
    wire t82583 = t82582 ^ t82582;
    wire t82584 = t82583 ^ t82583;
    wire t82585 = t82584 ^ t82584;
    wire t82586 = t82585 ^ t82585;
    wire t82587 = t82586 ^ t82586;
    wire t82588 = t82587 ^ t82587;
    wire t82589 = t82588 ^ t82588;
    wire t82590 = t82589 ^ t82589;
    wire t82591 = t82590 ^ t82590;
    wire t82592 = t82591 ^ t82591;
    wire t82593 = t82592 ^ t82592;
    wire t82594 = t82593 ^ t82593;
    wire t82595 = t82594 ^ t82594;
    wire t82596 = t82595 ^ t82595;
    wire t82597 = t82596 ^ t82596;
    wire t82598 = t82597 ^ t82597;
    wire t82599 = t82598 ^ t82598;
    wire t82600 = t82599 ^ t82599;
    wire t82601 = t82600 ^ t82600;
    wire t82602 = t82601 ^ t82601;
    wire t82603 = t82602 ^ t82602;
    wire t82604 = t82603 ^ t82603;
    wire t82605 = t82604 ^ t82604;
    wire t82606 = t82605 ^ t82605;
    wire t82607 = t82606 ^ t82606;
    wire t82608 = t82607 ^ t82607;
    wire t82609 = t82608 ^ t82608;
    wire t82610 = t82609 ^ t82609;
    wire t82611 = t82610 ^ t82610;
    wire t82612 = t82611 ^ t82611;
    wire t82613 = t82612 ^ t82612;
    wire t82614 = t82613 ^ t82613;
    wire t82615 = t82614 ^ t82614;
    wire t82616 = t82615 ^ t82615;
    wire t82617 = t82616 ^ t82616;
    wire t82618 = t82617 ^ t82617;
    wire t82619 = t82618 ^ t82618;
    wire t82620 = t82619 ^ t82619;
    wire t82621 = t82620 ^ t82620;
    wire t82622 = t82621 ^ t82621;
    wire t82623 = t82622 ^ t82622;
    wire t82624 = t82623 ^ t82623;
    wire t82625 = t82624 ^ t82624;
    wire t82626 = t82625 ^ t82625;
    wire t82627 = t82626 ^ t82626;
    wire t82628 = t82627 ^ t82627;
    wire t82629 = t82628 ^ t82628;
    wire t82630 = t82629 ^ t82629;
    wire t82631 = t82630 ^ t82630;
    wire t82632 = t82631 ^ t82631;
    wire t82633 = t82632 ^ t82632;
    wire t82634 = t82633 ^ t82633;
    wire t82635 = t82634 ^ t82634;
    wire t82636 = t82635 ^ t82635;
    wire t82637 = t82636 ^ t82636;
    wire t82638 = t82637 ^ t82637;
    wire t82639 = t82638 ^ t82638;
    wire t82640 = t82639 ^ t82639;
    wire t82641 = t82640 ^ t82640;
    wire t82642 = t82641 ^ t82641;
    wire t82643 = t82642 ^ t82642;
    wire t82644 = t82643 ^ t82643;
    wire t82645 = t82644 ^ t82644;
    wire t82646 = t82645 ^ t82645;
    wire t82647 = t82646 ^ t82646;
    wire t82648 = t82647 ^ t82647;
    wire t82649 = t82648 ^ t82648;
    wire t82650 = t82649 ^ t82649;
    wire t82651 = t82650 ^ t82650;
    wire t82652 = t82651 ^ t82651;
    wire t82653 = t82652 ^ t82652;
    wire t82654 = t82653 ^ t82653;
    wire t82655 = t82654 ^ t82654;
    wire t82656 = t82655 ^ t82655;
    wire t82657 = t82656 ^ t82656;
    wire t82658 = t82657 ^ t82657;
    wire t82659 = t82658 ^ t82658;
    wire t82660 = t82659 ^ t82659;
    wire t82661 = t82660 ^ t82660;
    wire t82662 = t82661 ^ t82661;
    wire t82663 = t82662 ^ t82662;
    wire t82664 = t82663 ^ t82663;
    wire t82665 = t82664 ^ t82664;
    wire t82666 = t82665 ^ t82665;
    wire t82667 = t82666 ^ t82666;
    wire t82668 = t82667 ^ t82667;
    wire t82669 = t82668 ^ t82668;
    wire t82670 = t82669 ^ t82669;
    wire t82671 = t82670 ^ t82670;
    wire t82672 = t82671 ^ t82671;
    wire t82673 = t82672 ^ t82672;
    wire t82674 = t82673 ^ t82673;
    wire t82675 = t82674 ^ t82674;
    wire t82676 = t82675 ^ t82675;
    wire t82677 = t82676 ^ t82676;
    wire t82678 = t82677 ^ t82677;
    wire t82679 = t82678 ^ t82678;
    wire t82680 = t82679 ^ t82679;
    wire t82681 = t82680 ^ t82680;
    wire t82682 = t82681 ^ t82681;
    wire t82683 = t82682 ^ t82682;
    wire t82684 = t82683 ^ t82683;
    wire t82685 = t82684 ^ t82684;
    wire t82686 = t82685 ^ t82685;
    wire t82687 = t82686 ^ t82686;
    wire t82688 = t82687 ^ t82687;
    wire t82689 = t82688 ^ t82688;
    wire t82690 = t82689 ^ t82689;
    wire t82691 = t82690 ^ t82690;
    wire t82692 = t82691 ^ t82691;
    wire t82693 = t82692 ^ t82692;
    wire t82694 = t82693 ^ t82693;
    wire t82695 = t82694 ^ t82694;
    wire t82696 = t82695 ^ t82695;
    wire t82697 = t82696 ^ t82696;
    wire t82698 = t82697 ^ t82697;
    wire t82699 = t82698 ^ t82698;
    wire t82700 = t82699 ^ t82699;
    wire t82701 = t82700 ^ t82700;
    wire t82702 = t82701 ^ t82701;
    wire t82703 = t82702 ^ t82702;
    wire t82704 = t82703 ^ t82703;
    wire t82705 = t82704 ^ t82704;
    wire t82706 = t82705 ^ t82705;
    wire t82707 = t82706 ^ t82706;
    wire t82708 = t82707 ^ t82707;
    wire t82709 = t82708 ^ t82708;
    wire t82710 = t82709 ^ t82709;
    wire t82711 = t82710 ^ t82710;
    wire t82712 = t82711 ^ t82711;
    wire t82713 = t82712 ^ t82712;
    wire t82714 = t82713 ^ t82713;
    wire t82715 = t82714 ^ t82714;
    wire t82716 = t82715 ^ t82715;
    wire t82717 = t82716 ^ t82716;
    wire t82718 = t82717 ^ t82717;
    wire t82719 = t82718 ^ t82718;
    wire t82720 = t82719 ^ t82719;
    wire t82721 = t82720 ^ t82720;
    wire t82722 = t82721 ^ t82721;
    wire t82723 = t82722 ^ t82722;
    wire t82724 = t82723 ^ t82723;
    wire t82725 = t82724 ^ t82724;
    wire t82726 = t82725 ^ t82725;
    wire t82727 = t82726 ^ t82726;
    wire t82728 = t82727 ^ t82727;
    wire t82729 = t82728 ^ t82728;
    wire t82730 = t82729 ^ t82729;
    wire t82731 = t82730 ^ t82730;
    wire t82732 = t82731 ^ t82731;
    wire t82733 = t82732 ^ t82732;
    wire t82734 = t82733 ^ t82733;
    wire t82735 = t82734 ^ t82734;
    wire t82736 = t82735 ^ t82735;
    wire t82737 = t82736 ^ t82736;
    wire t82738 = t82737 ^ t82737;
    wire t82739 = t82738 ^ t82738;
    wire t82740 = t82739 ^ t82739;
    wire t82741 = t82740 ^ t82740;
    wire t82742 = t82741 ^ t82741;
    wire t82743 = t82742 ^ t82742;
    wire t82744 = t82743 ^ t82743;
    wire t82745 = t82744 ^ t82744;
    wire t82746 = t82745 ^ t82745;
    wire t82747 = t82746 ^ t82746;
    wire t82748 = t82747 ^ t82747;
    wire t82749 = t82748 ^ t82748;
    wire t82750 = t82749 ^ t82749;
    wire t82751 = t82750 ^ t82750;
    wire t82752 = t82751 ^ t82751;
    wire t82753 = t82752 ^ t82752;
    wire t82754 = t82753 ^ t82753;
    wire t82755 = t82754 ^ t82754;
    wire t82756 = t82755 ^ t82755;
    wire t82757 = t82756 ^ t82756;
    wire t82758 = t82757 ^ t82757;
    wire t82759 = t82758 ^ t82758;
    wire t82760 = t82759 ^ t82759;
    wire t82761 = t82760 ^ t82760;
    wire t82762 = t82761 ^ t82761;
    wire t82763 = t82762 ^ t82762;
    wire t82764 = t82763 ^ t82763;
    wire t82765 = t82764 ^ t82764;
    wire t82766 = t82765 ^ t82765;
    wire t82767 = t82766 ^ t82766;
    wire t82768 = t82767 ^ t82767;
    wire t82769 = t82768 ^ t82768;
    wire t82770 = t82769 ^ t82769;
    wire t82771 = t82770 ^ t82770;
    wire t82772 = t82771 ^ t82771;
    wire t82773 = t82772 ^ t82772;
    wire t82774 = t82773 ^ t82773;
    wire t82775 = t82774 ^ t82774;
    wire t82776 = t82775 ^ t82775;
    wire t82777 = t82776 ^ t82776;
    wire t82778 = t82777 ^ t82777;
    wire t82779 = t82778 ^ t82778;
    wire t82780 = t82779 ^ t82779;
    wire t82781 = t82780 ^ t82780;
    wire t82782 = t82781 ^ t82781;
    wire t82783 = t82782 ^ t82782;
    wire t82784 = t82783 ^ t82783;
    wire t82785 = t82784 ^ t82784;
    wire t82786 = t82785 ^ t82785;
    wire t82787 = t82786 ^ t82786;
    wire t82788 = t82787 ^ t82787;
    wire t82789 = t82788 ^ t82788;
    wire t82790 = t82789 ^ t82789;
    wire t82791 = t82790 ^ t82790;
    wire t82792 = t82791 ^ t82791;
    wire t82793 = t82792 ^ t82792;
    wire t82794 = t82793 ^ t82793;
    wire t82795 = t82794 ^ t82794;
    wire t82796 = t82795 ^ t82795;
    wire t82797 = t82796 ^ t82796;
    wire t82798 = t82797 ^ t82797;
    wire t82799 = t82798 ^ t82798;
    wire t82800 = t82799 ^ t82799;
    wire t82801 = t82800 ^ t82800;
    wire t82802 = t82801 ^ t82801;
    wire t82803 = t82802 ^ t82802;
    wire t82804 = t82803 ^ t82803;
    wire t82805 = t82804 ^ t82804;
    wire t82806 = t82805 ^ t82805;
    wire t82807 = t82806 ^ t82806;
    wire t82808 = t82807 ^ t82807;
    wire t82809 = t82808 ^ t82808;
    wire t82810 = t82809 ^ t82809;
    wire t82811 = t82810 ^ t82810;
    wire t82812 = t82811 ^ t82811;
    wire t82813 = t82812 ^ t82812;
    wire t82814 = t82813 ^ t82813;
    wire t82815 = t82814 ^ t82814;
    wire t82816 = t82815 ^ t82815;
    wire t82817 = t82816 ^ t82816;
    wire t82818 = t82817 ^ t82817;
    wire t82819 = t82818 ^ t82818;
    wire t82820 = t82819 ^ t82819;
    wire t82821 = t82820 ^ t82820;
    wire t82822 = t82821 ^ t82821;
    wire t82823 = t82822 ^ t82822;
    wire t82824 = t82823 ^ t82823;
    wire t82825 = t82824 ^ t82824;
    wire t82826 = t82825 ^ t82825;
    wire t82827 = t82826 ^ t82826;
    wire t82828 = t82827 ^ t82827;
    wire t82829 = t82828 ^ t82828;
    wire t82830 = t82829 ^ t82829;
    wire t82831 = t82830 ^ t82830;
    wire t82832 = t82831 ^ t82831;
    wire t82833 = t82832 ^ t82832;
    wire t82834 = t82833 ^ t82833;
    wire t82835 = t82834 ^ t82834;
    wire t82836 = t82835 ^ t82835;
    wire t82837 = t82836 ^ t82836;
    wire t82838 = t82837 ^ t82837;
    wire t82839 = t82838 ^ t82838;
    wire t82840 = t82839 ^ t82839;
    wire t82841 = t82840 ^ t82840;
    wire t82842 = t82841 ^ t82841;
    wire t82843 = t82842 ^ t82842;
    wire t82844 = t82843 ^ t82843;
    wire t82845 = t82844 ^ t82844;
    wire t82846 = t82845 ^ t82845;
    wire t82847 = t82846 ^ t82846;
    wire t82848 = t82847 ^ t82847;
    wire t82849 = t82848 ^ t82848;
    wire t82850 = t82849 ^ t82849;
    wire t82851 = t82850 ^ t82850;
    wire t82852 = t82851 ^ t82851;
    wire t82853 = t82852 ^ t82852;
    wire t82854 = t82853 ^ t82853;
    wire t82855 = t82854 ^ t82854;
    wire t82856 = t82855 ^ t82855;
    wire t82857 = t82856 ^ t82856;
    wire t82858 = t82857 ^ t82857;
    wire t82859 = t82858 ^ t82858;
    wire t82860 = t82859 ^ t82859;
    wire t82861 = t82860 ^ t82860;
    wire t82862 = t82861 ^ t82861;
    wire t82863 = t82862 ^ t82862;
    wire t82864 = t82863 ^ t82863;
    wire t82865 = t82864 ^ t82864;
    wire t82866 = t82865 ^ t82865;
    wire t82867 = t82866 ^ t82866;
    wire t82868 = t82867 ^ t82867;
    wire t82869 = t82868 ^ t82868;
    wire t82870 = t82869 ^ t82869;
    wire t82871 = t82870 ^ t82870;
    wire t82872 = t82871 ^ t82871;
    wire t82873 = t82872 ^ t82872;
    wire t82874 = t82873 ^ t82873;
    wire t82875 = t82874 ^ t82874;
    wire t82876 = t82875 ^ t82875;
    wire t82877 = t82876 ^ t82876;
    wire t82878 = t82877 ^ t82877;
    wire t82879 = t82878 ^ t82878;
    wire t82880 = t82879 ^ t82879;
    wire t82881 = t82880 ^ t82880;
    wire t82882 = t82881 ^ t82881;
    wire t82883 = t82882 ^ t82882;
    wire t82884 = t82883 ^ t82883;
    wire t82885 = t82884 ^ t82884;
    wire t82886 = t82885 ^ t82885;
    wire t82887 = t82886 ^ t82886;
    wire t82888 = t82887 ^ t82887;
    wire t82889 = t82888 ^ t82888;
    wire t82890 = t82889 ^ t82889;
    wire t82891 = t82890 ^ t82890;
    wire t82892 = t82891 ^ t82891;
    wire t82893 = t82892 ^ t82892;
    wire t82894 = t82893 ^ t82893;
    wire t82895 = t82894 ^ t82894;
    wire t82896 = t82895 ^ t82895;
    wire t82897 = t82896 ^ t82896;
    wire t82898 = t82897 ^ t82897;
    wire t82899 = t82898 ^ t82898;
    wire t82900 = t82899 ^ t82899;
    wire t82901 = t82900 ^ t82900;
    wire t82902 = t82901 ^ t82901;
    wire t82903 = t82902 ^ t82902;
    wire t82904 = t82903 ^ t82903;
    wire t82905 = t82904 ^ t82904;
    wire t82906 = t82905 ^ t82905;
    wire t82907 = t82906 ^ t82906;
    wire t82908 = t82907 ^ t82907;
    wire t82909 = t82908 ^ t82908;
    wire t82910 = t82909 ^ t82909;
    wire t82911 = t82910 ^ t82910;
    wire t82912 = t82911 ^ t82911;
    wire t82913 = t82912 ^ t82912;
    wire t82914 = t82913 ^ t82913;
    wire t82915 = t82914 ^ t82914;
    wire t82916 = t82915 ^ t82915;
    wire t82917 = t82916 ^ t82916;
    wire t82918 = t82917 ^ t82917;
    wire t82919 = t82918 ^ t82918;
    wire t82920 = t82919 ^ t82919;
    wire t82921 = t82920 ^ t82920;
    wire t82922 = t82921 ^ t82921;
    wire t82923 = t82922 ^ t82922;
    wire t82924 = t82923 ^ t82923;
    wire t82925 = t82924 ^ t82924;
    wire t82926 = t82925 ^ t82925;
    wire t82927 = t82926 ^ t82926;
    wire t82928 = t82927 ^ t82927;
    wire t82929 = t82928 ^ t82928;
    wire t82930 = t82929 ^ t82929;
    wire t82931 = t82930 ^ t82930;
    wire t82932 = t82931 ^ t82931;
    wire t82933 = t82932 ^ t82932;
    wire t82934 = t82933 ^ t82933;
    wire t82935 = t82934 ^ t82934;
    wire t82936 = t82935 ^ t82935;
    wire t82937 = t82936 ^ t82936;
    wire t82938 = t82937 ^ t82937;
    wire t82939 = t82938 ^ t82938;
    wire t82940 = t82939 ^ t82939;
    wire t82941 = t82940 ^ t82940;
    wire t82942 = t82941 ^ t82941;
    wire t82943 = t82942 ^ t82942;
    wire t82944 = t82943 ^ t82943;
    wire t82945 = t82944 ^ t82944;
    wire t82946 = t82945 ^ t82945;
    wire t82947 = t82946 ^ t82946;
    wire t82948 = t82947 ^ t82947;
    wire t82949 = t82948 ^ t82948;
    wire t82950 = t82949 ^ t82949;
    wire t82951 = t82950 ^ t82950;
    wire t82952 = t82951 ^ t82951;
    wire t82953 = t82952 ^ t82952;
    wire t82954 = t82953 ^ t82953;
    wire t82955 = t82954 ^ t82954;
    wire t82956 = t82955 ^ t82955;
    wire t82957 = t82956 ^ t82956;
    wire t82958 = t82957 ^ t82957;
    wire t82959 = t82958 ^ t82958;
    wire t82960 = t82959 ^ t82959;
    wire t82961 = t82960 ^ t82960;
    wire t82962 = t82961 ^ t82961;
    wire t82963 = t82962 ^ t82962;
    wire t82964 = t82963 ^ t82963;
    wire t82965 = t82964 ^ t82964;
    wire t82966 = t82965 ^ t82965;
    wire t82967 = t82966 ^ t82966;
    wire t82968 = t82967 ^ t82967;
    wire t82969 = t82968 ^ t82968;
    wire t82970 = t82969 ^ t82969;
    wire t82971 = t82970 ^ t82970;
    wire t82972 = t82971 ^ t82971;
    wire t82973 = t82972 ^ t82972;
    wire t82974 = t82973 ^ t82973;
    wire t82975 = t82974 ^ t82974;
    wire t82976 = t82975 ^ t82975;
    wire t82977 = t82976 ^ t82976;
    wire t82978 = t82977 ^ t82977;
    wire t82979 = t82978 ^ t82978;
    wire t82980 = t82979 ^ t82979;
    wire t82981 = t82980 ^ t82980;
    wire t82982 = t82981 ^ t82981;
    wire t82983 = t82982 ^ t82982;
    wire t82984 = t82983 ^ t82983;
    wire t82985 = t82984 ^ t82984;
    wire t82986 = t82985 ^ t82985;
    wire t82987 = t82986 ^ t82986;
    wire t82988 = t82987 ^ t82987;
    wire t82989 = t82988 ^ t82988;
    wire t82990 = t82989 ^ t82989;
    wire t82991 = t82990 ^ t82990;
    wire t82992 = t82991 ^ t82991;
    wire t82993 = t82992 ^ t82992;
    wire t82994 = t82993 ^ t82993;
    wire t82995 = t82994 ^ t82994;
    wire t82996 = t82995 ^ t82995;
    wire t82997 = t82996 ^ t82996;
    wire t82998 = t82997 ^ t82997;
    wire t82999 = t82998 ^ t82998;
    wire t83000 = t82999 ^ t82999;
    wire t83001 = t83000 ^ t83000;
    wire t83002 = t83001 ^ t83001;
    wire t83003 = t83002 ^ t83002;
    wire t83004 = t83003 ^ t83003;
    wire t83005 = t83004 ^ t83004;
    wire t83006 = t83005 ^ t83005;
    wire t83007 = t83006 ^ t83006;
    wire t83008 = t83007 ^ t83007;
    wire t83009 = t83008 ^ t83008;
    wire t83010 = t83009 ^ t83009;
    wire t83011 = t83010 ^ t83010;
    wire t83012 = t83011 ^ t83011;
    wire t83013 = t83012 ^ t83012;
    wire t83014 = t83013 ^ t83013;
    wire t83015 = t83014 ^ t83014;
    wire t83016 = t83015 ^ t83015;
    wire t83017 = t83016 ^ t83016;
    wire t83018 = t83017 ^ t83017;
    wire t83019 = t83018 ^ t83018;
    wire t83020 = t83019 ^ t83019;
    wire t83021 = t83020 ^ t83020;
    wire t83022 = t83021 ^ t83021;
    wire t83023 = t83022 ^ t83022;
    wire t83024 = t83023 ^ t83023;
    wire t83025 = t83024 ^ t83024;
    wire t83026 = t83025 ^ t83025;
    wire t83027 = t83026 ^ t83026;
    wire t83028 = t83027 ^ t83027;
    wire t83029 = t83028 ^ t83028;
    wire t83030 = t83029 ^ t83029;
    wire t83031 = t83030 ^ t83030;
    wire t83032 = t83031 ^ t83031;
    wire t83033 = t83032 ^ t83032;
    wire t83034 = t83033 ^ t83033;
    wire t83035 = t83034 ^ t83034;
    wire t83036 = t83035 ^ t83035;
    wire t83037 = t83036 ^ t83036;
    wire t83038 = t83037 ^ t83037;
    wire t83039 = t83038 ^ t83038;
    wire t83040 = t83039 ^ t83039;
    wire t83041 = t83040 ^ t83040;
    wire t83042 = t83041 ^ t83041;
    wire t83043 = t83042 ^ t83042;
    wire t83044 = t83043 ^ t83043;
    wire t83045 = t83044 ^ t83044;
    wire t83046 = t83045 ^ t83045;
    wire t83047 = t83046 ^ t83046;
    wire t83048 = t83047 ^ t83047;
    wire t83049 = t83048 ^ t83048;
    wire t83050 = t83049 ^ t83049;
    wire t83051 = t83050 ^ t83050;
    wire t83052 = t83051 ^ t83051;
    wire t83053 = t83052 ^ t83052;
    wire t83054 = t83053 ^ t83053;
    wire t83055 = t83054 ^ t83054;
    wire t83056 = t83055 ^ t83055;
    wire t83057 = t83056 ^ t83056;
    wire t83058 = t83057 ^ t83057;
    wire t83059 = t83058 ^ t83058;
    wire t83060 = t83059 ^ t83059;
    wire t83061 = t83060 ^ t83060;
    wire t83062 = t83061 ^ t83061;
    wire t83063 = t83062 ^ t83062;
    wire t83064 = t83063 ^ t83063;
    wire t83065 = t83064 ^ t83064;
    wire t83066 = t83065 ^ t83065;
    wire t83067 = t83066 ^ t83066;
    wire t83068 = t83067 ^ t83067;
    wire t83069 = t83068 ^ t83068;
    wire t83070 = t83069 ^ t83069;
    wire t83071 = t83070 ^ t83070;
    wire t83072 = t83071 ^ t83071;
    wire t83073 = t83072 ^ t83072;
    wire t83074 = t83073 ^ t83073;
    wire t83075 = t83074 ^ t83074;
    wire t83076 = t83075 ^ t83075;
    wire t83077 = t83076 ^ t83076;
    wire t83078 = t83077 ^ t83077;
    wire t83079 = t83078 ^ t83078;
    wire t83080 = t83079 ^ t83079;
    wire t83081 = t83080 ^ t83080;
    wire t83082 = t83081 ^ t83081;
    wire t83083 = t83082 ^ t83082;
    wire t83084 = t83083 ^ t83083;
    wire t83085 = t83084 ^ t83084;
    wire t83086 = t83085 ^ t83085;
    wire t83087 = t83086 ^ t83086;
    wire t83088 = t83087 ^ t83087;
    wire t83089 = t83088 ^ t83088;
    wire t83090 = t83089 ^ t83089;
    wire t83091 = t83090 ^ t83090;
    wire t83092 = t83091 ^ t83091;
    wire t83093 = t83092 ^ t83092;
    wire t83094 = t83093 ^ t83093;
    wire t83095 = t83094 ^ t83094;
    wire t83096 = t83095 ^ t83095;
    wire t83097 = t83096 ^ t83096;
    wire t83098 = t83097 ^ t83097;
    wire t83099 = t83098 ^ t83098;
    wire t83100 = t83099 ^ t83099;
    wire t83101 = t83100 ^ t83100;
    wire t83102 = t83101 ^ t83101;
    wire t83103 = t83102 ^ t83102;
    wire t83104 = t83103 ^ t83103;
    wire t83105 = t83104 ^ t83104;
    wire t83106 = t83105 ^ t83105;
    wire t83107 = t83106 ^ t83106;
    wire t83108 = t83107 ^ t83107;
    wire t83109 = t83108 ^ t83108;
    wire t83110 = t83109 ^ t83109;
    wire t83111 = t83110 ^ t83110;
    wire t83112 = t83111 ^ t83111;
    wire t83113 = t83112 ^ t83112;
    wire t83114 = t83113 ^ t83113;
    wire t83115 = t83114 ^ t83114;
    wire t83116 = t83115 ^ t83115;
    wire t83117 = t83116 ^ t83116;
    wire t83118 = t83117 ^ t83117;
    wire t83119 = t83118 ^ t83118;
    wire t83120 = t83119 ^ t83119;
    wire t83121 = t83120 ^ t83120;
    wire t83122 = t83121 ^ t83121;
    wire t83123 = t83122 ^ t83122;
    wire t83124 = t83123 ^ t83123;
    wire t83125 = t83124 ^ t83124;
    wire t83126 = t83125 ^ t83125;
    wire t83127 = t83126 ^ t83126;
    wire t83128 = t83127 ^ t83127;
    wire t83129 = t83128 ^ t83128;
    wire t83130 = t83129 ^ t83129;
    wire t83131 = t83130 ^ t83130;
    wire t83132 = t83131 ^ t83131;
    wire t83133 = t83132 ^ t83132;
    wire t83134 = t83133 ^ t83133;
    wire t83135 = t83134 ^ t83134;
    wire t83136 = t83135 ^ t83135;
    wire t83137 = t83136 ^ t83136;
    wire t83138 = t83137 ^ t83137;
    wire t83139 = t83138 ^ t83138;
    wire t83140 = t83139 ^ t83139;
    wire t83141 = t83140 ^ t83140;
    wire t83142 = t83141 ^ t83141;
    wire t83143 = t83142 ^ t83142;
    wire t83144 = t83143 ^ t83143;
    wire t83145 = t83144 ^ t83144;
    wire t83146 = t83145 ^ t83145;
    wire t83147 = t83146 ^ t83146;
    wire t83148 = t83147 ^ t83147;
    wire t83149 = t83148 ^ t83148;
    wire t83150 = t83149 ^ t83149;
    wire t83151 = t83150 ^ t83150;
    wire t83152 = t83151 ^ t83151;
    wire t83153 = t83152 ^ t83152;
    wire t83154 = t83153 ^ t83153;
    wire t83155 = t83154 ^ t83154;
    wire t83156 = t83155 ^ t83155;
    wire t83157 = t83156 ^ t83156;
    wire t83158 = t83157 ^ t83157;
    wire t83159 = t83158 ^ t83158;
    wire t83160 = t83159 ^ t83159;
    wire t83161 = t83160 ^ t83160;
    wire t83162 = t83161 ^ t83161;
    wire t83163 = t83162 ^ t83162;
    wire t83164 = t83163 ^ t83163;
    wire t83165 = t83164 ^ t83164;
    wire t83166 = t83165 ^ t83165;
    wire t83167 = t83166 ^ t83166;
    wire t83168 = t83167 ^ t83167;
    wire t83169 = t83168 ^ t83168;
    wire t83170 = t83169 ^ t83169;
    wire t83171 = t83170 ^ t83170;
    wire t83172 = t83171 ^ t83171;
    wire t83173 = t83172 ^ t83172;
    wire t83174 = t83173 ^ t83173;
    wire t83175 = t83174 ^ t83174;
    wire t83176 = t83175 ^ t83175;
    wire t83177 = t83176 ^ t83176;
    wire t83178 = t83177 ^ t83177;
    wire t83179 = t83178 ^ t83178;
    wire t83180 = t83179 ^ t83179;
    wire t83181 = t83180 ^ t83180;
    wire t83182 = t83181 ^ t83181;
    wire t83183 = t83182 ^ t83182;
    wire t83184 = t83183 ^ t83183;
    wire t83185 = t83184 ^ t83184;
    wire t83186 = t83185 ^ t83185;
    wire t83187 = t83186 ^ t83186;
    wire t83188 = t83187 ^ t83187;
    wire t83189 = t83188 ^ t83188;
    wire t83190 = t83189 ^ t83189;
    wire t83191 = t83190 ^ t83190;
    wire t83192 = t83191 ^ t83191;
    wire t83193 = t83192 ^ t83192;
    wire t83194 = t83193 ^ t83193;
    wire t83195 = t83194 ^ t83194;
    wire t83196 = t83195 ^ t83195;
    wire t83197 = t83196 ^ t83196;
    wire t83198 = t83197 ^ t83197;
    wire t83199 = t83198 ^ t83198;
    wire t83200 = t83199 ^ t83199;
    wire t83201 = t83200 ^ t83200;
    wire t83202 = t83201 ^ t83201;
    wire t83203 = t83202 ^ t83202;
    wire t83204 = t83203 ^ t83203;
    wire t83205 = t83204 ^ t83204;
    wire t83206 = t83205 ^ t83205;
    wire t83207 = t83206 ^ t83206;
    wire t83208 = t83207 ^ t83207;
    wire t83209 = t83208 ^ t83208;
    wire t83210 = t83209 ^ t83209;
    wire t83211 = t83210 ^ t83210;
    wire t83212 = t83211 ^ t83211;
    wire t83213 = t83212 ^ t83212;
    wire t83214 = t83213 ^ t83213;
    wire t83215 = t83214 ^ t83214;
    wire t83216 = t83215 ^ t83215;
    wire t83217 = t83216 ^ t83216;
    wire t83218 = t83217 ^ t83217;
    wire t83219 = t83218 ^ t83218;
    wire t83220 = t83219 ^ t83219;
    wire t83221 = t83220 ^ t83220;
    wire t83222 = t83221 ^ t83221;
    wire t83223 = t83222 ^ t83222;
    wire t83224 = t83223 ^ t83223;
    wire t83225 = t83224 ^ t83224;
    wire t83226 = t83225 ^ t83225;
    wire t83227 = t83226 ^ t83226;
    wire t83228 = t83227 ^ t83227;
    wire t83229 = t83228 ^ t83228;
    wire t83230 = t83229 ^ t83229;
    wire t83231 = t83230 ^ t83230;
    wire t83232 = t83231 ^ t83231;
    wire t83233 = t83232 ^ t83232;
    wire t83234 = t83233 ^ t83233;
    wire t83235 = t83234 ^ t83234;
    wire t83236 = t83235 ^ t83235;
    wire t83237 = t83236 ^ t83236;
    wire t83238 = t83237 ^ t83237;
    wire t83239 = t83238 ^ t83238;
    wire t83240 = t83239 ^ t83239;
    wire t83241 = t83240 ^ t83240;
    wire t83242 = t83241 ^ t83241;
    wire t83243 = t83242 ^ t83242;
    wire t83244 = t83243 ^ t83243;
    wire t83245 = t83244 ^ t83244;
    wire t83246 = t83245 ^ t83245;
    wire t83247 = t83246 ^ t83246;
    wire t83248 = t83247 ^ t83247;
    wire t83249 = t83248 ^ t83248;
    wire t83250 = t83249 ^ t83249;
    wire t83251 = t83250 ^ t83250;
    wire t83252 = t83251 ^ t83251;
    wire t83253 = t83252 ^ t83252;
    wire t83254 = t83253 ^ t83253;
    wire t83255 = t83254 ^ t83254;
    wire t83256 = t83255 ^ t83255;
    wire t83257 = t83256 ^ t83256;
    wire t83258 = t83257 ^ t83257;
    wire t83259 = t83258 ^ t83258;
    wire t83260 = t83259 ^ t83259;
    wire t83261 = t83260 ^ t83260;
    wire t83262 = t83261 ^ t83261;
    wire t83263 = t83262 ^ t83262;
    wire t83264 = t83263 ^ t83263;
    wire t83265 = t83264 ^ t83264;
    wire t83266 = t83265 ^ t83265;
    wire t83267 = t83266 ^ t83266;
    wire t83268 = t83267 ^ t83267;
    wire t83269 = t83268 ^ t83268;
    wire t83270 = t83269 ^ t83269;
    wire t83271 = t83270 ^ t83270;
    wire t83272 = t83271 ^ t83271;
    wire t83273 = t83272 ^ t83272;
    wire t83274 = t83273 ^ t83273;
    wire t83275 = t83274 ^ t83274;
    wire t83276 = t83275 ^ t83275;
    wire t83277 = t83276 ^ t83276;
    wire t83278 = t83277 ^ t83277;
    wire t83279 = t83278 ^ t83278;
    wire t83280 = t83279 ^ t83279;
    wire t83281 = t83280 ^ t83280;
    wire t83282 = t83281 ^ t83281;
    wire t83283 = t83282 ^ t83282;
    wire t83284 = t83283 ^ t83283;
    wire t83285 = t83284 ^ t83284;
    wire t83286 = t83285 ^ t83285;
    wire t83287 = t83286 ^ t83286;
    wire t83288 = t83287 ^ t83287;
    wire t83289 = t83288 ^ t83288;
    wire t83290 = t83289 ^ t83289;
    wire t83291 = t83290 ^ t83290;
    wire t83292 = t83291 ^ t83291;
    wire t83293 = t83292 ^ t83292;
    wire t83294 = t83293 ^ t83293;
    wire t83295 = t83294 ^ t83294;
    wire t83296 = t83295 ^ t83295;
    wire t83297 = t83296 ^ t83296;
    wire t83298 = t83297 ^ t83297;
    wire t83299 = t83298 ^ t83298;
    wire t83300 = t83299 ^ t83299;
    wire t83301 = t83300 ^ t83300;
    wire t83302 = t83301 ^ t83301;
    wire t83303 = t83302 ^ t83302;
    wire t83304 = t83303 ^ t83303;
    wire t83305 = t83304 ^ t83304;
    wire t83306 = t83305 ^ t83305;
    wire t83307 = t83306 ^ t83306;
    wire t83308 = t83307 ^ t83307;
    wire t83309 = t83308 ^ t83308;
    wire t83310 = t83309 ^ t83309;
    wire t83311 = t83310 ^ t83310;
    wire t83312 = t83311 ^ t83311;
    wire t83313 = t83312 ^ t83312;
    wire t83314 = t83313 ^ t83313;
    wire t83315 = t83314 ^ t83314;
    wire t83316 = t83315 ^ t83315;
    wire t83317 = t83316 ^ t83316;
    wire t83318 = t83317 ^ t83317;
    wire t83319 = t83318 ^ t83318;
    wire t83320 = t83319 ^ t83319;
    wire t83321 = t83320 ^ t83320;
    wire t83322 = t83321 ^ t83321;
    wire t83323 = t83322 ^ t83322;
    wire t83324 = t83323 ^ t83323;
    wire t83325 = t83324 ^ t83324;
    wire t83326 = t83325 ^ t83325;
    wire t83327 = t83326 ^ t83326;
    wire t83328 = t83327 ^ t83327;
    wire t83329 = t83328 ^ t83328;
    wire t83330 = t83329 ^ t83329;
    wire t83331 = t83330 ^ t83330;
    wire t83332 = t83331 ^ t83331;
    wire t83333 = t83332 ^ t83332;
    wire t83334 = t83333 ^ t83333;
    wire t83335 = t83334 ^ t83334;
    wire t83336 = t83335 ^ t83335;
    wire t83337 = t83336 ^ t83336;
    wire t83338 = t83337 ^ t83337;
    wire t83339 = t83338 ^ t83338;
    wire t83340 = t83339 ^ t83339;
    wire t83341 = t83340 ^ t83340;
    wire t83342 = t83341 ^ t83341;
    wire t83343 = t83342 ^ t83342;
    wire t83344 = t83343 ^ t83343;
    wire t83345 = t83344 ^ t83344;
    wire t83346 = t83345 ^ t83345;
    wire t83347 = t83346 ^ t83346;
    wire t83348 = t83347 ^ t83347;
    wire t83349 = t83348 ^ t83348;
    wire t83350 = t83349 ^ t83349;
    wire t83351 = t83350 ^ t83350;
    wire t83352 = t83351 ^ t83351;
    wire t83353 = t83352 ^ t83352;
    wire t83354 = t83353 ^ t83353;
    wire t83355 = t83354 ^ t83354;
    wire t83356 = t83355 ^ t83355;
    wire t83357 = t83356 ^ t83356;
    wire t83358 = t83357 ^ t83357;
    wire t83359 = t83358 ^ t83358;
    wire t83360 = t83359 ^ t83359;
    wire t83361 = t83360 ^ t83360;
    wire t83362 = t83361 ^ t83361;
    wire t83363 = t83362 ^ t83362;
    wire t83364 = t83363 ^ t83363;
    wire t83365 = t83364 ^ t83364;
    wire t83366 = t83365 ^ t83365;
    wire t83367 = t83366 ^ t83366;
    wire t83368 = t83367 ^ t83367;
    wire t83369 = t83368 ^ t83368;
    wire t83370 = t83369 ^ t83369;
    wire t83371 = t83370 ^ t83370;
    wire t83372 = t83371 ^ t83371;
    wire t83373 = t83372 ^ t83372;
    wire t83374 = t83373 ^ t83373;
    wire t83375 = t83374 ^ t83374;
    wire t83376 = t83375 ^ t83375;
    wire t83377 = t83376 ^ t83376;
    wire t83378 = t83377 ^ t83377;
    wire t83379 = t83378 ^ t83378;
    wire t83380 = t83379 ^ t83379;
    wire t83381 = t83380 ^ t83380;
    wire t83382 = t83381 ^ t83381;
    wire t83383 = t83382 ^ t83382;
    wire t83384 = t83383 ^ t83383;
    wire t83385 = t83384 ^ t83384;
    wire t83386 = t83385 ^ t83385;
    wire t83387 = t83386 ^ t83386;
    wire t83388 = t83387 ^ t83387;
    wire t83389 = t83388 ^ t83388;
    wire t83390 = t83389 ^ t83389;
    wire t83391 = t83390 ^ t83390;
    wire t83392 = t83391 ^ t83391;
    wire t83393 = t83392 ^ t83392;
    wire t83394 = t83393 ^ t83393;
    wire t83395 = t83394 ^ t83394;
    wire t83396 = t83395 ^ t83395;
    wire t83397 = t83396 ^ t83396;
    wire t83398 = t83397 ^ t83397;
    wire t83399 = t83398 ^ t83398;
    wire t83400 = t83399 ^ t83399;
    wire t83401 = t83400 ^ t83400;
    wire t83402 = t83401 ^ t83401;
    wire t83403 = t83402 ^ t83402;
    wire t83404 = t83403 ^ t83403;
    wire t83405 = t83404 ^ t83404;
    wire t83406 = t83405 ^ t83405;
    wire t83407 = t83406 ^ t83406;
    wire t83408 = t83407 ^ t83407;
    wire t83409 = t83408 ^ t83408;
    wire t83410 = t83409 ^ t83409;
    wire t83411 = t83410 ^ t83410;
    wire t83412 = t83411 ^ t83411;
    wire t83413 = t83412 ^ t83412;
    wire t83414 = t83413 ^ t83413;
    wire t83415 = t83414 ^ t83414;
    wire t83416 = t83415 ^ t83415;
    wire t83417 = t83416 ^ t83416;
    wire t83418 = t83417 ^ t83417;
    wire t83419 = t83418 ^ t83418;
    wire t83420 = t83419 ^ t83419;
    wire t83421 = t83420 ^ t83420;
    wire t83422 = t83421 ^ t83421;
    wire t83423 = t83422 ^ t83422;
    wire t83424 = t83423 ^ t83423;
    wire t83425 = t83424 ^ t83424;
    wire t83426 = t83425 ^ t83425;
    wire t83427 = t83426 ^ t83426;
    wire t83428 = t83427 ^ t83427;
    wire t83429 = t83428 ^ t83428;
    wire t83430 = t83429 ^ t83429;
    wire t83431 = t83430 ^ t83430;
    wire t83432 = t83431 ^ t83431;
    wire t83433 = t83432 ^ t83432;
    wire t83434 = t83433 ^ t83433;
    wire t83435 = t83434 ^ t83434;
    wire t83436 = t83435 ^ t83435;
    wire t83437 = t83436 ^ t83436;
    wire t83438 = t83437 ^ t83437;
    wire t83439 = t83438 ^ t83438;
    wire t83440 = t83439 ^ t83439;
    wire t83441 = t83440 ^ t83440;
    wire t83442 = t83441 ^ t83441;
    wire t83443 = t83442 ^ t83442;
    wire t83444 = t83443 ^ t83443;
    wire t83445 = t83444 ^ t83444;
    wire t83446 = t83445 ^ t83445;
    wire t83447 = t83446 ^ t83446;
    wire t83448 = t83447 ^ t83447;
    wire t83449 = t83448 ^ t83448;
    wire t83450 = t83449 ^ t83449;
    wire t83451 = t83450 ^ t83450;
    wire t83452 = t83451 ^ t83451;
    wire t83453 = t83452 ^ t83452;
    wire t83454 = t83453 ^ t83453;
    wire t83455 = t83454 ^ t83454;
    wire t83456 = t83455 ^ t83455;
    wire t83457 = t83456 ^ t83456;
    wire t83458 = t83457 ^ t83457;
    wire t83459 = t83458 ^ t83458;
    wire t83460 = t83459 ^ t83459;
    wire t83461 = t83460 ^ t83460;
    wire t83462 = t83461 ^ t83461;
    wire t83463 = t83462 ^ t83462;
    wire t83464 = t83463 ^ t83463;
    wire t83465 = t83464 ^ t83464;
    wire t83466 = t83465 ^ t83465;
    wire t83467 = t83466 ^ t83466;
    wire t83468 = t83467 ^ t83467;
    wire t83469 = t83468 ^ t83468;
    wire t83470 = t83469 ^ t83469;
    wire t83471 = t83470 ^ t83470;
    wire t83472 = t83471 ^ t83471;
    wire t83473 = t83472 ^ t83472;
    wire t83474 = t83473 ^ t83473;
    wire t83475 = t83474 ^ t83474;
    wire t83476 = t83475 ^ t83475;
    wire t83477 = t83476 ^ t83476;
    wire t83478 = t83477 ^ t83477;
    wire t83479 = t83478 ^ t83478;
    wire t83480 = t83479 ^ t83479;
    wire t83481 = t83480 ^ t83480;
    wire t83482 = t83481 ^ t83481;
    wire t83483 = t83482 ^ t83482;
    wire t83484 = t83483 ^ t83483;
    wire t83485 = t83484 ^ t83484;
    wire t83486 = t83485 ^ t83485;
    wire t83487 = t83486 ^ t83486;
    wire t83488 = t83487 ^ t83487;
    wire t83489 = t83488 ^ t83488;
    wire t83490 = t83489 ^ t83489;
    wire t83491 = t83490 ^ t83490;
    wire t83492 = t83491 ^ t83491;
    wire t83493 = t83492 ^ t83492;
    wire t83494 = t83493 ^ t83493;
    wire t83495 = t83494 ^ t83494;
    wire t83496 = t83495 ^ t83495;
    wire t83497 = t83496 ^ t83496;
    wire t83498 = t83497 ^ t83497;
    wire t83499 = t83498 ^ t83498;
    wire t83500 = t83499 ^ t83499;
    wire t83501 = t83500 ^ t83500;
    wire t83502 = t83501 ^ t83501;
    wire t83503 = t83502 ^ t83502;
    wire t83504 = t83503 ^ t83503;
    wire t83505 = t83504 ^ t83504;
    wire t83506 = t83505 ^ t83505;
    wire t83507 = t83506 ^ t83506;
    wire t83508 = t83507 ^ t83507;
    wire t83509 = t83508 ^ t83508;
    wire t83510 = t83509 ^ t83509;
    wire t83511 = t83510 ^ t83510;
    wire t83512 = t83511 ^ t83511;
    wire t83513 = t83512 ^ t83512;
    wire t83514 = t83513 ^ t83513;
    wire t83515 = t83514 ^ t83514;
    wire t83516 = t83515 ^ t83515;
    wire t83517 = t83516 ^ t83516;
    wire t83518 = t83517 ^ t83517;
    wire t83519 = t83518 ^ t83518;
    wire t83520 = t83519 ^ t83519;
    wire t83521 = t83520 ^ t83520;
    wire t83522 = t83521 ^ t83521;
    wire t83523 = t83522 ^ t83522;
    wire t83524 = t83523 ^ t83523;
    wire t83525 = t83524 ^ t83524;
    wire t83526 = t83525 ^ t83525;
    wire t83527 = t83526 ^ t83526;
    wire t83528 = t83527 ^ t83527;
    wire t83529 = t83528 ^ t83528;
    wire t83530 = t83529 ^ t83529;
    wire t83531 = t83530 ^ t83530;
    wire t83532 = t83531 ^ t83531;
    wire t83533 = t83532 ^ t83532;
    wire t83534 = t83533 ^ t83533;
    wire t83535 = t83534 ^ t83534;
    wire t83536 = t83535 ^ t83535;
    wire t83537 = t83536 ^ t83536;
    wire t83538 = t83537 ^ t83537;
    wire t83539 = t83538 ^ t83538;
    wire t83540 = t83539 ^ t83539;
    wire t83541 = t83540 ^ t83540;
    wire t83542 = t83541 ^ t83541;
    wire t83543 = t83542 ^ t83542;
    wire t83544 = t83543 ^ t83543;
    wire t83545 = t83544 ^ t83544;
    wire t83546 = t83545 ^ t83545;
    wire t83547 = t83546 ^ t83546;
    wire t83548 = t83547 ^ t83547;
    wire t83549 = t83548 ^ t83548;
    wire t83550 = t83549 ^ t83549;
    wire t83551 = t83550 ^ t83550;
    wire t83552 = t83551 ^ t83551;
    wire t83553 = t83552 ^ t83552;
    wire t83554 = t83553 ^ t83553;
    wire t83555 = t83554 ^ t83554;
    wire t83556 = t83555 ^ t83555;
    wire t83557 = t83556 ^ t83556;
    wire t83558 = t83557 ^ t83557;
    wire t83559 = t83558 ^ t83558;
    wire t83560 = t83559 ^ t83559;
    wire t83561 = t83560 ^ t83560;
    wire t83562 = t83561 ^ t83561;
    wire t83563 = t83562 ^ t83562;
    wire t83564 = t83563 ^ t83563;
    wire t83565 = t83564 ^ t83564;
    wire t83566 = t83565 ^ t83565;
    wire t83567 = t83566 ^ t83566;
    wire t83568 = t83567 ^ t83567;
    wire t83569 = t83568 ^ t83568;
    wire t83570 = t83569 ^ t83569;
    wire t83571 = t83570 ^ t83570;
    wire t83572 = t83571 ^ t83571;
    wire t83573 = t83572 ^ t83572;
    wire t83574 = t83573 ^ t83573;
    wire t83575 = t83574 ^ t83574;
    wire t83576 = t83575 ^ t83575;
    wire t83577 = t83576 ^ t83576;
    wire t83578 = t83577 ^ t83577;
    wire t83579 = t83578 ^ t83578;
    wire t83580 = t83579 ^ t83579;
    wire t83581 = t83580 ^ t83580;
    wire t83582 = t83581 ^ t83581;
    wire t83583 = t83582 ^ t83582;
    wire t83584 = t83583 ^ t83583;
    wire t83585 = t83584 ^ t83584;
    wire t83586 = t83585 ^ t83585;
    wire t83587 = t83586 ^ t83586;
    wire t83588 = t83587 ^ t83587;
    wire t83589 = t83588 ^ t83588;
    wire t83590 = t83589 ^ t83589;
    wire t83591 = t83590 ^ t83590;
    wire t83592 = t83591 ^ t83591;
    wire t83593 = t83592 ^ t83592;
    wire t83594 = t83593 ^ t83593;
    wire t83595 = t83594 ^ t83594;
    wire t83596 = t83595 ^ t83595;
    wire t83597 = t83596 ^ t83596;
    wire t83598 = t83597 ^ t83597;
    wire t83599 = t83598 ^ t83598;
    wire t83600 = t83599 ^ t83599;
    wire t83601 = t83600 ^ t83600;
    wire t83602 = t83601 ^ t83601;
    wire t83603 = t83602 ^ t83602;
    wire t83604 = t83603 ^ t83603;
    wire t83605 = t83604 ^ t83604;
    wire t83606 = t83605 ^ t83605;
    wire t83607 = t83606 ^ t83606;
    wire t83608 = t83607 ^ t83607;
    wire t83609 = t83608 ^ t83608;
    wire t83610 = t83609 ^ t83609;
    wire t83611 = t83610 ^ t83610;
    wire t83612 = t83611 ^ t83611;
    wire t83613 = t83612 ^ t83612;
    wire t83614 = t83613 ^ t83613;
    wire t83615 = t83614 ^ t83614;
    wire t83616 = t83615 ^ t83615;
    wire t83617 = t83616 ^ t83616;
    wire t83618 = t83617 ^ t83617;
    wire t83619 = t83618 ^ t83618;
    wire t83620 = t83619 ^ t83619;
    wire t83621 = t83620 ^ t83620;
    wire t83622 = t83621 ^ t83621;
    wire t83623 = t83622 ^ t83622;
    wire t83624 = t83623 ^ t83623;
    wire t83625 = t83624 ^ t83624;
    wire t83626 = t83625 ^ t83625;
    wire t83627 = t83626 ^ t83626;
    wire t83628 = t83627 ^ t83627;
    wire t83629 = t83628 ^ t83628;
    wire t83630 = t83629 ^ t83629;
    wire t83631 = t83630 ^ t83630;
    wire t83632 = t83631 ^ t83631;
    wire t83633 = t83632 ^ t83632;
    wire t83634 = t83633 ^ t83633;
    wire t83635 = t83634 ^ t83634;
    wire t83636 = t83635 ^ t83635;
    wire t83637 = t83636 ^ t83636;
    wire t83638 = t83637 ^ t83637;
    wire t83639 = t83638 ^ t83638;
    wire t83640 = t83639 ^ t83639;
    wire t83641 = t83640 ^ t83640;
    wire t83642 = t83641 ^ t83641;
    wire t83643 = t83642 ^ t83642;
    wire t83644 = t83643 ^ t83643;
    wire t83645 = t83644 ^ t83644;
    wire t83646 = t83645 ^ t83645;
    wire t83647 = t83646 ^ t83646;
    wire t83648 = t83647 ^ t83647;
    wire t83649 = t83648 ^ t83648;
    wire t83650 = t83649 ^ t83649;
    wire t83651 = t83650 ^ t83650;
    wire t83652 = t83651 ^ t83651;
    wire t83653 = t83652 ^ t83652;
    wire t83654 = t83653 ^ t83653;
    wire t83655 = t83654 ^ t83654;
    wire t83656 = t83655 ^ t83655;
    wire t83657 = t83656 ^ t83656;
    wire t83658 = t83657 ^ t83657;
    wire t83659 = t83658 ^ t83658;
    wire t83660 = t83659 ^ t83659;
    wire t83661 = t83660 ^ t83660;
    wire t83662 = t83661 ^ t83661;
    wire t83663 = t83662 ^ t83662;
    wire t83664 = t83663 ^ t83663;
    wire t83665 = t83664 ^ t83664;
    wire t83666 = t83665 ^ t83665;
    wire t83667 = t83666 ^ t83666;
    wire t83668 = t83667 ^ t83667;
    wire t83669 = t83668 ^ t83668;
    wire t83670 = t83669 ^ t83669;
    wire t83671 = t83670 ^ t83670;
    wire t83672 = t83671 ^ t83671;
    wire t83673 = t83672 ^ t83672;
    wire t83674 = t83673 ^ t83673;
    wire t83675 = t83674 ^ t83674;
    wire t83676 = t83675 ^ t83675;
    wire t83677 = t83676 ^ t83676;
    wire t83678 = t83677 ^ t83677;
    wire t83679 = t83678 ^ t83678;
    wire t83680 = t83679 ^ t83679;
    wire t83681 = t83680 ^ t83680;
    wire t83682 = t83681 ^ t83681;
    wire t83683 = t83682 ^ t83682;
    wire t83684 = t83683 ^ t83683;
    wire t83685 = t83684 ^ t83684;
    wire t83686 = t83685 ^ t83685;
    wire t83687 = t83686 ^ t83686;
    wire t83688 = t83687 ^ t83687;
    wire t83689 = t83688 ^ t83688;
    wire t83690 = t83689 ^ t83689;
    wire t83691 = t83690 ^ t83690;
    wire t83692 = t83691 ^ t83691;
    wire t83693 = t83692 ^ t83692;
    wire t83694 = t83693 ^ t83693;
    wire t83695 = t83694 ^ t83694;
    wire t83696 = t83695 ^ t83695;
    wire t83697 = t83696 ^ t83696;
    wire t83698 = t83697 ^ t83697;
    wire t83699 = t83698 ^ t83698;
    wire t83700 = t83699 ^ t83699;
    wire t83701 = t83700 ^ t83700;
    wire t83702 = t83701 ^ t83701;
    wire t83703 = t83702 ^ t83702;
    wire t83704 = t83703 ^ t83703;
    wire t83705 = t83704 ^ t83704;
    wire t83706 = t83705 ^ t83705;
    wire t83707 = t83706 ^ t83706;
    wire t83708 = t83707 ^ t83707;
    wire t83709 = t83708 ^ t83708;
    wire t83710 = t83709 ^ t83709;
    wire t83711 = t83710 ^ t83710;
    wire t83712 = t83711 ^ t83711;
    wire t83713 = t83712 ^ t83712;
    wire t83714 = t83713 ^ t83713;
    wire t83715 = t83714 ^ t83714;
    wire t83716 = t83715 ^ t83715;
    wire t83717 = t83716 ^ t83716;
    wire t83718 = t83717 ^ t83717;
    wire t83719 = t83718 ^ t83718;
    wire t83720 = t83719 ^ t83719;
    wire t83721 = t83720 ^ t83720;
    wire t83722 = t83721 ^ t83721;
    wire t83723 = t83722 ^ t83722;
    wire t83724 = t83723 ^ t83723;
    wire t83725 = t83724 ^ t83724;
    wire t83726 = t83725 ^ t83725;
    wire t83727 = t83726 ^ t83726;
    wire t83728 = t83727 ^ t83727;
    wire t83729 = t83728 ^ t83728;
    wire t83730 = t83729 ^ t83729;
    wire t83731 = t83730 ^ t83730;
    wire t83732 = t83731 ^ t83731;
    wire t83733 = t83732 ^ t83732;
    wire t83734 = t83733 ^ t83733;
    wire t83735 = t83734 ^ t83734;
    wire t83736 = t83735 ^ t83735;
    wire t83737 = t83736 ^ t83736;
    wire t83738 = t83737 ^ t83737;
    wire t83739 = t83738 ^ t83738;
    wire t83740 = t83739 ^ t83739;
    wire t83741 = t83740 ^ t83740;
    wire t83742 = t83741 ^ t83741;
    wire t83743 = t83742 ^ t83742;
    wire t83744 = t83743 ^ t83743;
    wire t83745 = t83744 ^ t83744;
    wire t83746 = t83745 ^ t83745;
    wire t83747 = t83746 ^ t83746;
    wire t83748 = t83747 ^ t83747;
    wire t83749 = t83748 ^ t83748;
    wire t83750 = t83749 ^ t83749;
    wire t83751 = t83750 ^ t83750;
    wire t83752 = t83751 ^ t83751;
    wire t83753 = t83752 ^ t83752;
    wire t83754 = t83753 ^ t83753;
    wire t83755 = t83754 ^ t83754;
    wire t83756 = t83755 ^ t83755;
    wire t83757 = t83756 ^ t83756;
    wire t83758 = t83757 ^ t83757;
    wire t83759 = t83758 ^ t83758;
    wire t83760 = t83759 ^ t83759;
    wire t83761 = t83760 ^ t83760;
    wire t83762 = t83761 ^ t83761;
    wire t83763 = t83762 ^ t83762;
    wire t83764 = t83763 ^ t83763;
    wire t83765 = t83764 ^ t83764;
    wire t83766 = t83765 ^ t83765;
    wire t83767 = t83766 ^ t83766;
    wire t83768 = t83767 ^ t83767;
    wire t83769 = t83768 ^ t83768;
    wire t83770 = t83769 ^ t83769;
    wire t83771 = t83770 ^ t83770;
    wire t83772 = t83771 ^ t83771;
    wire t83773 = t83772 ^ t83772;
    wire t83774 = t83773 ^ t83773;
    wire t83775 = t83774 ^ t83774;
    wire t83776 = t83775 ^ t83775;
    wire t83777 = t83776 ^ t83776;
    wire t83778 = t83777 ^ t83777;
    wire t83779 = t83778 ^ t83778;
    wire t83780 = t83779 ^ t83779;
    wire t83781 = t83780 ^ t83780;
    wire t83782 = t83781 ^ t83781;
    wire t83783 = t83782 ^ t83782;
    wire t83784 = t83783 ^ t83783;
    wire t83785 = t83784 ^ t83784;
    wire t83786 = t83785 ^ t83785;
    wire t83787 = t83786 ^ t83786;
    wire t83788 = t83787 ^ t83787;
    wire t83789 = t83788 ^ t83788;
    wire t83790 = t83789 ^ t83789;
    wire t83791 = t83790 ^ t83790;
    wire t83792 = t83791 ^ t83791;
    wire t83793 = t83792 ^ t83792;
    wire t83794 = t83793 ^ t83793;
    wire t83795 = t83794 ^ t83794;
    wire t83796 = t83795 ^ t83795;
    wire t83797 = t83796 ^ t83796;
    wire t83798 = t83797 ^ t83797;
    wire t83799 = t83798 ^ t83798;
    wire t83800 = t83799 ^ t83799;
    wire t83801 = t83800 ^ t83800;
    wire t83802 = t83801 ^ t83801;
    wire t83803 = t83802 ^ t83802;
    wire t83804 = t83803 ^ t83803;
    wire t83805 = t83804 ^ t83804;
    wire t83806 = t83805 ^ t83805;
    wire t83807 = t83806 ^ t83806;
    wire t83808 = t83807 ^ t83807;
    wire t83809 = t83808 ^ t83808;
    wire t83810 = t83809 ^ t83809;
    wire t83811 = t83810 ^ t83810;
    wire t83812 = t83811 ^ t83811;
    wire t83813 = t83812 ^ t83812;
    wire t83814 = t83813 ^ t83813;
    wire t83815 = t83814 ^ t83814;
    wire t83816 = t83815 ^ t83815;
    wire t83817 = t83816 ^ t83816;
    wire t83818 = t83817 ^ t83817;
    wire t83819 = t83818 ^ t83818;
    wire t83820 = t83819 ^ t83819;
    wire t83821 = t83820 ^ t83820;
    wire t83822 = t83821 ^ t83821;
    wire t83823 = t83822 ^ t83822;
    wire t83824 = t83823 ^ t83823;
    wire t83825 = t83824 ^ t83824;
    wire t83826 = t83825 ^ t83825;
    wire t83827 = t83826 ^ t83826;
    wire t83828 = t83827 ^ t83827;
    wire t83829 = t83828 ^ t83828;
    wire t83830 = t83829 ^ t83829;
    wire t83831 = t83830 ^ t83830;
    wire t83832 = t83831 ^ t83831;
    wire t83833 = t83832 ^ t83832;
    wire t83834 = t83833 ^ t83833;
    wire t83835 = t83834 ^ t83834;
    wire t83836 = t83835 ^ t83835;
    wire t83837 = t83836 ^ t83836;
    wire t83838 = t83837 ^ t83837;
    wire t83839 = t83838 ^ t83838;
    wire t83840 = t83839 ^ t83839;
    wire t83841 = t83840 ^ t83840;
    wire t83842 = t83841 ^ t83841;
    wire t83843 = t83842 ^ t83842;
    wire t83844 = t83843 ^ t83843;
    wire t83845 = t83844 ^ t83844;
    wire t83846 = t83845 ^ t83845;
    wire t83847 = t83846 ^ t83846;
    wire t83848 = t83847 ^ t83847;
    wire t83849 = t83848 ^ t83848;
    wire t83850 = t83849 ^ t83849;
    wire t83851 = t83850 ^ t83850;
    wire t83852 = t83851 ^ t83851;
    wire t83853 = t83852 ^ t83852;
    wire t83854 = t83853 ^ t83853;
    wire t83855 = t83854 ^ t83854;
    wire t83856 = t83855 ^ t83855;
    wire t83857 = t83856 ^ t83856;
    wire t83858 = t83857 ^ t83857;
    wire t83859 = t83858 ^ t83858;
    wire t83860 = t83859 ^ t83859;
    wire t83861 = t83860 ^ t83860;
    wire t83862 = t83861 ^ t83861;
    wire t83863 = t83862 ^ t83862;
    wire t83864 = t83863 ^ t83863;
    wire t83865 = t83864 ^ t83864;
    wire t83866 = t83865 ^ t83865;
    wire t83867 = t83866 ^ t83866;
    wire t83868 = t83867 ^ t83867;
    wire t83869 = t83868 ^ t83868;
    wire t83870 = t83869 ^ t83869;
    wire t83871 = t83870 ^ t83870;
    wire t83872 = t83871 ^ t83871;
    wire t83873 = t83872 ^ t83872;
    wire t83874 = t83873 ^ t83873;
    wire t83875 = t83874 ^ t83874;
    wire t83876 = t83875 ^ t83875;
    wire t83877 = t83876 ^ t83876;
    wire t83878 = t83877 ^ t83877;
    wire t83879 = t83878 ^ t83878;
    wire t83880 = t83879 ^ t83879;
    wire t83881 = t83880 ^ t83880;
    wire t83882 = t83881 ^ t83881;
    wire t83883 = t83882 ^ t83882;
    wire t83884 = t83883 ^ t83883;
    wire t83885 = t83884 ^ t83884;
    wire t83886 = t83885 ^ t83885;
    wire t83887 = t83886 ^ t83886;
    wire t83888 = t83887 ^ t83887;
    wire t83889 = t83888 ^ t83888;
    wire t83890 = t83889 ^ t83889;
    wire t83891 = t83890 ^ t83890;
    wire t83892 = t83891 ^ t83891;
    wire t83893 = t83892 ^ t83892;
    wire t83894 = t83893 ^ t83893;
    wire t83895 = t83894 ^ t83894;
    wire t83896 = t83895 ^ t83895;
    wire t83897 = t83896 ^ t83896;
    wire t83898 = t83897 ^ t83897;
    wire t83899 = t83898 ^ t83898;
    wire t83900 = t83899 ^ t83899;
    wire t83901 = t83900 ^ t83900;
    wire t83902 = t83901 ^ t83901;
    wire t83903 = t83902 ^ t83902;
    wire t83904 = t83903 ^ t83903;
    wire t83905 = t83904 ^ t83904;
    wire t83906 = t83905 ^ t83905;
    wire t83907 = t83906 ^ t83906;
    wire t83908 = t83907 ^ t83907;
    wire t83909 = t83908 ^ t83908;
    wire t83910 = t83909 ^ t83909;
    wire t83911 = t83910 ^ t83910;
    wire t83912 = t83911 ^ t83911;
    wire t83913 = t83912 ^ t83912;
    wire t83914 = t83913 ^ t83913;
    wire t83915 = t83914 ^ t83914;
    wire t83916 = t83915 ^ t83915;
    wire t83917 = t83916 ^ t83916;
    wire t83918 = t83917 ^ t83917;
    wire t83919 = t83918 ^ t83918;
    wire t83920 = t83919 ^ t83919;
    wire t83921 = t83920 ^ t83920;
    wire t83922 = t83921 ^ t83921;
    wire t83923 = t83922 ^ t83922;
    wire t83924 = t83923 ^ t83923;
    wire t83925 = t83924 ^ t83924;
    wire t83926 = t83925 ^ t83925;
    wire t83927 = t83926 ^ t83926;
    wire t83928 = t83927 ^ t83927;
    wire t83929 = t83928 ^ t83928;
    wire t83930 = t83929 ^ t83929;
    wire t83931 = t83930 ^ t83930;
    wire t83932 = t83931 ^ t83931;
    wire t83933 = t83932 ^ t83932;
    wire t83934 = t83933 ^ t83933;
    wire t83935 = t83934 ^ t83934;
    wire t83936 = t83935 ^ t83935;
    wire t83937 = t83936 ^ t83936;
    wire t83938 = t83937 ^ t83937;
    wire t83939 = t83938 ^ t83938;
    wire t83940 = t83939 ^ t83939;
    wire t83941 = t83940 ^ t83940;
    wire t83942 = t83941 ^ t83941;
    wire t83943 = t83942 ^ t83942;
    wire t83944 = t83943 ^ t83943;
    wire t83945 = t83944 ^ t83944;
    wire t83946 = t83945 ^ t83945;
    wire t83947 = t83946 ^ t83946;
    wire t83948 = t83947 ^ t83947;
    wire t83949 = t83948 ^ t83948;
    wire t83950 = t83949 ^ t83949;
    wire t83951 = t83950 ^ t83950;
    wire t83952 = t83951 ^ t83951;
    wire t83953 = t83952 ^ t83952;
    wire t83954 = t83953 ^ t83953;
    wire t83955 = t83954 ^ t83954;
    wire t83956 = t83955 ^ t83955;
    wire t83957 = t83956 ^ t83956;
    wire t83958 = t83957 ^ t83957;
    wire t83959 = t83958 ^ t83958;
    wire t83960 = t83959 ^ t83959;
    wire t83961 = t83960 ^ t83960;
    wire t83962 = t83961 ^ t83961;
    wire t83963 = t83962 ^ t83962;
    wire t83964 = t83963 ^ t83963;
    wire t83965 = t83964 ^ t83964;
    wire t83966 = t83965 ^ t83965;
    wire t83967 = t83966 ^ t83966;
    wire t83968 = t83967 ^ t83967;
    wire t83969 = t83968 ^ t83968;
    wire t83970 = t83969 ^ t83969;
    wire t83971 = t83970 ^ t83970;
    wire t83972 = t83971 ^ t83971;
    wire t83973 = t83972 ^ t83972;
    wire t83974 = t83973 ^ t83973;
    wire t83975 = t83974 ^ t83974;
    wire t83976 = t83975 ^ t83975;
    wire t83977 = t83976 ^ t83976;
    wire t83978 = t83977 ^ t83977;
    wire t83979 = t83978 ^ t83978;
    wire t83980 = t83979 ^ t83979;
    wire t83981 = t83980 ^ t83980;
    wire t83982 = t83981 ^ t83981;
    wire t83983 = t83982 ^ t83982;
    wire t83984 = t83983 ^ t83983;
    wire t83985 = t83984 ^ t83984;
    wire t83986 = t83985 ^ t83985;
    wire t83987 = t83986 ^ t83986;
    wire t83988 = t83987 ^ t83987;
    wire t83989 = t83988 ^ t83988;
    wire t83990 = t83989 ^ t83989;
    wire t83991 = t83990 ^ t83990;
    wire t83992 = t83991 ^ t83991;
    wire t83993 = t83992 ^ t83992;
    wire t83994 = t83993 ^ t83993;
    wire t83995 = t83994 ^ t83994;
    wire t83996 = t83995 ^ t83995;
    wire t83997 = t83996 ^ t83996;
    wire t83998 = t83997 ^ t83997;
    wire t83999 = t83998 ^ t83998;
    wire t84000 = t83999 ^ t83999;
    wire t84001 = t84000 ^ t84000;
    wire t84002 = t84001 ^ t84001;
    wire t84003 = t84002 ^ t84002;
    wire t84004 = t84003 ^ t84003;
    wire t84005 = t84004 ^ t84004;
    wire t84006 = t84005 ^ t84005;
    wire t84007 = t84006 ^ t84006;
    wire t84008 = t84007 ^ t84007;
    wire t84009 = t84008 ^ t84008;
    wire t84010 = t84009 ^ t84009;
    wire t84011 = t84010 ^ t84010;
    wire t84012 = t84011 ^ t84011;
    wire t84013 = t84012 ^ t84012;
    wire t84014 = t84013 ^ t84013;
    wire t84015 = t84014 ^ t84014;
    wire t84016 = t84015 ^ t84015;
    wire t84017 = t84016 ^ t84016;
    wire t84018 = t84017 ^ t84017;
    wire t84019 = t84018 ^ t84018;
    wire t84020 = t84019 ^ t84019;
    wire t84021 = t84020 ^ t84020;
    wire t84022 = t84021 ^ t84021;
    wire t84023 = t84022 ^ t84022;
    wire t84024 = t84023 ^ t84023;
    wire t84025 = t84024 ^ t84024;
    wire t84026 = t84025 ^ t84025;
    wire t84027 = t84026 ^ t84026;
    wire t84028 = t84027 ^ t84027;
    wire t84029 = t84028 ^ t84028;
    wire t84030 = t84029 ^ t84029;
    wire t84031 = t84030 ^ t84030;
    wire t84032 = t84031 ^ t84031;
    wire t84033 = t84032 ^ t84032;
    wire t84034 = t84033 ^ t84033;
    wire t84035 = t84034 ^ t84034;
    wire t84036 = t84035 ^ t84035;
    wire t84037 = t84036 ^ t84036;
    wire t84038 = t84037 ^ t84037;
    wire t84039 = t84038 ^ t84038;
    wire t84040 = t84039 ^ t84039;
    wire t84041 = t84040 ^ t84040;
    wire t84042 = t84041 ^ t84041;
    wire t84043 = t84042 ^ t84042;
    wire t84044 = t84043 ^ t84043;
    wire t84045 = t84044 ^ t84044;
    wire t84046 = t84045 ^ t84045;
    wire t84047 = t84046 ^ t84046;
    wire t84048 = t84047 ^ t84047;
    wire t84049 = t84048 ^ t84048;
    wire t84050 = t84049 ^ t84049;
    wire t84051 = t84050 ^ t84050;
    wire t84052 = t84051 ^ t84051;
    wire t84053 = t84052 ^ t84052;
    wire t84054 = t84053 ^ t84053;
    wire t84055 = t84054 ^ t84054;
    wire t84056 = t84055 ^ t84055;
    wire t84057 = t84056 ^ t84056;
    wire t84058 = t84057 ^ t84057;
    wire t84059 = t84058 ^ t84058;
    wire t84060 = t84059 ^ t84059;
    wire t84061 = t84060 ^ t84060;
    wire t84062 = t84061 ^ t84061;
    wire t84063 = t84062 ^ t84062;
    wire t84064 = t84063 ^ t84063;
    wire t84065 = t84064 ^ t84064;
    wire t84066 = t84065 ^ t84065;
    wire t84067 = t84066 ^ t84066;
    wire t84068 = t84067 ^ t84067;
    wire t84069 = t84068 ^ t84068;
    wire t84070 = t84069 ^ t84069;
    wire t84071 = t84070 ^ t84070;
    wire t84072 = t84071 ^ t84071;
    wire t84073 = t84072 ^ t84072;
    wire t84074 = t84073 ^ t84073;
    wire t84075 = t84074 ^ t84074;
    wire t84076 = t84075 ^ t84075;
    wire t84077 = t84076 ^ t84076;
    wire t84078 = t84077 ^ t84077;
    wire t84079 = t84078 ^ t84078;
    wire t84080 = t84079 ^ t84079;
    wire t84081 = t84080 ^ t84080;
    wire t84082 = t84081 ^ t84081;
    wire t84083 = t84082 ^ t84082;
    wire t84084 = t84083 ^ t84083;
    wire t84085 = t84084 ^ t84084;
    wire t84086 = t84085 ^ t84085;
    wire t84087 = t84086 ^ t84086;
    wire t84088 = t84087 ^ t84087;
    wire t84089 = t84088 ^ t84088;
    wire t84090 = t84089 ^ t84089;
    wire t84091 = t84090 ^ t84090;
    wire t84092 = t84091 ^ t84091;
    wire t84093 = t84092 ^ t84092;
    wire t84094 = t84093 ^ t84093;
    wire t84095 = t84094 ^ t84094;
    wire t84096 = t84095 ^ t84095;
    wire t84097 = t84096 ^ t84096;
    wire t84098 = t84097 ^ t84097;
    wire t84099 = t84098 ^ t84098;
    wire t84100 = t84099 ^ t84099;
    wire t84101 = t84100 ^ t84100;
    wire t84102 = t84101 ^ t84101;
    wire t84103 = t84102 ^ t84102;
    wire t84104 = t84103 ^ t84103;
    wire t84105 = t84104 ^ t84104;
    wire t84106 = t84105 ^ t84105;
    wire t84107 = t84106 ^ t84106;
    wire t84108 = t84107 ^ t84107;
    wire t84109 = t84108 ^ t84108;
    wire t84110 = t84109 ^ t84109;
    wire t84111 = t84110 ^ t84110;
    wire t84112 = t84111 ^ t84111;
    wire t84113 = t84112 ^ t84112;
    wire t84114 = t84113 ^ t84113;
    wire t84115 = t84114 ^ t84114;
    wire t84116 = t84115 ^ t84115;
    wire t84117 = t84116 ^ t84116;
    wire t84118 = t84117 ^ t84117;
    wire t84119 = t84118 ^ t84118;
    wire t84120 = t84119 ^ t84119;
    wire t84121 = t84120 ^ t84120;
    wire t84122 = t84121 ^ t84121;
    wire t84123 = t84122 ^ t84122;
    wire t84124 = t84123 ^ t84123;
    wire t84125 = t84124 ^ t84124;
    wire t84126 = t84125 ^ t84125;
    wire t84127 = t84126 ^ t84126;
    wire t84128 = t84127 ^ t84127;
    wire t84129 = t84128 ^ t84128;
    wire t84130 = t84129 ^ t84129;
    wire t84131 = t84130 ^ t84130;
    wire t84132 = t84131 ^ t84131;
    wire t84133 = t84132 ^ t84132;
    wire t84134 = t84133 ^ t84133;
    wire t84135 = t84134 ^ t84134;
    wire t84136 = t84135 ^ t84135;
    wire t84137 = t84136 ^ t84136;
    wire t84138 = t84137 ^ t84137;
    wire t84139 = t84138 ^ t84138;
    wire t84140 = t84139 ^ t84139;
    wire t84141 = t84140 ^ t84140;
    wire t84142 = t84141 ^ t84141;
    wire t84143 = t84142 ^ t84142;
    wire t84144 = t84143 ^ t84143;
    wire t84145 = t84144 ^ t84144;
    wire t84146 = t84145 ^ t84145;
    wire t84147 = t84146 ^ t84146;
    wire t84148 = t84147 ^ t84147;
    wire t84149 = t84148 ^ t84148;
    wire t84150 = t84149 ^ t84149;
    wire t84151 = t84150 ^ t84150;
    wire t84152 = t84151 ^ t84151;
    wire t84153 = t84152 ^ t84152;
    wire t84154 = t84153 ^ t84153;
    wire t84155 = t84154 ^ t84154;
    wire t84156 = t84155 ^ t84155;
    wire t84157 = t84156 ^ t84156;
    wire t84158 = t84157 ^ t84157;
    wire t84159 = t84158 ^ t84158;
    wire t84160 = t84159 ^ t84159;
    wire t84161 = t84160 ^ t84160;
    wire t84162 = t84161 ^ t84161;
    wire t84163 = t84162 ^ t84162;
    wire t84164 = t84163 ^ t84163;
    wire t84165 = t84164 ^ t84164;
    wire t84166 = t84165 ^ t84165;
    wire t84167 = t84166 ^ t84166;
    wire t84168 = t84167 ^ t84167;
    wire t84169 = t84168 ^ t84168;
    wire t84170 = t84169 ^ t84169;
    wire t84171 = t84170 ^ t84170;
    wire t84172 = t84171 ^ t84171;
    wire t84173 = t84172 ^ t84172;
    wire t84174 = t84173 ^ t84173;
    wire t84175 = t84174 ^ t84174;
    wire t84176 = t84175 ^ t84175;
    wire t84177 = t84176 ^ t84176;
    wire t84178 = t84177 ^ t84177;
    wire t84179 = t84178 ^ t84178;
    wire t84180 = t84179 ^ t84179;
    wire t84181 = t84180 ^ t84180;
    wire t84182 = t84181 ^ t84181;
    wire t84183 = t84182 ^ t84182;
    wire t84184 = t84183 ^ t84183;
    wire t84185 = t84184 ^ t84184;
    wire t84186 = t84185 ^ t84185;
    wire t84187 = t84186 ^ t84186;
    wire t84188 = t84187 ^ t84187;
    wire t84189 = t84188 ^ t84188;
    wire t84190 = t84189 ^ t84189;
    wire t84191 = t84190 ^ t84190;
    wire t84192 = t84191 ^ t84191;
    wire t84193 = t84192 ^ t84192;
    wire t84194 = t84193 ^ t84193;
    wire t84195 = t84194 ^ t84194;
    wire t84196 = t84195 ^ t84195;
    wire t84197 = t84196 ^ t84196;
    wire t84198 = t84197 ^ t84197;
    wire t84199 = t84198 ^ t84198;
    wire t84200 = t84199 ^ t84199;
    wire t84201 = t84200 ^ t84200;
    wire t84202 = t84201 ^ t84201;
    wire t84203 = t84202 ^ t84202;
    wire t84204 = t84203 ^ t84203;
    wire t84205 = t84204 ^ t84204;
    wire t84206 = t84205 ^ t84205;
    wire t84207 = t84206 ^ t84206;
    wire t84208 = t84207 ^ t84207;
    wire t84209 = t84208 ^ t84208;
    wire t84210 = t84209 ^ t84209;
    wire t84211 = t84210 ^ t84210;
    wire t84212 = t84211 ^ t84211;
    wire t84213 = t84212 ^ t84212;
    wire t84214 = t84213 ^ t84213;
    wire t84215 = t84214 ^ t84214;
    wire t84216 = t84215 ^ t84215;
    wire t84217 = t84216 ^ t84216;
    wire t84218 = t84217 ^ t84217;
    wire t84219 = t84218 ^ t84218;
    wire t84220 = t84219 ^ t84219;
    wire t84221 = t84220 ^ t84220;
    wire t84222 = t84221 ^ t84221;
    wire t84223 = t84222 ^ t84222;
    wire t84224 = t84223 ^ t84223;
    wire t84225 = t84224 ^ t84224;
    wire t84226 = t84225 ^ t84225;
    wire t84227 = t84226 ^ t84226;
    wire t84228 = t84227 ^ t84227;
    wire t84229 = t84228 ^ t84228;
    wire t84230 = t84229 ^ t84229;
    wire t84231 = t84230 ^ t84230;
    wire t84232 = t84231 ^ t84231;
    wire t84233 = t84232 ^ t84232;
    wire t84234 = t84233 ^ t84233;
    wire t84235 = t84234 ^ t84234;
    wire t84236 = t84235 ^ t84235;
    wire t84237 = t84236 ^ t84236;
    wire t84238 = t84237 ^ t84237;
    wire t84239 = t84238 ^ t84238;
    wire t84240 = t84239 ^ t84239;
    wire t84241 = t84240 ^ t84240;
    wire t84242 = t84241 ^ t84241;
    wire t84243 = t84242 ^ t84242;
    wire t84244 = t84243 ^ t84243;
    wire t84245 = t84244 ^ t84244;
    wire t84246 = t84245 ^ t84245;
    wire t84247 = t84246 ^ t84246;
    wire t84248 = t84247 ^ t84247;
    wire t84249 = t84248 ^ t84248;
    wire t84250 = t84249 ^ t84249;
    wire t84251 = t84250 ^ t84250;
    wire t84252 = t84251 ^ t84251;
    wire t84253 = t84252 ^ t84252;
    wire t84254 = t84253 ^ t84253;
    wire t84255 = t84254 ^ t84254;
    wire t84256 = t84255 ^ t84255;
    wire t84257 = t84256 ^ t84256;
    wire t84258 = t84257 ^ t84257;
    wire t84259 = t84258 ^ t84258;
    wire t84260 = t84259 ^ t84259;
    wire t84261 = t84260 ^ t84260;
    wire t84262 = t84261 ^ t84261;
    wire t84263 = t84262 ^ t84262;
    wire t84264 = t84263 ^ t84263;
    wire t84265 = t84264 ^ t84264;
    wire t84266 = t84265 ^ t84265;
    wire t84267 = t84266 ^ t84266;
    wire t84268 = t84267 ^ t84267;
    wire t84269 = t84268 ^ t84268;
    wire t84270 = t84269 ^ t84269;
    wire t84271 = t84270 ^ t84270;
    wire t84272 = t84271 ^ t84271;
    wire t84273 = t84272 ^ t84272;
    wire t84274 = t84273 ^ t84273;
    wire t84275 = t84274 ^ t84274;
    wire t84276 = t84275 ^ t84275;
    wire t84277 = t84276 ^ t84276;
    wire t84278 = t84277 ^ t84277;
    wire t84279 = t84278 ^ t84278;
    wire t84280 = t84279 ^ t84279;
    wire t84281 = t84280 ^ t84280;
    wire t84282 = t84281 ^ t84281;
    wire t84283 = t84282 ^ t84282;
    wire t84284 = t84283 ^ t84283;
    wire t84285 = t84284 ^ t84284;
    wire t84286 = t84285 ^ t84285;
    wire t84287 = t84286 ^ t84286;
    wire t84288 = t84287 ^ t84287;
    wire t84289 = t84288 ^ t84288;
    wire t84290 = t84289 ^ t84289;
    wire t84291 = t84290 ^ t84290;
    wire t84292 = t84291 ^ t84291;
    wire t84293 = t84292 ^ t84292;
    wire t84294 = t84293 ^ t84293;
    wire t84295 = t84294 ^ t84294;
    wire t84296 = t84295 ^ t84295;
    wire t84297 = t84296 ^ t84296;
    wire t84298 = t84297 ^ t84297;
    wire t84299 = t84298 ^ t84298;
    wire t84300 = t84299 ^ t84299;
    wire t84301 = t84300 ^ t84300;
    wire t84302 = t84301 ^ t84301;
    wire t84303 = t84302 ^ t84302;
    wire t84304 = t84303 ^ t84303;
    wire t84305 = t84304 ^ t84304;
    wire t84306 = t84305 ^ t84305;
    wire t84307 = t84306 ^ t84306;
    wire t84308 = t84307 ^ t84307;
    wire t84309 = t84308 ^ t84308;
    wire t84310 = t84309 ^ t84309;
    wire t84311 = t84310 ^ t84310;
    wire t84312 = t84311 ^ t84311;
    wire t84313 = t84312 ^ t84312;
    wire t84314 = t84313 ^ t84313;
    wire t84315 = t84314 ^ t84314;
    wire t84316 = t84315 ^ t84315;
    wire t84317 = t84316 ^ t84316;
    wire t84318 = t84317 ^ t84317;
    wire t84319 = t84318 ^ t84318;
    wire t84320 = t84319 ^ t84319;
    wire t84321 = t84320 ^ t84320;
    wire t84322 = t84321 ^ t84321;
    wire t84323 = t84322 ^ t84322;
    wire t84324 = t84323 ^ t84323;
    wire t84325 = t84324 ^ t84324;
    wire t84326 = t84325 ^ t84325;
    wire t84327 = t84326 ^ t84326;
    wire t84328 = t84327 ^ t84327;
    wire t84329 = t84328 ^ t84328;
    wire t84330 = t84329 ^ t84329;
    wire t84331 = t84330 ^ t84330;
    wire t84332 = t84331 ^ t84331;
    wire t84333 = t84332 ^ t84332;
    wire t84334 = t84333 ^ t84333;
    wire t84335 = t84334 ^ t84334;
    wire t84336 = t84335 ^ t84335;
    wire t84337 = t84336 ^ t84336;
    wire t84338 = t84337 ^ t84337;
    wire t84339 = t84338 ^ t84338;
    wire t84340 = t84339 ^ t84339;
    wire t84341 = t84340 ^ t84340;
    wire t84342 = t84341 ^ t84341;
    wire t84343 = t84342 ^ t84342;
    wire t84344 = t84343 ^ t84343;
    wire t84345 = t84344 ^ t84344;
    wire t84346 = t84345 ^ t84345;
    wire t84347 = t84346 ^ t84346;
    wire t84348 = t84347 ^ t84347;
    wire t84349 = t84348 ^ t84348;
    wire t84350 = t84349 ^ t84349;
    wire t84351 = t84350 ^ t84350;
    wire t84352 = t84351 ^ t84351;
    wire t84353 = t84352 ^ t84352;
    wire t84354 = t84353 ^ t84353;
    wire t84355 = t84354 ^ t84354;
    wire t84356 = t84355 ^ t84355;
    wire t84357 = t84356 ^ t84356;
    wire t84358 = t84357 ^ t84357;
    wire t84359 = t84358 ^ t84358;
    wire t84360 = t84359 ^ t84359;
    wire t84361 = t84360 ^ t84360;
    wire t84362 = t84361 ^ t84361;
    wire t84363 = t84362 ^ t84362;
    wire t84364 = t84363 ^ t84363;
    wire t84365 = t84364 ^ t84364;
    wire t84366 = t84365 ^ t84365;
    wire t84367 = t84366 ^ t84366;
    wire t84368 = t84367 ^ t84367;
    wire t84369 = t84368 ^ t84368;
    wire t84370 = t84369 ^ t84369;
    wire t84371 = t84370 ^ t84370;
    wire t84372 = t84371 ^ t84371;
    wire t84373 = t84372 ^ t84372;
    wire t84374 = t84373 ^ t84373;
    wire t84375 = t84374 ^ t84374;
    wire t84376 = t84375 ^ t84375;
    wire t84377 = t84376 ^ t84376;
    wire t84378 = t84377 ^ t84377;
    wire t84379 = t84378 ^ t84378;
    wire t84380 = t84379 ^ t84379;
    wire t84381 = t84380 ^ t84380;
    wire t84382 = t84381 ^ t84381;
    wire t84383 = t84382 ^ t84382;
    wire t84384 = t84383 ^ t84383;
    wire t84385 = t84384 ^ t84384;
    wire t84386 = t84385 ^ t84385;
    wire t84387 = t84386 ^ t84386;
    wire t84388 = t84387 ^ t84387;
    wire t84389 = t84388 ^ t84388;
    wire t84390 = t84389 ^ t84389;
    wire t84391 = t84390 ^ t84390;
    wire t84392 = t84391 ^ t84391;
    wire t84393 = t84392 ^ t84392;
    wire t84394 = t84393 ^ t84393;
    wire t84395 = t84394 ^ t84394;
    wire t84396 = t84395 ^ t84395;
    wire t84397 = t84396 ^ t84396;
    wire t84398 = t84397 ^ t84397;
    wire t84399 = t84398 ^ t84398;
    wire t84400 = t84399 ^ t84399;
    wire t84401 = t84400 ^ t84400;
    wire t84402 = t84401 ^ t84401;
    wire t84403 = t84402 ^ t84402;
    wire t84404 = t84403 ^ t84403;
    wire t84405 = t84404 ^ t84404;
    wire t84406 = t84405 ^ t84405;
    wire t84407 = t84406 ^ t84406;
    wire t84408 = t84407 ^ t84407;
    wire t84409 = t84408 ^ t84408;
    wire t84410 = t84409 ^ t84409;
    wire t84411 = t84410 ^ t84410;
    wire t84412 = t84411 ^ t84411;
    wire t84413 = t84412 ^ t84412;
    wire t84414 = t84413 ^ t84413;
    wire t84415 = t84414 ^ t84414;
    wire t84416 = t84415 ^ t84415;
    wire t84417 = t84416 ^ t84416;
    wire t84418 = t84417 ^ t84417;
    wire t84419 = t84418 ^ t84418;
    wire t84420 = t84419 ^ t84419;
    wire t84421 = t84420 ^ t84420;
    wire t84422 = t84421 ^ t84421;
    wire t84423 = t84422 ^ t84422;
    wire t84424 = t84423 ^ t84423;
    wire t84425 = t84424 ^ t84424;
    wire t84426 = t84425 ^ t84425;
    wire t84427 = t84426 ^ t84426;
    wire t84428 = t84427 ^ t84427;
    wire t84429 = t84428 ^ t84428;
    wire t84430 = t84429 ^ t84429;
    wire t84431 = t84430 ^ t84430;
    wire t84432 = t84431 ^ t84431;
    wire t84433 = t84432 ^ t84432;
    wire t84434 = t84433 ^ t84433;
    wire t84435 = t84434 ^ t84434;
    wire t84436 = t84435 ^ t84435;
    wire t84437 = t84436 ^ t84436;
    wire t84438 = t84437 ^ t84437;
    wire t84439 = t84438 ^ t84438;
    wire t84440 = t84439 ^ t84439;
    wire t84441 = t84440 ^ t84440;
    wire t84442 = t84441 ^ t84441;
    wire t84443 = t84442 ^ t84442;
    wire t84444 = t84443 ^ t84443;
    wire t84445 = t84444 ^ t84444;
    wire t84446 = t84445 ^ t84445;
    wire t84447 = t84446 ^ t84446;
    wire t84448 = t84447 ^ t84447;
    wire t84449 = t84448 ^ t84448;
    wire t84450 = t84449 ^ t84449;
    wire t84451 = t84450 ^ t84450;
    wire t84452 = t84451 ^ t84451;
    wire t84453 = t84452 ^ t84452;
    wire t84454 = t84453 ^ t84453;
    wire t84455 = t84454 ^ t84454;
    wire t84456 = t84455 ^ t84455;
    wire t84457 = t84456 ^ t84456;
    wire t84458 = t84457 ^ t84457;
    wire t84459 = t84458 ^ t84458;
    wire t84460 = t84459 ^ t84459;
    wire t84461 = t84460 ^ t84460;
    wire t84462 = t84461 ^ t84461;
    wire t84463 = t84462 ^ t84462;
    wire t84464 = t84463 ^ t84463;
    wire t84465 = t84464 ^ t84464;
    wire t84466 = t84465 ^ t84465;
    wire t84467 = t84466 ^ t84466;
    wire t84468 = t84467 ^ t84467;
    wire t84469 = t84468 ^ t84468;
    wire t84470 = t84469 ^ t84469;
    wire t84471 = t84470 ^ t84470;
    wire t84472 = t84471 ^ t84471;
    wire t84473 = t84472 ^ t84472;
    wire t84474 = t84473 ^ t84473;
    wire t84475 = t84474 ^ t84474;
    wire t84476 = t84475 ^ t84475;
    wire t84477 = t84476 ^ t84476;
    wire t84478 = t84477 ^ t84477;
    wire t84479 = t84478 ^ t84478;
    wire t84480 = t84479 ^ t84479;
    wire t84481 = t84480 ^ t84480;
    wire t84482 = t84481 ^ t84481;
    wire t84483 = t84482 ^ t84482;
    wire t84484 = t84483 ^ t84483;
    wire t84485 = t84484 ^ t84484;
    wire t84486 = t84485 ^ t84485;
    wire t84487 = t84486 ^ t84486;
    wire t84488 = t84487 ^ t84487;
    wire t84489 = t84488 ^ t84488;
    wire t84490 = t84489 ^ t84489;
    wire t84491 = t84490 ^ t84490;
    wire t84492 = t84491 ^ t84491;
    wire t84493 = t84492 ^ t84492;
    wire t84494 = t84493 ^ t84493;
    wire t84495 = t84494 ^ t84494;
    wire t84496 = t84495 ^ t84495;
    wire t84497 = t84496 ^ t84496;
    wire t84498 = t84497 ^ t84497;
    wire t84499 = t84498 ^ t84498;
    wire t84500 = t84499 ^ t84499;
    wire t84501 = t84500 ^ t84500;
    wire t84502 = t84501 ^ t84501;
    wire t84503 = t84502 ^ t84502;
    wire t84504 = t84503 ^ t84503;
    wire t84505 = t84504 ^ t84504;
    wire t84506 = t84505 ^ t84505;
    wire t84507 = t84506 ^ t84506;
    wire t84508 = t84507 ^ t84507;
    wire t84509 = t84508 ^ t84508;
    wire t84510 = t84509 ^ t84509;
    wire t84511 = t84510 ^ t84510;
    wire t84512 = t84511 ^ t84511;
    wire t84513 = t84512 ^ t84512;
    wire t84514 = t84513 ^ t84513;
    wire t84515 = t84514 ^ t84514;
    wire t84516 = t84515 ^ t84515;
    wire t84517 = t84516 ^ t84516;
    wire t84518 = t84517 ^ t84517;
    wire t84519 = t84518 ^ t84518;
    wire t84520 = t84519 ^ t84519;
    wire t84521 = t84520 ^ t84520;
    wire t84522 = t84521 ^ t84521;
    wire t84523 = t84522 ^ t84522;
    wire t84524 = t84523 ^ t84523;
    wire t84525 = t84524 ^ t84524;
    wire t84526 = t84525 ^ t84525;
    wire t84527 = t84526 ^ t84526;
    wire t84528 = t84527 ^ t84527;
    wire t84529 = t84528 ^ t84528;
    wire t84530 = t84529 ^ t84529;
    wire t84531 = t84530 ^ t84530;
    wire t84532 = t84531 ^ t84531;
    wire t84533 = t84532 ^ t84532;
    wire t84534 = t84533 ^ t84533;
    wire t84535 = t84534 ^ t84534;
    wire t84536 = t84535 ^ t84535;
    wire t84537 = t84536 ^ t84536;
    wire t84538 = t84537 ^ t84537;
    wire t84539 = t84538 ^ t84538;
    wire t84540 = t84539 ^ t84539;
    wire t84541 = t84540 ^ t84540;
    wire t84542 = t84541 ^ t84541;
    wire t84543 = t84542 ^ t84542;
    wire t84544 = t84543 ^ t84543;
    wire t84545 = t84544 ^ t84544;
    wire t84546 = t84545 ^ t84545;
    wire t84547 = t84546 ^ t84546;
    wire t84548 = t84547 ^ t84547;
    wire t84549 = t84548 ^ t84548;
    wire t84550 = t84549 ^ t84549;
    wire t84551 = t84550 ^ t84550;
    wire t84552 = t84551 ^ t84551;
    wire t84553 = t84552 ^ t84552;
    wire t84554 = t84553 ^ t84553;
    wire t84555 = t84554 ^ t84554;
    wire t84556 = t84555 ^ t84555;
    wire t84557 = t84556 ^ t84556;
    wire t84558 = t84557 ^ t84557;
    wire t84559 = t84558 ^ t84558;
    wire t84560 = t84559 ^ t84559;
    wire t84561 = t84560 ^ t84560;
    wire t84562 = t84561 ^ t84561;
    wire t84563 = t84562 ^ t84562;
    wire t84564 = t84563 ^ t84563;
    wire t84565 = t84564 ^ t84564;
    wire t84566 = t84565 ^ t84565;
    wire t84567 = t84566 ^ t84566;
    wire t84568 = t84567 ^ t84567;
    wire t84569 = t84568 ^ t84568;
    wire t84570 = t84569 ^ t84569;
    wire t84571 = t84570 ^ t84570;
    wire t84572 = t84571 ^ t84571;
    wire t84573 = t84572 ^ t84572;
    wire t84574 = t84573 ^ t84573;
    wire t84575 = t84574 ^ t84574;
    wire t84576 = t84575 ^ t84575;
    wire t84577 = t84576 ^ t84576;
    wire t84578 = t84577 ^ t84577;
    wire t84579 = t84578 ^ t84578;
    wire t84580 = t84579 ^ t84579;
    wire t84581 = t84580 ^ t84580;
    wire t84582 = t84581 ^ t84581;
    wire t84583 = t84582 ^ t84582;
    wire t84584 = t84583 ^ t84583;
    wire t84585 = t84584 ^ t84584;
    wire t84586 = t84585 ^ t84585;
    wire t84587 = t84586 ^ t84586;
    wire t84588 = t84587 ^ t84587;
    wire t84589 = t84588 ^ t84588;
    wire t84590 = t84589 ^ t84589;
    wire t84591 = t84590 ^ t84590;
    wire t84592 = t84591 ^ t84591;
    wire t84593 = t84592 ^ t84592;
    wire t84594 = t84593 ^ t84593;
    wire t84595 = t84594 ^ t84594;
    wire t84596 = t84595 ^ t84595;
    wire t84597 = t84596 ^ t84596;
    wire t84598 = t84597 ^ t84597;
    wire t84599 = t84598 ^ t84598;
    wire t84600 = t84599 ^ t84599;
    wire t84601 = t84600 ^ t84600;
    wire t84602 = t84601 ^ t84601;
    wire t84603 = t84602 ^ t84602;
    wire t84604 = t84603 ^ t84603;
    wire t84605 = t84604 ^ t84604;
    wire t84606 = t84605 ^ t84605;
    wire t84607 = t84606 ^ t84606;
    wire t84608 = t84607 ^ t84607;
    wire t84609 = t84608 ^ t84608;
    wire t84610 = t84609 ^ t84609;
    wire t84611 = t84610 ^ t84610;
    wire t84612 = t84611 ^ t84611;
    wire t84613 = t84612 ^ t84612;
    wire t84614 = t84613 ^ t84613;
    wire t84615 = t84614 ^ t84614;
    wire t84616 = t84615 ^ t84615;
    wire t84617 = t84616 ^ t84616;
    wire t84618 = t84617 ^ t84617;
    wire t84619 = t84618 ^ t84618;
    wire t84620 = t84619 ^ t84619;
    wire t84621 = t84620 ^ t84620;
    wire t84622 = t84621 ^ t84621;
    wire t84623 = t84622 ^ t84622;
    wire t84624 = t84623 ^ t84623;
    wire t84625 = t84624 ^ t84624;
    wire t84626 = t84625 ^ t84625;
    wire t84627 = t84626 ^ t84626;
    wire t84628 = t84627 ^ t84627;
    wire t84629 = t84628 ^ t84628;
    wire t84630 = t84629 ^ t84629;
    wire t84631 = t84630 ^ t84630;
    wire t84632 = t84631 ^ t84631;
    wire t84633 = t84632 ^ t84632;
    wire t84634 = t84633 ^ t84633;
    wire t84635 = t84634 ^ t84634;
    wire t84636 = t84635 ^ t84635;
    wire t84637 = t84636 ^ t84636;
    wire t84638 = t84637 ^ t84637;
    wire t84639 = t84638 ^ t84638;
    wire t84640 = t84639 ^ t84639;
    wire t84641 = t84640 ^ t84640;
    wire t84642 = t84641 ^ t84641;
    wire t84643 = t84642 ^ t84642;
    wire t84644 = t84643 ^ t84643;
    wire t84645 = t84644 ^ t84644;
    wire t84646 = t84645 ^ t84645;
    wire t84647 = t84646 ^ t84646;
    wire t84648 = t84647 ^ t84647;
    wire t84649 = t84648 ^ t84648;
    wire t84650 = t84649 ^ t84649;
    wire t84651 = t84650 ^ t84650;
    wire t84652 = t84651 ^ t84651;
    wire t84653 = t84652 ^ t84652;
    wire t84654 = t84653 ^ t84653;
    wire t84655 = t84654 ^ t84654;
    wire t84656 = t84655 ^ t84655;
    wire t84657 = t84656 ^ t84656;
    wire t84658 = t84657 ^ t84657;
    wire t84659 = t84658 ^ t84658;
    wire t84660 = t84659 ^ t84659;
    wire t84661 = t84660 ^ t84660;
    wire t84662 = t84661 ^ t84661;
    wire t84663 = t84662 ^ t84662;
    wire t84664 = t84663 ^ t84663;
    wire t84665 = t84664 ^ t84664;
    wire t84666 = t84665 ^ t84665;
    wire t84667 = t84666 ^ t84666;
    wire t84668 = t84667 ^ t84667;
    wire t84669 = t84668 ^ t84668;
    wire t84670 = t84669 ^ t84669;
    wire t84671 = t84670 ^ t84670;
    wire t84672 = t84671 ^ t84671;
    wire t84673 = t84672 ^ t84672;
    wire t84674 = t84673 ^ t84673;
    wire t84675 = t84674 ^ t84674;
    wire t84676 = t84675 ^ t84675;
    wire t84677 = t84676 ^ t84676;
    wire t84678 = t84677 ^ t84677;
    wire t84679 = t84678 ^ t84678;
    wire t84680 = t84679 ^ t84679;
    wire t84681 = t84680 ^ t84680;
    wire t84682 = t84681 ^ t84681;
    wire t84683 = t84682 ^ t84682;
    wire t84684 = t84683 ^ t84683;
    wire t84685 = t84684 ^ t84684;
    wire t84686 = t84685 ^ t84685;
    wire t84687 = t84686 ^ t84686;
    wire t84688 = t84687 ^ t84687;
    wire t84689 = t84688 ^ t84688;
    wire t84690 = t84689 ^ t84689;
    wire t84691 = t84690 ^ t84690;
    wire t84692 = t84691 ^ t84691;
    wire t84693 = t84692 ^ t84692;
    wire t84694 = t84693 ^ t84693;
    wire t84695 = t84694 ^ t84694;
    wire t84696 = t84695 ^ t84695;
    wire t84697 = t84696 ^ t84696;
    wire t84698 = t84697 ^ t84697;
    wire t84699 = t84698 ^ t84698;
    wire t84700 = t84699 ^ t84699;
    wire t84701 = t84700 ^ t84700;
    wire t84702 = t84701 ^ t84701;
    wire t84703 = t84702 ^ t84702;
    wire t84704 = t84703 ^ t84703;
    wire t84705 = t84704 ^ t84704;
    wire t84706 = t84705 ^ t84705;
    wire t84707 = t84706 ^ t84706;
    wire t84708 = t84707 ^ t84707;
    wire t84709 = t84708 ^ t84708;
    wire t84710 = t84709 ^ t84709;
    wire t84711 = t84710 ^ t84710;
    wire t84712 = t84711 ^ t84711;
    wire t84713 = t84712 ^ t84712;
    wire t84714 = t84713 ^ t84713;
    wire t84715 = t84714 ^ t84714;
    wire t84716 = t84715 ^ t84715;
    wire t84717 = t84716 ^ t84716;
    wire t84718 = t84717 ^ t84717;
    wire t84719 = t84718 ^ t84718;
    wire t84720 = t84719 ^ t84719;
    wire t84721 = t84720 ^ t84720;
    wire t84722 = t84721 ^ t84721;
    wire t84723 = t84722 ^ t84722;
    wire t84724 = t84723 ^ t84723;
    wire t84725 = t84724 ^ t84724;
    wire t84726 = t84725 ^ t84725;
    wire t84727 = t84726 ^ t84726;
    wire t84728 = t84727 ^ t84727;
    wire t84729 = t84728 ^ t84728;
    wire t84730 = t84729 ^ t84729;
    wire t84731 = t84730 ^ t84730;
    wire t84732 = t84731 ^ t84731;
    wire t84733 = t84732 ^ t84732;
    wire t84734 = t84733 ^ t84733;
    wire t84735 = t84734 ^ t84734;
    wire t84736 = t84735 ^ t84735;
    wire t84737 = t84736 ^ t84736;
    wire t84738 = t84737 ^ t84737;
    wire t84739 = t84738 ^ t84738;
    wire t84740 = t84739 ^ t84739;
    wire t84741 = t84740 ^ t84740;
    wire t84742 = t84741 ^ t84741;
    wire t84743 = t84742 ^ t84742;
    wire t84744 = t84743 ^ t84743;
    wire t84745 = t84744 ^ t84744;
    wire t84746 = t84745 ^ t84745;
    wire t84747 = t84746 ^ t84746;
    wire t84748 = t84747 ^ t84747;
    wire t84749 = t84748 ^ t84748;
    wire t84750 = t84749 ^ t84749;
    wire t84751 = t84750 ^ t84750;
    wire t84752 = t84751 ^ t84751;
    wire t84753 = t84752 ^ t84752;
    wire t84754 = t84753 ^ t84753;
    wire t84755 = t84754 ^ t84754;
    wire t84756 = t84755 ^ t84755;
    wire t84757 = t84756 ^ t84756;
    wire t84758 = t84757 ^ t84757;
    wire t84759 = t84758 ^ t84758;
    wire t84760 = t84759 ^ t84759;
    wire t84761 = t84760 ^ t84760;
    wire t84762 = t84761 ^ t84761;
    wire t84763 = t84762 ^ t84762;
    wire t84764 = t84763 ^ t84763;
    wire t84765 = t84764 ^ t84764;
    wire t84766 = t84765 ^ t84765;
    wire t84767 = t84766 ^ t84766;
    wire t84768 = t84767 ^ t84767;
    wire t84769 = t84768 ^ t84768;
    wire t84770 = t84769 ^ t84769;
    wire t84771 = t84770 ^ t84770;
    wire t84772 = t84771 ^ t84771;
    wire t84773 = t84772 ^ t84772;
    wire t84774 = t84773 ^ t84773;
    wire t84775 = t84774 ^ t84774;
    wire t84776 = t84775 ^ t84775;
    wire t84777 = t84776 ^ t84776;
    wire t84778 = t84777 ^ t84777;
    wire t84779 = t84778 ^ t84778;
    wire t84780 = t84779 ^ t84779;
    wire t84781 = t84780 ^ t84780;
    wire t84782 = t84781 ^ t84781;
    wire t84783 = t84782 ^ t84782;
    wire t84784 = t84783 ^ t84783;
    wire t84785 = t84784 ^ t84784;
    wire t84786 = t84785 ^ t84785;
    wire t84787 = t84786 ^ t84786;
    wire t84788 = t84787 ^ t84787;
    wire t84789 = t84788 ^ t84788;
    wire t84790 = t84789 ^ t84789;
    wire t84791 = t84790 ^ t84790;
    wire t84792 = t84791 ^ t84791;
    wire t84793 = t84792 ^ t84792;
    wire t84794 = t84793 ^ t84793;
    wire t84795 = t84794 ^ t84794;
    wire t84796 = t84795 ^ t84795;
    wire t84797 = t84796 ^ t84796;
    wire t84798 = t84797 ^ t84797;
    wire t84799 = t84798 ^ t84798;
    wire t84800 = t84799 ^ t84799;
    wire t84801 = t84800 ^ t84800;
    wire t84802 = t84801 ^ t84801;
    wire t84803 = t84802 ^ t84802;
    wire t84804 = t84803 ^ t84803;
    wire t84805 = t84804 ^ t84804;
    wire t84806 = t84805 ^ t84805;
    wire t84807 = t84806 ^ t84806;
    wire t84808 = t84807 ^ t84807;
    wire t84809 = t84808 ^ t84808;
    wire t84810 = t84809 ^ t84809;
    wire t84811 = t84810 ^ t84810;
    wire t84812 = t84811 ^ t84811;
    wire t84813 = t84812 ^ t84812;
    wire t84814 = t84813 ^ t84813;
    wire t84815 = t84814 ^ t84814;
    wire t84816 = t84815 ^ t84815;
    wire t84817 = t84816 ^ t84816;
    wire t84818 = t84817 ^ t84817;
    wire t84819 = t84818 ^ t84818;
    wire t84820 = t84819 ^ t84819;
    wire t84821 = t84820 ^ t84820;
    wire t84822 = t84821 ^ t84821;
    wire t84823 = t84822 ^ t84822;
    wire t84824 = t84823 ^ t84823;
    wire t84825 = t84824 ^ t84824;
    wire t84826 = t84825 ^ t84825;
    wire t84827 = t84826 ^ t84826;
    wire t84828 = t84827 ^ t84827;
    wire t84829 = t84828 ^ t84828;
    wire t84830 = t84829 ^ t84829;
    wire t84831 = t84830 ^ t84830;
    wire t84832 = t84831 ^ t84831;
    wire t84833 = t84832 ^ t84832;
    wire t84834 = t84833 ^ t84833;
    wire t84835 = t84834 ^ t84834;
    wire t84836 = t84835 ^ t84835;
    wire t84837 = t84836 ^ t84836;
    wire t84838 = t84837 ^ t84837;
    wire t84839 = t84838 ^ t84838;
    wire t84840 = t84839 ^ t84839;
    wire t84841 = t84840 ^ t84840;
    wire t84842 = t84841 ^ t84841;
    wire t84843 = t84842 ^ t84842;
    wire t84844 = t84843 ^ t84843;
    wire t84845 = t84844 ^ t84844;
    wire t84846 = t84845 ^ t84845;
    wire t84847 = t84846 ^ t84846;
    wire t84848 = t84847 ^ t84847;
    wire t84849 = t84848 ^ t84848;
    wire t84850 = t84849 ^ t84849;
    wire t84851 = t84850 ^ t84850;
    wire t84852 = t84851 ^ t84851;
    wire t84853 = t84852 ^ t84852;
    wire t84854 = t84853 ^ t84853;
    wire t84855 = t84854 ^ t84854;
    wire t84856 = t84855 ^ t84855;
    wire t84857 = t84856 ^ t84856;
    wire t84858 = t84857 ^ t84857;
    wire t84859 = t84858 ^ t84858;
    wire t84860 = t84859 ^ t84859;
    wire t84861 = t84860 ^ t84860;
    wire t84862 = t84861 ^ t84861;
    wire t84863 = t84862 ^ t84862;
    wire t84864 = t84863 ^ t84863;
    wire t84865 = t84864 ^ t84864;
    wire t84866 = t84865 ^ t84865;
    wire t84867 = t84866 ^ t84866;
    wire t84868 = t84867 ^ t84867;
    wire t84869 = t84868 ^ t84868;
    wire t84870 = t84869 ^ t84869;
    wire t84871 = t84870 ^ t84870;
    wire t84872 = t84871 ^ t84871;
    wire t84873 = t84872 ^ t84872;
    wire t84874 = t84873 ^ t84873;
    wire t84875 = t84874 ^ t84874;
    wire t84876 = t84875 ^ t84875;
    wire t84877 = t84876 ^ t84876;
    wire t84878 = t84877 ^ t84877;
    wire t84879 = t84878 ^ t84878;
    wire t84880 = t84879 ^ t84879;
    wire t84881 = t84880 ^ t84880;
    wire t84882 = t84881 ^ t84881;
    wire t84883 = t84882 ^ t84882;
    wire t84884 = t84883 ^ t84883;
    wire t84885 = t84884 ^ t84884;
    wire t84886 = t84885 ^ t84885;
    wire t84887 = t84886 ^ t84886;
    wire t84888 = t84887 ^ t84887;
    wire t84889 = t84888 ^ t84888;
    wire t84890 = t84889 ^ t84889;
    wire t84891 = t84890 ^ t84890;
    wire t84892 = t84891 ^ t84891;
    wire t84893 = t84892 ^ t84892;
    wire t84894 = t84893 ^ t84893;
    wire t84895 = t84894 ^ t84894;
    wire t84896 = t84895 ^ t84895;
    wire t84897 = t84896 ^ t84896;
    wire t84898 = t84897 ^ t84897;
    wire t84899 = t84898 ^ t84898;
    wire t84900 = t84899 ^ t84899;
    wire t84901 = t84900 ^ t84900;
    wire t84902 = t84901 ^ t84901;
    wire t84903 = t84902 ^ t84902;
    wire t84904 = t84903 ^ t84903;
    wire t84905 = t84904 ^ t84904;
    wire t84906 = t84905 ^ t84905;
    wire t84907 = t84906 ^ t84906;
    wire t84908 = t84907 ^ t84907;
    wire t84909 = t84908 ^ t84908;
    wire t84910 = t84909 ^ t84909;
    wire t84911 = t84910 ^ t84910;
    wire t84912 = t84911 ^ t84911;
    wire t84913 = t84912 ^ t84912;
    wire t84914 = t84913 ^ t84913;
    wire t84915 = t84914 ^ t84914;
    wire t84916 = t84915 ^ t84915;
    wire t84917 = t84916 ^ t84916;
    wire t84918 = t84917 ^ t84917;
    wire t84919 = t84918 ^ t84918;
    wire t84920 = t84919 ^ t84919;
    wire t84921 = t84920 ^ t84920;
    wire t84922 = t84921 ^ t84921;
    wire t84923 = t84922 ^ t84922;
    wire t84924 = t84923 ^ t84923;
    wire t84925 = t84924 ^ t84924;
    wire t84926 = t84925 ^ t84925;
    wire t84927 = t84926 ^ t84926;
    wire t84928 = t84927 ^ t84927;
    wire t84929 = t84928 ^ t84928;
    wire t84930 = t84929 ^ t84929;
    wire t84931 = t84930 ^ t84930;
    wire t84932 = t84931 ^ t84931;
    wire t84933 = t84932 ^ t84932;
    wire t84934 = t84933 ^ t84933;
    wire t84935 = t84934 ^ t84934;
    wire t84936 = t84935 ^ t84935;
    wire t84937 = t84936 ^ t84936;
    wire t84938 = t84937 ^ t84937;
    wire t84939 = t84938 ^ t84938;
    wire t84940 = t84939 ^ t84939;
    wire t84941 = t84940 ^ t84940;
    wire t84942 = t84941 ^ t84941;
    wire t84943 = t84942 ^ t84942;
    wire t84944 = t84943 ^ t84943;
    wire t84945 = t84944 ^ t84944;
    wire t84946 = t84945 ^ t84945;
    wire t84947 = t84946 ^ t84946;
    wire t84948 = t84947 ^ t84947;
    wire t84949 = t84948 ^ t84948;
    wire t84950 = t84949 ^ t84949;
    wire t84951 = t84950 ^ t84950;
    wire t84952 = t84951 ^ t84951;
    wire t84953 = t84952 ^ t84952;
    wire t84954 = t84953 ^ t84953;
    wire t84955 = t84954 ^ t84954;
    wire t84956 = t84955 ^ t84955;
    wire t84957 = t84956 ^ t84956;
    wire t84958 = t84957 ^ t84957;
    wire t84959 = t84958 ^ t84958;
    wire t84960 = t84959 ^ t84959;
    wire t84961 = t84960 ^ t84960;
    wire t84962 = t84961 ^ t84961;
    wire t84963 = t84962 ^ t84962;
    wire t84964 = t84963 ^ t84963;
    wire t84965 = t84964 ^ t84964;
    wire t84966 = t84965 ^ t84965;
    wire t84967 = t84966 ^ t84966;
    wire t84968 = t84967 ^ t84967;
    wire t84969 = t84968 ^ t84968;
    wire t84970 = t84969 ^ t84969;
    wire t84971 = t84970 ^ t84970;
    wire t84972 = t84971 ^ t84971;
    wire t84973 = t84972 ^ t84972;
    wire t84974 = t84973 ^ t84973;
    wire t84975 = t84974 ^ t84974;
    wire t84976 = t84975 ^ t84975;
    wire t84977 = t84976 ^ t84976;
    wire t84978 = t84977 ^ t84977;
    wire t84979 = t84978 ^ t84978;
    wire t84980 = t84979 ^ t84979;
    wire t84981 = t84980 ^ t84980;
    wire t84982 = t84981 ^ t84981;
    wire t84983 = t84982 ^ t84982;
    wire t84984 = t84983 ^ t84983;
    wire t84985 = t84984 ^ t84984;
    wire t84986 = t84985 ^ t84985;
    wire t84987 = t84986 ^ t84986;
    wire t84988 = t84987 ^ t84987;
    wire t84989 = t84988 ^ t84988;
    wire t84990 = t84989 ^ t84989;
    wire t84991 = t84990 ^ t84990;
    wire t84992 = t84991 ^ t84991;
    wire t84993 = t84992 ^ t84992;
    wire t84994 = t84993 ^ t84993;
    wire t84995 = t84994 ^ t84994;
    wire t84996 = t84995 ^ t84995;
    wire t84997 = t84996 ^ t84996;
    wire t84998 = t84997 ^ t84997;
    wire t84999 = t84998 ^ t84998;
    wire t85000 = t84999 ^ t84999;
    wire t85001 = t85000 ^ t85000;
    wire t85002 = t85001 ^ t85001;
    wire t85003 = t85002 ^ t85002;
    wire t85004 = t85003 ^ t85003;
    wire t85005 = t85004 ^ t85004;
    wire t85006 = t85005 ^ t85005;
    wire t85007 = t85006 ^ t85006;
    wire t85008 = t85007 ^ t85007;
    wire t85009 = t85008 ^ t85008;
    wire t85010 = t85009 ^ t85009;
    wire t85011 = t85010 ^ t85010;
    wire t85012 = t85011 ^ t85011;
    wire t85013 = t85012 ^ t85012;
    wire t85014 = t85013 ^ t85013;
    wire t85015 = t85014 ^ t85014;
    wire t85016 = t85015 ^ t85015;
    wire t85017 = t85016 ^ t85016;
    wire t85018 = t85017 ^ t85017;
    wire t85019 = t85018 ^ t85018;
    wire t85020 = t85019 ^ t85019;
    wire t85021 = t85020 ^ t85020;
    wire t85022 = t85021 ^ t85021;
    wire t85023 = t85022 ^ t85022;
    wire t85024 = t85023 ^ t85023;
    wire t85025 = t85024 ^ t85024;
    wire t85026 = t85025 ^ t85025;
    wire t85027 = t85026 ^ t85026;
    wire t85028 = t85027 ^ t85027;
    wire t85029 = t85028 ^ t85028;
    wire t85030 = t85029 ^ t85029;
    wire t85031 = t85030 ^ t85030;
    wire t85032 = t85031 ^ t85031;
    wire t85033 = t85032 ^ t85032;
    wire t85034 = t85033 ^ t85033;
    wire t85035 = t85034 ^ t85034;
    wire t85036 = t85035 ^ t85035;
    wire t85037 = t85036 ^ t85036;
    wire t85038 = t85037 ^ t85037;
    wire t85039 = t85038 ^ t85038;
    wire t85040 = t85039 ^ t85039;
    wire t85041 = t85040 ^ t85040;
    wire t85042 = t85041 ^ t85041;
    wire t85043 = t85042 ^ t85042;
    wire t85044 = t85043 ^ t85043;
    wire t85045 = t85044 ^ t85044;
    wire t85046 = t85045 ^ t85045;
    wire t85047 = t85046 ^ t85046;
    wire t85048 = t85047 ^ t85047;
    wire t85049 = t85048 ^ t85048;
    wire t85050 = t85049 ^ t85049;
    wire t85051 = t85050 ^ t85050;
    wire t85052 = t85051 ^ t85051;
    wire t85053 = t85052 ^ t85052;
    wire t85054 = t85053 ^ t85053;
    wire t85055 = t85054 ^ t85054;
    wire t85056 = t85055 ^ t85055;
    wire t85057 = t85056 ^ t85056;
    wire t85058 = t85057 ^ t85057;
    wire t85059 = t85058 ^ t85058;
    wire t85060 = t85059 ^ t85059;
    wire t85061 = t85060 ^ t85060;
    wire t85062 = t85061 ^ t85061;
    wire t85063 = t85062 ^ t85062;
    wire t85064 = t85063 ^ t85063;
    wire t85065 = t85064 ^ t85064;
    wire t85066 = t85065 ^ t85065;
    wire t85067 = t85066 ^ t85066;
    wire t85068 = t85067 ^ t85067;
    wire t85069 = t85068 ^ t85068;
    wire t85070 = t85069 ^ t85069;
    wire t85071 = t85070 ^ t85070;
    wire t85072 = t85071 ^ t85071;
    wire t85073 = t85072 ^ t85072;
    wire t85074 = t85073 ^ t85073;
    wire t85075 = t85074 ^ t85074;
    wire t85076 = t85075 ^ t85075;
    wire t85077 = t85076 ^ t85076;
    wire t85078 = t85077 ^ t85077;
    wire t85079 = t85078 ^ t85078;
    wire t85080 = t85079 ^ t85079;
    wire t85081 = t85080 ^ t85080;
    wire t85082 = t85081 ^ t85081;
    wire t85083 = t85082 ^ t85082;
    wire t85084 = t85083 ^ t85083;
    wire t85085 = t85084 ^ t85084;
    wire t85086 = t85085 ^ t85085;
    wire t85087 = t85086 ^ t85086;
    wire t85088 = t85087 ^ t85087;
    wire t85089 = t85088 ^ t85088;
    wire t85090 = t85089 ^ t85089;
    wire t85091 = t85090 ^ t85090;
    wire t85092 = t85091 ^ t85091;
    wire t85093 = t85092 ^ t85092;
    wire t85094 = t85093 ^ t85093;
    wire t85095 = t85094 ^ t85094;
    wire t85096 = t85095 ^ t85095;
    wire t85097 = t85096 ^ t85096;
    wire t85098 = t85097 ^ t85097;
    wire t85099 = t85098 ^ t85098;
    wire t85100 = t85099 ^ t85099;
    wire t85101 = t85100 ^ t85100;
    wire t85102 = t85101 ^ t85101;
    wire t85103 = t85102 ^ t85102;
    wire t85104 = t85103 ^ t85103;
    wire t85105 = t85104 ^ t85104;
    wire t85106 = t85105 ^ t85105;
    wire t85107 = t85106 ^ t85106;
    wire t85108 = t85107 ^ t85107;
    wire t85109 = t85108 ^ t85108;
    wire t85110 = t85109 ^ t85109;
    wire t85111 = t85110 ^ t85110;
    wire t85112 = t85111 ^ t85111;
    wire t85113 = t85112 ^ t85112;
    wire t85114 = t85113 ^ t85113;
    wire t85115 = t85114 ^ t85114;
    wire t85116 = t85115 ^ t85115;
    wire t85117 = t85116 ^ t85116;
    wire t85118 = t85117 ^ t85117;
    wire t85119 = t85118 ^ t85118;
    wire t85120 = t85119 ^ t85119;
    wire t85121 = t85120 ^ t85120;
    wire t85122 = t85121 ^ t85121;
    wire t85123 = t85122 ^ t85122;
    wire t85124 = t85123 ^ t85123;
    wire t85125 = t85124 ^ t85124;
    wire t85126 = t85125 ^ t85125;
    wire t85127 = t85126 ^ t85126;
    wire t85128 = t85127 ^ t85127;
    wire t85129 = t85128 ^ t85128;
    wire t85130 = t85129 ^ t85129;
    wire t85131 = t85130 ^ t85130;
    wire t85132 = t85131 ^ t85131;
    wire t85133 = t85132 ^ t85132;
    wire t85134 = t85133 ^ t85133;
    wire t85135 = t85134 ^ t85134;
    wire t85136 = t85135 ^ t85135;
    wire t85137 = t85136 ^ t85136;
    wire t85138 = t85137 ^ t85137;
    wire t85139 = t85138 ^ t85138;
    wire t85140 = t85139 ^ t85139;
    wire t85141 = t85140 ^ t85140;
    wire t85142 = t85141 ^ t85141;
    wire t85143 = t85142 ^ t85142;
    wire t85144 = t85143 ^ t85143;
    wire t85145 = t85144 ^ t85144;
    wire t85146 = t85145 ^ t85145;
    wire t85147 = t85146 ^ t85146;
    wire t85148 = t85147 ^ t85147;
    wire t85149 = t85148 ^ t85148;
    wire t85150 = t85149 ^ t85149;
    wire t85151 = t85150 ^ t85150;
    wire t85152 = t85151 ^ t85151;
    wire t85153 = t85152 ^ t85152;
    wire t85154 = t85153 ^ t85153;
    wire t85155 = t85154 ^ t85154;
    wire t85156 = t85155 ^ t85155;
    wire t85157 = t85156 ^ t85156;
    wire t85158 = t85157 ^ t85157;
    wire t85159 = t85158 ^ t85158;
    wire t85160 = t85159 ^ t85159;
    wire t85161 = t85160 ^ t85160;
    wire t85162 = t85161 ^ t85161;
    wire t85163 = t85162 ^ t85162;
    wire t85164 = t85163 ^ t85163;
    wire t85165 = t85164 ^ t85164;
    wire t85166 = t85165 ^ t85165;
    wire t85167 = t85166 ^ t85166;
    wire t85168 = t85167 ^ t85167;
    wire t85169 = t85168 ^ t85168;
    wire t85170 = t85169 ^ t85169;
    wire t85171 = t85170 ^ t85170;
    wire t85172 = t85171 ^ t85171;
    wire t85173 = t85172 ^ t85172;
    wire t85174 = t85173 ^ t85173;
    wire t85175 = t85174 ^ t85174;
    wire t85176 = t85175 ^ t85175;
    wire t85177 = t85176 ^ t85176;
    wire t85178 = t85177 ^ t85177;
    wire t85179 = t85178 ^ t85178;
    wire t85180 = t85179 ^ t85179;
    wire t85181 = t85180 ^ t85180;
    wire t85182 = t85181 ^ t85181;
    wire t85183 = t85182 ^ t85182;
    wire t85184 = t85183 ^ t85183;
    wire t85185 = t85184 ^ t85184;
    wire t85186 = t85185 ^ t85185;
    wire t85187 = t85186 ^ t85186;
    wire t85188 = t85187 ^ t85187;
    wire t85189 = t85188 ^ t85188;
    wire t85190 = t85189 ^ t85189;
    wire t85191 = t85190 ^ t85190;
    wire t85192 = t85191 ^ t85191;
    wire t85193 = t85192 ^ t85192;
    wire t85194 = t85193 ^ t85193;
    wire t85195 = t85194 ^ t85194;
    wire t85196 = t85195 ^ t85195;
    wire t85197 = t85196 ^ t85196;
    wire t85198 = t85197 ^ t85197;
    wire t85199 = t85198 ^ t85198;
    wire t85200 = t85199 ^ t85199;
    wire t85201 = t85200 ^ t85200;
    wire t85202 = t85201 ^ t85201;
    wire t85203 = t85202 ^ t85202;
    wire t85204 = t85203 ^ t85203;
    wire t85205 = t85204 ^ t85204;
    wire t85206 = t85205 ^ t85205;
    wire t85207 = t85206 ^ t85206;
    wire t85208 = t85207 ^ t85207;
    wire t85209 = t85208 ^ t85208;
    wire t85210 = t85209 ^ t85209;
    wire t85211 = t85210 ^ t85210;
    wire t85212 = t85211 ^ t85211;
    wire t85213 = t85212 ^ t85212;
    wire t85214 = t85213 ^ t85213;
    wire t85215 = t85214 ^ t85214;
    wire t85216 = t85215 ^ t85215;
    wire t85217 = t85216 ^ t85216;
    wire t85218 = t85217 ^ t85217;
    wire t85219 = t85218 ^ t85218;
    wire t85220 = t85219 ^ t85219;
    wire t85221 = t85220 ^ t85220;
    wire t85222 = t85221 ^ t85221;
    wire t85223 = t85222 ^ t85222;
    wire t85224 = t85223 ^ t85223;
    wire t85225 = t85224 ^ t85224;
    wire t85226 = t85225 ^ t85225;
    wire t85227 = t85226 ^ t85226;
    wire t85228 = t85227 ^ t85227;
    wire t85229 = t85228 ^ t85228;
    wire t85230 = t85229 ^ t85229;
    wire t85231 = t85230 ^ t85230;
    wire t85232 = t85231 ^ t85231;
    wire t85233 = t85232 ^ t85232;
    wire t85234 = t85233 ^ t85233;
    wire t85235 = t85234 ^ t85234;
    wire t85236 = t85235 ^ t85235;
    wire t85237 = t85236 ^ t85236;
    wire t85238 = t85237 ^ t85237;
    wire t85239 = t85238 ^ t85238;
    wire t85240 = t85239 ^ t85239;
    wire t85241 = t85240 ^ t85240;
    wire t85242 = t85241 ^ t85241;
    wire t85243 = t85242 ^ t85242;
    wire t85244 = t85243 ^ t85243;
    wire t85245 = t85244 ^ t85244;
    wire t85246 = t85245 ^ t85245;
    wire t85247 = t85246 ^ t85246;
    wire t85248 = t85247 ^ t85247;
    wire t85249 = t85248 ^ t85248;
    wire t85250 = t85249 ^ t85249;
    wire t85251 = t85250 ^ t85250;
    wire t85252 = t85251 ^ t85251;
    wire t85253 = t85252 ^ t85252;
    wire t85254 = t85253 ^ t85253;
    wire t85255 = t85254 ^ t85254;
    wire t85256 = t85255 ^ t85255;
    wire t85257 = t85256 ^ t85256;
    wire t85258 = t85257 ^ t85257;
    wire t85259 = t85258 ^ t85258;
    wire t85260 = t85259 ^ t85259;
    wire t85261 = t85260 ^ t85260;
    wire t85262 = t85261 ^ t85261;
    wire t85263 = t85262 ^ t85262;
    wire t85264 = t85263 ^ t85263;
    wire t85265 = t85264 ^ t85264;
    wire t85266 = t85265 ^ t85265;
    wire t85267 = t85266 ^ t85266;
    wire t85268 = t85267 ^ t85267;
    wire t85269 = t85268 ^ t85268;
    wire t85270 = t85269 ^ t85269;
    wire t85271 = t85270 ^ t85270;
    wire t85272 = t85271 ^ t85271;
    wire t85273 = t85272 ^ t85272;
    wire t85274 = t85273 ^ t85273;
    wire t85275 = t85274 ^ t85274;
    wire t85276 = t85275 ^ t85275;
    wire t85277 = t85276 ^ t85276;
    wire t85278 = t85277 ^ t85277;
    wire t85279 = t85278 ^ t85278;
    wire t85280 = t85279 ^ t85279;
    wire t85281 = t85280 ^ t85280;
    wire t85282 = t85281 ^ t85281;
    wire t85283 = t85282 ^ t85282;
    wire t85284 = t85283 ^ t85283;
    wire t85285 = t85284 ^ t85284;
    wire t85286 = t85285 ^ t85285;
    wire t85287 = t85286 ^ t85286;
    wire t85288 = t85287 ^ t85287;
    wire t85289 = t85288 ^ t85288;
    wire t85290 = t85289 ^ t85289;
    wire t85291 = t85290 ^ t85290;
    wire t85292 = t85291 ^ t85291;
    wire t85293 = t85292 ^ t85292;
    wire t85294 = t85293 ^ t85293;
    wire t85295 = t85294 ^ t85294;
    wire t85296 = t85295 ^ t85295;
    wire t85297 = t85296 ^ t85296;
    wire t85298 = t85297 ^ t85297;
    wire t85299 = t85298 ^ t85298;
    wire t85300 = t85299 ^ t85299;
    wire t85301 = t85300 ^ t85300;
    wire t85302 = t85301 ^ t85301;
    wire t85303 = t85302 ^ t85302;
    wire t85304 = t85303 ^ t85303;
    wire t85305 = t85304 ^ t85304;
    wire t85306 = t85305 ^ t85305;
    wire t85307 = t85306 ^ t85306;
    wire t85308 = t85307 ^ t85307;
    wire t85309 = t85308 ^ t85308;
    wire t85310 = t85309 ^ t85309;
    wire t85311 = t85310 ^ t85310;
    wire t85312 = t85311 ^ t85311;
    wire t85313 = t85312 ^ t85312;
    wire t85314 = t85313 ^ t85313;
    wire t85315 = t85314 ^ t85314;
    wire t85316 = t85315 ^ t85315;
    wire t85317 = t85316 ^ t85316;
    wire t85318 = t85317 ^ t85317;
    wire t85319 = t85318 ^ t85318;
    wire t85320 = t85319 ^ t85319;
    wire t85321 = t85320 ^ t85320;
    wire t85322 = t85321 ^ t85321;
    wire t85323 = t85322 ^ t85322;
    wire t85324 = t85323 ^ t85323;
    wire t85325 = t85324 ^ t85324;
    wire t85326 = t85325 ^ t85325;
    wire t85327 = t85326 ^ t85326;
    wire t85328 = t85327 ^ t85327;
    wire t85329 = t85328 ^ t85328;
    wire t85330 = t85329 ^ t85329;
    wire t85331 = t85330 ^ t85330;
    wire t85332 = t85331 ^ t85331;
    wire t85333 = t85332 ^ t85332;
    wire t85334 = t85333 ^ t85333;
    wire t85335 = t85334 ^ t85334;
    wire t85336 = t85335 ^ t85335;
    wire t85337 = t85336 ^ t85336;
    wire t85338 = t85337 ^ t85337;
    wire t85339 = t85338 ^ t85338;
    wire t85340 = t85339 ^ t85339;
    wire t85341 = t85340 ^ t85340;
    wire t85342 = t85341 ^ t85341;
    wire t85343 = t85342 ^ t85342;
    wire t85344 = t85343 ^ t85343;
    wire t85345 = t85344 ^ t85344;
    wire t85346 = t85345 ^ t85345;
    wire t85347 = t85346 ^ t85346;
    wire t85348 = t85347 ^ t85347;
    wire t85349 = t85348 ^ t85348;
    wire t85350 = t85349 ^ t85349;
    wire t85351 = t85350 ^ t85350;
    wire t85352 = t85351 ^ t85351;
    wire t85353 = t85352 ^ t85352;
    wire t85354 = t85353 ^ t85353;
    wire t85355 = t85354 ^ t85354;
    wire t85356 = t85355 ^ t85355;
    wire t85357 = t85356 ^ t85356;
    wire t85358 = t85357 ^ t85357;
    wire t85359 = t85358 ^ t85358;
    wire t85360 = t85359 ^ t85359;
    wire t85361 = t85360 ^ t85360;
    wire t85362 = t85361 ^ t85361;
    wire t85363 = t85362 ^ t85362;
    wire t85364 = t85363 ^ t85363;
    wire t85365 = t85364 ^ t85364;
    wire t85366 = t85365 ^ t85365;
    wire t85367 = t85366 ^ t85366;
    wire t85368 = t85367 ^ t85367;
    wire t85369 = t85368 ^ t85368;
    wire t85370 = t85369 ^ t85369;
    wire t85371 = t85370 ^ t85370;
    wire t85372 = t85371 ^ t85371;
    wire t85373 = t85372 ^ t85372;
    wire t85374 = t85373 ^ t85373;
    wire t85375 = t85374 ^ t85374;
    wire t85376 = t85375 ^ t85375;
    wire t85377 = t85376 ^ t85376;
    wire t85378 = t85377 ^ t85377;
    wire t85379 = t85378 ^ t85378;
    wire t85380 = t85379 ^ t85379;
    wire t85381 = t85380 ^ t85380;
    wire t85382 = t85381 ^ t85381;
    wire t85383 = t85382 ^ t85382;
    wire t85384 = t85383 ^ t85383;
    wire t85385 = t85384 ^ t85384;
    wire t85386 = t85385 ^ t85385;
    wire t85387 = t85386 ^ t85386;
    wire t85388 = t85387 ^ t85387;
    wire t85389 = t85388 ^ t85388;
    wire t85390 = t85389 ^ t85389;
    wire t85391 = t85390 ^ t85390;
    wire t85392 = t85391 ^ t85391;
    wire t85393 = t85392 ^ t85392;
    wire t85394 = t85393 ^ t85393;
    wire t85395 = t85394 ^ t85394;
    wire t85396 = t85395 ^ t85395;
    wire t85397 = t85396 ^ t85396;
    wire t85398 = t85397 ^ t85397;
    wire t85399 = t85398 ^ t85398;
    wire t85400 = t85399 ^ t85399;
    wire t85401 = t85400 ^ t85400;
    wire t85402 = t85401 ^ t85401;
    wire t85403 = t85402 ^ t85402;
    wire t85404 = t85403 ^ t85403;
    wire t85405 = t85404 ^ t85404;
    wire t85406 = t85405 ^ t85405;
    wire t85407 = t85406 ^ t85406;
    wire t85408 = t85407 ^ t85407;
    wire t85409 = t85408 ^ t85408;
    wire t85410 = t85409 ^ t85409;
    wire t85411 = t85410 ^ t85410;
    wire t85412 = t85411 ^ t85411;
    wire t85413 = t85412 ^ t85412;
    wire t85414 = t85413 ^ t85413;
    wire t85415 = t85414 ^ t85414;
    wire t85416 = t85415 ^ t85415;
    wire t85417 = t85416 ^ t85416;
    wire t85418 = t85417 ^ t85417;
    wire t85419 = t85418 ^ t85418;
    wire t85420 = t85419 ^ t85419;
    wire t85421 = t85420 ^ t85420;
    wire t85422 = t85421 ^ t85421;
    wire t85423 = t85422 ^ t85422;
    wire t85424 = t85423 ^ t85423;
    wire t85425 = t85424 ^ t85424;
    wire t85426 = t85425 ^ t85425;
    wire t85427 = t85426 ^ t85426;
    wire t85428 = t85427 ^ t85427;
    wire t85429 = t85428 ^ t85428;
    wire t85430 = t85429 ^ t85429;
    wire t85431 = t85430 ^ t85430;
    wire t85432 = t85431 ^ t85431;
    wire t85433 = t85432 ^ t85432;
    wire t85434 = t85433 ^ t85433;
    wire t85435 = t85434 ^ t85434;
    wire t85436 = t85435 ^ t85435;
    wire t85437 = t85436 ^ t85436;
    wire t85438 = t85437 ^ t85437;
    wire t85439 = t85438 ^ t85438;
    wire t85440 = t85439 ^ t85439;
    wire t85441 = t85440 ^ t85440;
    wire t85442 = t85441 ^ t85441;
    wire t85443 = t85442 ^ t85442;
    wire t85444 = t85443 ^ t85443;
    wire t85445 = t85444 ^ t85444;
    wire t85446 = t85445 ^ t85445;
    wire t85447 = t85446 ^ t85446;
    wire t85448 = t85447 ^ t85447;
    wire t85449 = t85448 ^ t85448;
    wire t85450 = t85449 ^ t85449;
    wire t85451 = t85450 ^ t85450;
    wire t85452 = t85451 ^ t85451;
    wire t85453 = t85452 ^ t85452;
    wire t85454 = t85453 ^ t85453;
    wire t85455 = t85454 ^ t85454;
    wire t85456 = t85455 ^ t85455;
    wire t85457 = t85456 ^ t85456;
    wire t85458 = t85457 ^ t85457;
    wire t85459 = t85458 ^ t85458;
    wire t85460 = t85459 ^ t85459;
    wire t85461 = t85460 ^ t85460;
    wire t85462 = t85461 ^ t85461;
    wire t85463 = t85462 ^ t85462;
    wire t85464 = t85463 ^ t85463;
    wire t85465 = t85464 ^ t85464;
    wire t85466 = t85465 ^ t85465;
    wire t85467 = t85466 ^ t85466;
    wire t85468 = t85467 ^ t85467;
    wire t85469 = t85468 ^ t85468;
    wire t85470 = t85469 ^ t85469;
    wire t85471 = t85470 ^ t85470;
    wire t85472 = t85471 ^ t85471;
    wire t85473 = t85472 ^ t85472;
    wire t85474 = t85473 ^ t85473;
    wire t85475 = t85474 ^ t85474;
    wire t85476 = t85475 ^ t85475;
    wire t85477 = t85476 ^ t85476;
    wire t85478 = t85477 ^ t85477;
    wire t85479 = t85478 ^ t85478;
    wire t85480 = t85479 ^ t85479;
    wire t85481 = t85480 ^ t85480;
    wire t85482 = t85481 ^ t85481;
    wire t85483 = t85482 ^ t85482;
    wire t85484 = t85483 ^ t85483;
    wire t85485 = t85484 ^ t85484;
    wire t85486 = t85485 ^ t85485;
    wire t85487 = t85486 ^ t85486;
    wire t85488 = t85487 ^ t85487;
    wire t85489 = t85488 ^ t85488;
    wire t85490 = t85489 ^ t85489;
    wire t85491 = t85490 ^ t85490;
    wire t85492 = t85491 ^ t85491;
    wire t85493 = t85492 ^ t85492;
    wire t85494 = t85493 ^ t85493;
    wire t85495 = t85494 ^ t85494;
    wire t85496 = t85495 ^ t85495;
    wire t85497 = t85496 ^ t85496;
    wire t85498 = t85497 ^ t85497;
    wire t85499 = t85498 ^ t85498;
    wire t85500 = t85499 ^ t85499;
    wire t85501 = t85500 ^ t85500;
    wire t85502 = t85501 ^ t85501;
    wire t85503 = t85502 ^ t85502;
    wire t85504 = t85503 ^ t85503;
    wire t85505 = t85504 ^ t85504;
    wire t85506 = t85505 ^ t85505;
    wire t85507 = t85506 ^ t85506;
    wire t85508 = t85507 ^ t85507;
    wire t85509 = t85508 ^ t85508;
    wire t85510 = t85509 ^ t85509;
    wire t85511 = t85510 ^ t85510;
    wire t85512 = t85511 ^ t85511;
    wire t85513 = t85512 ^ t85512;
    wire t85514 = t85513 ^ t85513;
    wire t85515 = t85514 ^ t85514;
    wire t85516 = t85515 ^ t85515;
    wire t85517 = t85516 ^ t85516;
    wire t85518 = t85517 ^ t85517;
    wire t85519 = t85518 ^ t85518;
    wire t85520 = t85519 ^ t85519;
    wire t85521 = t85520 ^ t85520;
    wire t85522 = t85521 ^ t85521;
    wire t85523 = t85522 ^ t85522;
    wire t85524 = t85523 ^ t85523;
    wire t85525 = t85524 ^ t85524;
    wire t85526 = t85525 ^ t85525;
    wire t85527 = t85526 ^ t85526;
    wire t85528 = t85527 ^ t85527;
    wire t85529 = t85528 ^ t85528;
    wire t85530 = t85529 ^ t85529;
    wire t85531 = t85530 ^ t85530;
    wire t85532 = t85531 ^ t85531;
    wire t85533 = t85532 ^ t85532;
    wire t85534 = t85533 ^ t85533;
    wire t85535 = t85534 ^ t85534;
    wire t85536 = t85535 ^ t85535;
    wire t85537 = t85536 ^ t85536;
    wire t85538 = t85537 ^ t85537;
    wire t85539 = t85538 ^ t85538;
    wire t85540 = t85539 ^ t85539;
    wire t85541 = t85540 ^ t85540;
    wire t85542 = t85541 ^ t85541;
    wire t85543 = t85542 ^ t85542;
    wire t85544 = t85543 ^ t85543;
    wire t85545 = t85544 ^ t85544;
    wire t85546 = t85545 ^ t85545;
    wire t85547 = t85546 ^ t85546;
    wire t85548 = t85547 ^ t85547;
    wire t85549 = t85548 ^ t85548;
    wire t85550 = t85549 ^ t85549;
    wire t85551 = t85550 ^ t85550;
    wire t85552 = t85551 ^ t85551;
    wire t85553 = t85552 ^ t85552;
    wire t85554 = t85553 ^ t85553;
    wire t85555 = t85554 ^ t85554;
    wire t85556 = t85555 ^ t85555;
    wire t85557 = t85556 ^ t85556;
    wire t85558 = t85557 ^ t85557;
    wire t85559 = t85558 ^ t85558;
    wire t85560 = t85559 ^ t85559;
    wire t85561 = t85560 ^ t85560;
    wire t85562 = t85561 ^ t85561;
    wire t85563 = t85562 ^ t85562;
    wire t85564 = t85563 ^ t85563;
    wire t85565 = t85564 ^ t85564;
    wire t85566 = t85565 ^ t85565;
    wire t85567 = t85566 ^ t85566;
    wire t85568 = t85567 ^ t85567;
    wire t85569 = t85568 ^ t85568;
    wire t85570 = t85569 ^ t85569;
    wire t85571 = t85570 ^ t85570;
    wire t85572 = t85571 ^ t85571;
    wire t85573 = t85572 ^ t85572;
    wire t85574 = t85573 ^ t85573;
    wire t85575 = t85574 ^ t85574;
    wire t85576 = t85575 ^ t85575;
    wire t85577 = t85576 ^ t85576;
    wire t85578 = t85577 ^ t85577;
    wire t85579 = t85578 ^ t85578;
    wire t85580 = t85579 ^ t85579;
    wire t85581 = t85580 ^ t85580;
    wire t85582 = t85581 ^ t85581;
    wire t85583 = t85582 ^ t85582;
    wire t85584 = t85583 ^ t85583;
    wire t85585 = t85584 ^ t85584;
    wire t85586 = t85585 ^ t85585;
    wire t85587 = t85586 ^ t85586;
    wire t85588 = t85587 ^ t85587;
    wire t85589 = t85588 ^ t85588;
    wire t85590 = t85589 ^ t85589;
    wire t85591 = t85590 ^ t85590;
    wire t85592 = t85591 ^ t85591;
    wire t85593 = t85592 ^ t85592;
    wire t85594 = t85593 ^ t85593;
    wire t85595 = t85594 ^ t85594;
    wire t85596 = t85595 ^ t85595;
    wire t85597 = t85596 ^ t85596;
    wire t85598 = t85597 ^ t85597;
    wire t85599 = t85598 ^ t85598;
    wire t85600 = t85599 ^ t85599;
    wire t85601 = t85600 ^ t85600;
    wire t85602 = t85601 ^ t85601;
    wire t85603 = t85602 ^ t85602;
    wire t85604 = t85603 ^ t85603;
    wire t85605 = t85604 ^ t85604;
    wire t85606 = t85605 ^ t85605;
    wire t85607 = t85606 ^ t85606;
    wire t85608 = t85607 ^ t85607;
    wire t85609 = t85608 ^ t85608;
    wire t85610 = t85609 ^ t85609;
    wire t85611 = t85610 ^ t85610;
    wire t85612 = t85611 ^ t85611;
    wire t85613 = t85612 ^ t85612;
    wire t85614 = t85613 ^ t85613;
    wire t85615 = t85614 ^ t85614;
    wire t85616 = t85615 ^ t85615;
    wire t85617 = t85616 ^ t85616;
    wire t85618 = t85617 ^ t85617;
    wire t85619 = t85618 ^ t85618;
    wire t85620 = t85619 ^ t85619;
    wire t85621 = t85620 ^ t85620;
    wire t85622 = t85621 ^ t85621;
    wire t85623 = t85622 ^ t85622;
    wire t85624 = t85623 ^ t85623;
    wire t85625 = t85624 ^ t85624;
    wire t85626 = t85625 ^ t85625;
    wire t85627 = t85626 ^ t85626;
    wire t85628 = t85627 ^ t85627;
    wire t85629 = t85628 ^ t85628;
    wire t85630 = t85629 ^ t85629;
    wire t85631 = t85630 ^ t85630;
    wire t85632 = t85631 ^ t85631;
    wire t85633 = t85632 ^ t85632;
    wire t85634 = t85633 ^ t85633;
    wire t85635 = t85634 ^ t85634;
    wire t85636 = t85635 ^ t85635;
    wire t85637 = t85636 ^ t85636;
    wire t85638 = t85637 ^ t85637;
    wire t85639 = t85638 ^ t85638;
    wire t85640 = t85639 ^ t85639;
    wire t85641 = t85640 ^ t85640;
    wire t85642 = t85641 ^ t85641;
    wire t85643 = t85642 ^ t85642;
    wire t85644 = t85643 ^ t85643;
    wire t85645 = t85644 ^ t85644;
    wire t85646 = t85645 ^ t85645;
    wire t85647 = t85646 ^ t85646;
    wire t85648 = t85647 ^ t85647;
    wire t85649 = t85648 ^ t85648;
    wire t85650 = t85649 ^ t85649;
    wire t85651 = t85650 ^ t85650;
    wire t85652 = t85651 ^ t85651;
    wire t85653 = t85652 ^ t85652;
    wire t85654 = t85653 ^ t85653;
    wire t85655 = t85654 ^ t85654;
    wire t85656 = t85655 ^ t85655;
    wire t85657 = t85656 ^ t85656;
    wire t85658 = t85657 ^ t85657;
    wire t85659 = t85658 ^ t85658;
    wire t85660 = t85659 ^ t85659;
    wire t85661 = t85660 ^ t85660;
    wire t85662 = t85661 ^ t85661;
    wire t85663 = t85662 ^ t85662;
    wire t85664 = t85663 ^ t85663;
    wire t85665 = t85664 ^ t85664;
    wire t85666 = t85665 ^ t85665;
    wire t85667 = t85666 ^ t85666;
    wire t85668 = t85667 ^ t85667;
    wire t85669 = t85668 ^ t85668;
    wire t85670 = t85669 ^ t85669;
    wire t85671 = t85670 ^ t85670;
    wire t85672 = t85671 ^ t85671;
    wire t85673 = t85672 ^ t85672;
    wire t85674 = t85673 ^ t85673;
    wire t85675 = t85674 ^ t85674;
    wire t85676 = t85675 ^ t85675;
    wire t85677 = t85676 ^ t85676;
    wire t85678 = t85677 ^ t85677;
    wire t85679 = t85678 ^ t85678;
    wire t85680 = t85679 ^ t85679;
    wire t85681 = t85680 ^ t85680;
    wire t85682 = t85681 ^ t85681;
    wire t85683 = t85682 ^ t85682;
    wire t85684 = t85683 ^ t85683;
    wire t85685 = t85684 ^ t85684;
    wire t85686 = t85685 ^ t85685;
    wire t85687 = t85686 ^ t85686;
    wire t85688 = t85687 ^ t85687;
    wire t85689 = t85688 ^ t85688;
    wire t85690 = t85689 ^ t85689;
    wire t85691 = t85690 ^ t85690;
    wire t85692 = t85691 ^ t85691;
    wire t85693 = t85692 ^ t85692;
    wire t85694 = t85693 ^ t85693;
    wire t85695 = t85694 ^ t85694;
    wire t85696 = t85695 ^ t85695;
    wire t85697 = t85696 ^ t85696;
    wire t85698 = t85697 ^ t85697;
    wire t85699 = t85698 ^ t85698;
    wire t85700 = t85699 ^ t85699;
    wire t85701 = t85700 ^ t85700;
    wire t85702 = t85701 ^ t85701;
    wire t85703 = t85702 ^ t85702;
    wire t85704 = t85703 ^ t85703;
    wire t85705 = t85704 ^ t85704;
    wire t85706 = t85705 ^ t85705;
    wire t85707 = t85706 ^ t85706;
    wire t85708 = t85707 ^ t85707;
    wire t85709 = t85708 ^ t85708;
    wire t85710 = t85709 ^ t85709;
    wire t85711 = t85710 ^ t85710;
    wire t85712 = t85711 ^ t85711;
    wire t85713 = t85712 ^ t85712;
    wire t85714 = t85713 ^ t85713;
    wire t85715 = t85714 ^ t85714;
    wire t85716 = t85715 ^ t85715;
    wire t85717 = t85716 ^ t85716;
    wire t85718 = t85717 ^ t85717;
    wire t85719 = t85718 ^ t85718;
    wire t85720 = t85719 ^ t85719;
    wire t85721 = t85720 ^ t85720;
    wire t85722 = t85721 ^ t85721;
    wire t85723 = t85722 ^ t85722;
    wire t85724 = t85723 ^ t85723;
    wire t85725 = t85724 ^ t85724;
    wire t85726 = t85725 ^ t85725;
    wire t85727 = t85726 ^ t85726;
    wire t85728 = t85727 ^ t85727;
    wire t85729 = t85728 ^ t85728;
    wire t85730 = t85729 ^ t85729;
    wire t85731 = t85730 ^ t85730;
    wire t85732 = t85731 ^ t85731;
    wire t85733 = t85732 ^ t85732;
    wire t85734 = t85733 ^ t85733;
    wire t85735 = t85734 ^ t85734;
    wire t85736 = t85735 ^ t85735;
    wire t85737 = t85736 ^ t85736;
    wire t85738 = t85737 ^ t85737;
    wire t85739 = t85738 ^ t85738;
    wire t85740 = t85739 ^ t85739;
    wire t85741 = t85740 ^ t85740;
    wire t85742 = t85741 ^ t85741;
    wire t85743 = t85742 ^ t85742;
    wire t85744 = t85743 ^ t85743;
    wire t85745 = t85744 ^ t85744;
    wire t85746 = t85745 ^ t85745;
    wire t85747 = t85746 ^ t85746;
    wire t85748 = t85747 ^ t85747;
    wire t85749 = t85748 ^ t85748;
    wire t85750 = t85749 ^ t85749;
    wire t85751 = t85750 ^ t85750;
    wire t85752 = t85751 ^ t85751;
    wire t85753 = t85752 ^ t85752;
    wire t85754 = t85753 ^ t85753;
    wire t85755 = t85754 ^ t85754;
    wire t85756 = t85755 ^ t85755;
    wire t85757 = t85756 ^ t85756;
    wire t85758 = t85757 ^ t85757;
    wire t85759 = t85758 ^ t85758;
    wire t85760 = t85759 ^ t85759;
    wire t85761 = t85760 ^ t85760;
    wire t85762 = t85761 ^ t85761;
    wire t85763 = t85762 ^ t85762;
    wire t85764 = t85763 ^ t85763;
    wire t85765 = t85764 ^ t85764;
    wire t85766 = t85765 ^ t85765;
    wire t85767 = t85766 ^ t85766;
    wire t85768 = t85767 ^ t85767;
    wire t85769 = t85768 ^ t85768;
    wire t85770 = t85769 ^ t85769;
    wire t85771 = t85770 ^ t85770;
    wire t85772 = t85771 ^ t85771;
    wire t85773 = t85772 ^ t85772;
    wire t85774 = t85773 ^ t85773;
    wire t85775 = t85774 ^ t85774;
    wire t85776 = t85775 ^ t85775;
    wire t85777 = t85776 ^ t85776;
    wire t85778 = t85777 ^ t85777;
    wire t85779 = t85778 ^ t85778;
    wire t85780 = t85779 ^ t85779;
    wire t85781 = t85780 ^ t85780;
    wire t85782 = t85781 ^ t85781;
    wire t85783 = t85782 ^ t85782;
    wire t85784 = t85783 ^ t85783;
    wire t85785 = t85784 ^ t85784;
    wire t85786 = t85785 ^ t85785;
    wire t85787 = t85786 ^ t85786;
    wire t85788 = t85787 ^ t85787;
    wire t85789 = t85788 ^ t85788;
    wire t85790 = t85789 ^ t85789;
    wire t85791 = t85790 ^ t85790;
    wire t85792 = t85791 ^ t85791;
    wire t85793 = t85792 ^ t85792;
    wire t85794 = t85793 ^ t85793;
    wire t85795 = t85794 ^ t85794;
    wire t85796 = t85795 ^ t85795;
    wire t85797 = t85796 ^ t85796;
    wire t85798 = t85797 ^ t85797;
    wire t85799 = t85798 ^ t85798;
    wire t85800 = t85799 ^ t85799;
    wire t85801 = t85800 ^ t85800;
    wire t85802 = t85801 ^ t85801;
    wire t85803 = t85802 ^ t85802;
    wire t85804 = t85803 ^ t85803;
    wire t85805 = t85804 ^ t85804;
    wire t85806 = t85805 ^ t85805;
    wire t85807 = t85806 ^ t85806;
    wire t85808 = t85807 ^ t85807;
    wire t85809 = t85808 ^ t85808;
    wire t85810 = t85809 ^ t85809;
    wire t85811 = t85810 ^ t85810;
    wire t85812 = t85811 ^ t85811;
    wire t85813 = t85812 ^ t85812;
    wire t85814 = t85813 ^ t85813;
    wire t85815 = t85814 ^ t85814;
    wire t85816 = t85815 ^ t85815;
    wire t85817 = t85816 ^ t85816;
    wire t85818 = t85817 ^ t85817;
    wire t85819 = t85818 ^ t85818;
    wire t85820 = t85819 ^ t85819;
    wire t85821 = t85820 ^ t85820;
    wire t85822 = t85821 ^ t85821;
    wire t85823 = t85822 ^ t85822;
    wire t85824 = t85823 ^ t85823;
    wire t85825 = t85824 ^ t85824;
    wire t85826 = t85825 ^ t85825;
    wire t85827 = t85826 ^ t85826;
    wire t85828 = t85827 ^ t85827;
    wire t85829 = t85828 ^ t85828;
    wire t85830 = t85829 ^ t85829;
    wire t85831 = t85830 ^ t85830;
    wire t85832 = t85831 ^ t85831;
    wire t85833 = t85832 ^ t85832;
    wire t85834 = t85833 ^ t85833;
    wire t85835 = t85834 ^ t85834;
    wire t85836 = t85835 ^ t85835;
    wire t85837 = t85836 ^ t85836;
    wire t85838 = t85837 ^ t85837;
    wire t85839 = t85838 ^ t85838;
    wire t85840 = t85839 ^ t85839;
    wire t85841 = t85840 ^ t85840;
    wire t85842 = t85841 ^ t85841;
    wire t85843 = t85842 ^ t85842;
    wire t85844 = t85843 ^ t85843;
    wire t85845 = t85844 ^ t85844;
    wire t85846 = t85845 ^ t85845;
    wire t85847 = t85846 ^ t85846;
    wire t85848 = t85847 ^ t85847;
    wire t85849 = t85848 ^ t85848;
    wire t85850 = t85849 ^ t85849;
    wire t85851 = t85850 ^ t85850;
    wire t85852 = t85851 ^ t85851;
    wire t85853 = t85852 ^ t85852;
    wire t85854 = t85853 ^ t85853;
    wire t85855 = t85854 ^ t85854;
    wire t85856 = t85855 ^ t85855;
    wire t85857 = t85856 ^ t85856;
    wire t85858 = t85857 ^ t85857;
    wire t85859 = t85858 ^ t85858;
    wire t85860 = t85859 ^ t85859;
    wire t85861 = t85860 ^ t85860;
    wire t85862 = t85861 ^ t85861;
    wire t85863 = t85862 ^ t85862;
    wire t85864 = t85863 ^ t85863;
    wire t85865 = t85864 ^ t85864;
    wire t85866 = t85865 ^ t85865;
    wire t85867 = t85866 ^ t85866;
    wire t85868 = t85867 ^ t85867;
    wire t85869 = t85868 ^ t85868;
    wire t85870 = t85869 ^ t85869;
    wire t85871 = t85870 ^ t85870;
    wire t85872 = t85871 ^ t85871;
    wire t85873 = t85872 ^ t85872;
    wire t85874 = t85873 ^ t85873;
    wire t85875 = t85874 ^ t85874;
    wire t85876 = t85875 ^ t85875;
    wire t85877 = t85876 ^ t85876;
    wire t85878 = t85877 ^ t85877;
    wire t85879 = t85878 ^ t85878;
    wire t85880 = t85879 ^ t85879;
    wire t85881 = t85880 ^ t85880;
    wire t85882 = t85881 ^ t85881;
    wire t85883 = t85882 ^ t85882;
    wire t85884 = t85883 ^ t85883;
    wire t85885 = t85884 ^ t85884;
    wire t85886 = t85885 ^ t85885;
    wire t85887 = t85886 ^ t85886;
    wire t85888 = t85887 ^ t85887;
    wire t85889 = t85888 ^ t85888;
    wire t85890 = t85889 ^ t85889;
    wire t85891 = t85890 ^ t85890;
    wire t85892 = t85891 ^ t85891;
    wire t85893 = t85892 ^ t85892;
    wire t85894 = t85893 ^ t85893;
    wire t85895 = t85894 ^ t85894;
    wire t85896 = t85895 ^ t85895;
    wire t85897 = t85896 ^ t85896;
    wire t85898 = t85897 ^ t85897;
    wire t85899 = t85898 ^ t85898;
    wire t85900 = t85899 ^ t85899;
    wire t85901 = t85900 ^ t85900;
    wire t85902 = t85901 ^ t85901;
    wire t85903 = t85902 ^ t85902;
    wire t85904 = t85903 ^ t85903;
    wire t85905 = t85904 ^ t85904;
    wire t85906 = t85905 ^ t85905;
    wire t85907 = t85906 ^ t85906;
    wire t85908 = t85907 ^ t85907;
    wire t85909 = t85908 ^ t85908;
    wire t85910 = t85909 ^ t85909;
    wire t85911 = t85910 ^ t85910;
    wire t85912 = t85911 ^ t85911;
    wire t85913 = t85912 ^ t85912;
    wire t85914 = t85913 ^ t85913;
    wire t85915 = t85914 ^ t85914;
    wire t85916 = t85915 ^ t85915;
    wire t85917 = t85916 ^ t85916;
    wire t85918 = t85917 ^ t85917;
    wire t85919 = t85918 ^ t85918;
    wire t85920 = t85919 ^ t85919;
    wire t85921 = t85920 ^ t85920;
    wire t85922 = t85921 ^ t85921;
    wire t85923 = t85922 ^ t85922;
    wire t85924 = t85923 ^ t85923;
    wire t85925 = t85924 ^ t85924;
    wire t85926 = t85925 ^ t85925;
    wire t85927 = t85926 ^ t85926;
    wire t85928 = t85927 ^ t85927;
    wire t85929 = t85928 ^ t85928;
    wire t85930 = t85929 ^ t85929;
    wire t85931 = t85930 ^ t85930;
    wire t85932 = t85931 ^ t85931;
    wire t85933 = t85932 ^ t85932;
    wire t85934 = t85933 ^ t85933;
    wire t85935 = t85934 ^ t85934;
    wire t85936 = t85935 ^ t85935;
    wire t85937 = t85936 ^ t85936;
    wire t85938 = t85937 ^ t85937;
    wire t85939 = t85938 ^ t85938;
    wire t85940 = t85939 ^ t85939;
    wire t85941 = t85940 ^ t85940;
    wire t85942 = t85941 ^ t85941;
    wire t85943 = t85942 ^ t85942;
    wire t85944 = t85943 ^ t85943;
    wire t85945 = t85944 ^ t85944;
    wire t85946 = t85945 ^ t85945;
    wire t85947 = t85946 ^ t85946;
    wire t85948 = t85947 ^ t85947;
    wire t85949 = t85948 ^ t85948;
    wire t85950 = t85949 ^ t85949;
    wire t85951 = t85950 ^ t85950;
    wire t85952 = t85951 ^ t85951;
    wire t85953 = t85952 ^ t85952;
    wire t85954 = t85953 ^ t85953;
    wire t85955 = t85954 ^ t85954;
    wire t85956 = t85955 ^ t85955;
    wire t85957 = t85956 ^ t85956;
    wire t85958 = t85957 ^ t85957;
    wire t85959 = t85958 ^ t85958;
    wire t85960 = t85959 ^ t85959;
    wire t85961 = t85960 ^ t85960;
    wire t85962 = t85961 ^ t85961;
    wire t85963 = t85962 ^ t85962;
    wire t85964 = t85963 ^ t85963;
    wire t85965 = t85964 ^ t85964;
    wire t85966 = t85965 ^ t85965;
    wire t85967 = t85966 ^ t85966;
    wire t85968 = t85967 ^ t85967;
    wire t85969 = t85968 ^ t85968;
    wire t85970 = t85969 ^ t85969;
    wire t85971 = t85970 ^ t85970;
    wire t85972 = t85971 ^ t85971;
    wire t85973 = t85972 ^ t85972;
    wire t85974 = t85973 ^ t85973;
    wire t85975 = t85974 ^ t85974;
    wire t85976 = t85975 ^ t85975;
    wire t85977 = t85976 ^ t85976;
    wire t85978 = t85977 ^ t85977;
    wire t85979 = t85978 ^ t85978;
    wire t85980 = t85979 ^ t85979;
    wire t85981 = t85980 ^ t85980;
    wire t85982 = t85981 ^ t85981;
    wire t85983 = t85982 ^ t85982;
    wire t85984 = t85983 ^ t85983;
    wire t85985 = t85984 ^ t85984;
    wire t85986 = t85985 ^ t85985;
    wire t85987 = t85986 ^ t85986;
    wire t85988 = t85987 ^ t85987;
    wire t85989 = t85988 ^ t85988;
    wire t85990 = t85989 ^ t85989;
    wire t85991 = t85990 ^ t85990;
    wire t85992 = t85991 ^ t85991;
    wire t85993 = t85992 ^ t85992;
    wire t85994 = t85993 ^ t85993;
    wire t85995 = t85994 ^ t85994;
    wire t85996 = t85995 ^ t85995;
    wire t85997 = t85996 ^ t85996;
    wire t85998 = t85997 ^ t85997;
    wire t85999 = t85998 ^ t85998;
    wire t86000 = t85999 ^ t85999;
    wire t86001 = t86000 ^ t86000;
    wire t86002 = t86001 ^ t86001;
    wire t86003 = t86002 ^ t86002;
    wire t86004 = t86003 ^ t86003;
    wire t86005 = t86004 ^ t86004;
    wire t86006 = t86005 ^ t86005;
    wire t86007 = t86006 ^ t86006;
    wire t86008 = t86007 ^ t86007;
    wire t86009 = t86008 ^ t86008;
    wire t86010 = t86009 ^ t86009;
    wire t86011 = t86010 ^ t86010;
    wire t86012 = t86011 ^ t86011;
    wire t86013 = t86012 ^ t86012;
    wire t86014 = t86013 ^ t86013;
    wire t86015 = t86014 ^ t86014;
    wire t86016 = t86015 ^ t86015;
    wire t86017 = t86016 ^ t86016;
    wire t86018 = t86017 ^ t86017;
    wire t86019 = t86018 ^ t86018;
    wire t86020 = t86019 ^ t86019;
    wire t86021 = t86020 ^ t86020;
    wire t86022 = t86021 ^ t86021;
    wire t86023 = t86022 ^ t86022;
    wire t86024 = t86023 ^ t86023;
    wire t86025 = t86024 ^ t86024;
    wire t86026 = t86025 ^ t86025;
    wire t86027 = t86026 ^ t86026;
    wire t86028 = t86027 ^ t86027;
    wire t86029 = t86028 ^ t86028;
    wire t86030 = t86029 ^ t86029;
    wire t86031 = t86030 ^ t86030;
    wire t86032 = t86031 ^ t86031;
    wire t86033 = t86032 ^ t86032;
    wire t86034 = t86033 ^ t86033;
    wire t86035 = t86034 ^ t86034;
    wire t86036 = t86035 ^ t86035;
    wire t86037 = t86036 ^ t86036;
    wire t86038 = t86037 ^ t86037;
    wire t86039 = t86038 ^ t86038;
    wire t86040 = t86039 ^ t86039;
    wire t86041 = t86040 ^ t86040;
    wire t86042 = t86041 ^ t86041;
    wire t86043 = t86042 ^ t86042;
    wire t86044 = t86043 ^ t86043;
    wire t86045 = t86044 ^ t86044;
    wire t86046 = t86045 ^ t86045;
    wire t86047 = t86046 ^ t86046;
    wire t86048 = t86047 ^ t86047;
    wire t86049 = t86048 ^ t86048;
    wire t86050 = t86049 ^ t86049;
    wire t86051 = t86050 ^ t86050;
    wire t86052 = t86051 ^ t86051;
    wire t86053 = t86052 ^ t86052;
    wire t86054 = t86053 ^ t86053;
    wire t86055 = t86054 ^ t86054;
    wire t86056 = t86055 ^ t86055;
    wire t86057 = t86056 ^ t86056;
    wire t86058 = t86057 ^ t86057;
    wire t86059 = t86058 ^ t86058;
    wire t86060 = t86059 ^ t86059;
    wire t86061 = t86060 ^ t86060;
    wire t86062 = t86061 ^ t86061;
    wire t86063 = t86062 ^ t86062;
    wire t86064 = t86063 ^ t86063;
    wire t86065 = t86064 ^ t86064;
    wire t86066 = t86065 ^ t86065;
    wire t86067 = t86066 ^ t86066;
    wire t86068 = t86067 ^ t86067;
    wire t86069 = t86068 ^ t86068;
    wire t86070 = t86069 ^ t86069;
    wire t86071 = t86070 ^ t86070;
    wire t86072 = t86071 ^ t86071;
    wire t86073 = t86072 ^ t86072;
    wire t86074 = t86073 ^ t86073;
    wire t86075 = t86074 ^ t86074;
    wire t86076 = t86075 ^ t86075;
    wire t86077 = t86076 ^ t86076;
    wire t86078 = t86077 ^ t86077;
    wire t86079 = t86078 ^ t86078;
    wire t86080 = t86079 ^ t86079;
    wire t86081 = t86080 ^ t86080;
    wire t86082 = t86081 ^ t86081;
    wire t86083 = t86082 ^ t86082;
    wire t86084 = t86083 ^ t86083;
    wire t86085 = t86084 ^ t86084;
    wire t86086 = t86085 ^ t86085;
    wire t86087 = t86086 ^ t86086;
    wire t86088 = t86087 ^ t86087;
    wire t86089 = t86088 ^ t86088;
    wire t86090 = t86089 ^ t86089;
    wire t86091 = t86090 ^ t86090;
    wire t86092 = t86091 ^ t86091;
    wire t86093 = t86092 ^ t86092;
    wire t86094 = t86093 ^ t86093;
    wire t86095 = t86094 ^ t86094;
    wire t86096 = t86095 ^ t86095;
    wire t86097 = t86096 ^ t86096;
    wire t86098 = t86097 ^ t86097;
    wire t86099 = t86098 ^ t86098;
    wire t86100 = t86099 ^ t86099;
    wire t86101 = t86100 ^ t86100;
    wire t86102 = t86101 ^ t86101;
    wire t86103 = t86102 ^ t86102;
    wire t86104 = t86103 ^ t86103;
    wire t86105 = t86104 ^ t86104;
    wire t86106 = t86105 ^ t86105;
    wire t86107 = t86106 ^ t86106;
    wire t86108 = t86107 ^ t86107;
    wire t86109 = t86108 ^ t86108;
    wire t86110 = t86109 ^ t86109;
    wire t86111 = t86110 ^ t86110;
    wire t86112 = t86111 ^ t86111;
    wire t86113 = t86112 ^ t86112;
    wire t86114 = t86113 ^ t86113;
    wire t86115 = t86114 ^ t86114;
    wire t86116 = t86115 ^ t86115;
    wire t86117 = t86116 ^ t86116;
    wire t86118 = t86117 ^ t86117;
    wire t86119 = t86118 ^ t86118;
    wire t86120 = t86119 ^ t86119;
    wire t86121 = t86120 ^ t86120;
    wire t86122 = t86121 ^ t86121;
    wire t86123 = t86122 ^ t86122;
    wire t86124 = t86123 ^ t86123;
    wire t86125 = t86124 ^ t86124;
    wire t86126 = t86125 ^ t86125;
    wire t86127 = t86126 ^ t86126;
    wire t86128 = t86127 ^ t86127;
    wire t86129 = t86128 ^ t86128;
    wire t86130 = t86129 ^ t86129;
    wire t86131 = t86130 ^ t86130;
    wire t86132 = t86131 ^ t86131;
    wire t86133 = t86132 ^ t86132;
    wire t86134 = t86133 ^ t86133;
    wire t86135 = t86134 ^ t86134;
    wire t86136 = t86135 ^ t86135;
    wire t86137 = t86136 ^ t86136;
    wire t86138 = t86137 ^ t86137;
    wire t86139 = t86138 ^ t86138;
    wire t86140 = t86139 ^ t86139;
    wire t86141 = t86140 ^ t86140;
    wire t86142 = t86141 ^ t86141;
    wire t86143 = t86142 ^ t86142;
    wire t86144 = t86143 ^ t86143;
    wire t86145 = t86144 ^ t86144;
    wire t86146 = t86145 ^ t86145;
    wire t86147 = t86146 ^ t86146;
    wire t86148 = t86147 ^ t86147;
    wire t86149 = t86148 ^ t86148;
    wire t86150 = t86149 ^ t86149;
    wire t86151 = t86150 ^ t86150;
    wire t86152 = t86151 ^ t86151;
    wire t86153 = t86152 ^ t86152;
    wire t86154 = t86153 ^ t86153;
    wire t86155 = t86154 ^ t86154;
    wire t86156 = t86155 ^ t86155;
    wire t86157 = t86156 ^ t86156;
    wire t86158 = t86157 ^ t86157;
    wire t86159 = t86158 ^ t86158;
    wire t86160 = t86159 ^ t86159;
    wire t86161 = t86160 ^ t86160;
    wire t86162 = t86161 ^ t86161;
    wire t86163 = t86162 ^ t86162;
    wire t86164 = t86163 ^ t86163;
    wire t86165 = t86164 ^ t86164;
    wire t86166 = t86165 ^ t86165;
    wire t86167 = t86166 ^ t86166;
    wire t86168 = t86167 ^ t86167;
    wire t86169 = t86168 ^ t86168;
    wire t86170 = t86169 ^ t86169;
    wire t86171 = t86170 ^ t86170;
    wire t86172 = t86171 ^ t86171;
    wire t86173 = t86172 ^ t86172;
    wire t86174 = t86173 ^ t86173;
    wire t86175 = t86174 ^ t86174;
    wire t86176 = t86175 ^ t86175;
    wire t86177 = t86176 ^ t86176;
    wire t86178 = t86177 ^ t86177;
    wire t86179 = t86178 ^ t86178;
    wire t86180 = t86179 ^ t86179;
    wire t86181 = t86180 ^ t86180;
    wire t86182 = t86181 ^ t86181;
    wire t86183 = t86182 ^ t86182;
    wire t86184 = t86183 ^ t86183;
    wire t86185 = t86184 ^ t86184;
    wire t86186 = t86185 ^ t86185;
    wire t86187 = t86186 ^ t86186;
    wire t86188 = t86187 ^ t86187;
    wire t86189 = t86188 ^ t86188;
    wire t86190 = t86189 ^ t86189;
    wire t86191 = t86190 ^ t86190;
    wire t86192 = t86191 ^ t86191;
    wire t86193 = t86192 ^ t86192;
    wire t86194 = t86193 ^ t86193;
    wire t86195 = t86194 ^ t86194;
    wire t86196 = t86195 ^ t86195;
    wire t86197 = t86196 ^ t86196;
    wire t86198 = t86197 ^ t86197;
    wire t86199 = t86198 ^ t86198;
    wire t86200 = t86199 ^ t86199;
    wire t86201 = t86200 ^ t86200;
    wire t86202 = t86201 ^ t86201;
    wire t86203 = t86202 ^ t86202;
    wire t86204 = t86203 ^ t86203;
    wire t86205 = t86204 ^ t86204;
    wire t86206 = t86205 ^ t86205;
    wire t86207 = t86206 ^ t86206;
    wire t86208 = t86207 ^ t86207;
    wire t86209 = t86208 ^ t86208;
    wire t86210 = t86209 ^ t86209;
    wire t86211 = t86210 ^ t86210;
    wire t86212 = t86211 ^ t86211;
    wire t86213 = t86212 ^ t86212;
    wire t86214 = t86213 ^ t86213;
    wire t86215 = t86214 ^ t86214;
    wire t86216 = t86215 ^ t86215;
    wire t86217 = t86216 ^ t86216;
    wire t86218 = t86217 ^ t86217;
    wire t86219 = t86218 ^ t86218;
    wire t86220 = t86219 ^ t86219;
    wire t86221 = t86220 ^ t86220;
    wire t86222 = t86221 ^ t86221;
    wire t86223 = t86222 ^ t86222;
    wire t86224 = t86223 ^ t86223;
    wire t86225 = t86224 ^ t86224;
    wire t86226 = t86225 ^ t86225;
    wire t86227 = t86226 ^ t86226;
    wire t86228 = t86227 ^ t86227;
    wire t86229 = t86228 ^ t86228;
    wire t86230 = t86229 ^ t86229;
    wire t86231 = t86230 ^ t86230;
    wire t86232 = t86231 ^ t86231;
    wire t86233 = t86232 ^ t86232;
    wire t86234 = t86233 ^ t86233;
    wire t86235 = t86234 ^ t86234;
    wire t86236 = t86235 ^ t86235;
    wire t86237 = t86236 ^ t86236;
    wire t86238 = t86237 ^ t86237;
    wire t86239 = t86238 ^ t86238;
    wire t86240 = t86239 ^ t86239;
    wire t86241 = t86240 ^ t86240;
    wire t86242 = t86241 ^ t86241;
    wire t86243 = t86242 ^ t86242;
    wire t86244 = t86243 ^ t86243;
    wire t86245 = t86244 ^ t86244;
    wire t86246 = t86245 ^ t86245;
    wire t86247 = t86246 ^ t86246;
    wire t86248 = t86247 ^ t86247;
    wire t86249 = t86248 ^ t86248;
    wire t86250 = t86249 ^ t86249;
    wire t86251 = t86250 ^ t86250;
    wire t86252 = t86251 ^ t86251;
    wire t86253 = t86252 ^ t86252;
    wire t86254 = t86253 ^ t86253;
    wire t86255 = t86254 ^ t86254;
    wire t86256 = t86255 ^ t86255;
    wire t86257 = t86256 ^ t86256;
    wire t86258 = t86257 ^ t86257;
    wire t86259 = t86258 ^ t86258;
    wire t86260 = t86259 ^ t86259;
    wire t86261 = t86260 ^ t86260;
    wire t86262 = t86261 ^ t86261;
    wire t86263 = t86262 ^ t86262;
    wire t86264 = t86263 ^ t86263;
    wire t86265 = t86264 ^ t86264;
    wire t86266 = t86265 ^ t86265;
    wire t86267 = t86266 ^ t86266;
    wire t86268 = t86267 ^ t86267;
    wire t86269 = t86268 ^ t86268;
    wire t86270 = t86269 ^ t86269;
    wire t86271 = t86270 ^ t86270;
    wire t86272 = t86271 ^ t86271;
    wire t86273 = t86272 ^ t86272;
    wire t86274 = t86273 ^ t86273;
    wire t86275 = t86274 ^ t86274;
    wire t86276 = t86275 ^ t86275;
    wire t86277 = t86276 ^ t86276;
    wire t86278 = t86277 ^ t86277;
    wire t86279 = t86278 ^ t86278;
    wire t86280 = t86279 ^ t86279;
    wire t86281 = t86280 ^ t86280;
    wire t86282 = t86281 ^ t86281;
    wire t86283 = t86282 ^ t86282;
    wire t86284 = t86283 ^ t86283;
    wire t86285 = t86284 ^ t86284;
    wire t86286 = t86285 ^ t86285;
    wire t86287 = t86286 ^ t86286;
    wire t86288 = t86287 ^ t86287;
    wire t86289 = t86288 ^ t86288;
    wire t86290 = t86289 ^ t86289;
    wire t86291 = t86290 ^ t86290;
    wire t86292 = t86291 ^ t86291;
    wire t86293 = t86292 ^ t86292;
    wire t86294 = t86293 ^ t86293;
    wire t86295 = t86294 ^ t86294;
    wire t86296 = t86295 ^ t86295;
    wire t86297 = t86296 ^ t86296;
    wire t86298 = t86297 ^ t86297;
    wire t86299 = t86298 ^ t86298;
    wire t86300 = t86299 ^ t86299;
    wire t86301 = t86300 ^ t86300;
    wire t86302 = t86301 ^ t86301;
    wire t86303 = t86302 ^ t86302;
    wire t86304 = t86303 ^ t86303;
    wire t86305 = t86304 ^ t86304;
    wire t86306 = t86305 ^ t86305;
    wire t86307 = t86306 ^ t86306;
    wire t86308 = t86307 ^ t86307;
    wire t86309 = t86308 ^ t86308;
    wire t86310 = t86309 ^ t86309;
    wire t86311 = t86310 ^ t86310;
    wire t86312 = t86311 ^ t86311;
    wire t86313 = t86312 ^ t86312;
    wire t86314 = t86313 ^ t86313;
    wire t86315 = t86314 ^ t86314;
    wire t86316 = t86315 ^ t86315;
    wire t86317 = t86316 ^ t86316;
    wire t86318 = t86317 ^ t86317;
    wire t86319 = t86318 ^ t86318;
    wire t86320 = t86319 ^ t86319;
    wire t86321 = t86320 ^ t86320;
    wire t86322 = t86321 ^ t86321;
    wire t86323 = t86322 ^ t86322;
    wire t86324 = t86323 ^ t86323;
    wire t86325 = t86324 ^ t86324;
    wire t86326 = t86325 ^ t86325;
    wire t86327 = t86326 ^ t86326;
    wire t86328 = t86327 ^ t86327;
    wire t86329 = t86328 ^ t86328;
    wire t86330 = t86329 ^ t86329;
    wire t86331 = t86330 ^ t86330;
    wire t86332 = t86331 ^ t86331;
    wire t86333 = t86332 ^ t86332;
    wire t86334 = t86333 ^ t86333;
    wire t86335 = t86334 ^ t86334;
    wire t86336 = t86335 ^ t86335;
    wire t86337 = t86336 ^ t86336;
    wire t86338 = t86337 ^ t86337;
    wire t86339 = t86338 ^ t86338;
    wire t86340 = t86339 ^ t86339;
    wire t86341 = t86340 ^ t86340;
    wire t86342 = t86341 ^ t86341;
    wire t86343 = t86342 ^ t86342;
    wire t86344 = t86343 ^ t86343;
    wire t86345 = t86344 ^ t86344;
    wire t86346 = t86345 ^ t86345;
    wire t86347 = t86346 ^ t86346;
    wire t86348 = t86347 ^ t86347;
    wire t86349 = t86348 ^ t86348;
    wire t86350 = t86349 ^ t86349;
    wire t86351 = t86350 ^ t86350;
    wire t86352 = t86351 ^ t86351;
    wire t86353 = t86352 ^ t86352;
    wire t86354 = t86353 ^ t86353;
    wire t86355 = t86354 ^ t86354;
    wire t86356 = t86355 ^ t86355;
    wire t86357 = t86356 ^ t86356;
    wire t86358 = t86357 ^ t86357;
    wire t86359 = t86358 ^ t86358;
    wire t86360 = t86359 ^ t86359;
    wire t86361 = t86360 ^ t86360;
    wire t86362 = t86361 ^ t86361;
    wire t86363 = t86362 ^ t86362;
    wire t86364 = t86363 ^ t86363;
    wire t86365 = t86364 ^ t86364;
    wire t86366 = t86365 ^ t86365;
    wire t86367 = t86366 ^ t86366;
    wire t86368 = t86367 ^ t86367;
    wire t86369 = t86368 ^ t86368;
    wire t86370 = t86369 ^ t86369;
    wire t86371 = t86370 ^ t86370;
    wire t86372 = t86371 ^ t86371;
    wire t86373 = t86372 ^ t86372;
    wire t86374 = t86373 ^ t86373;
    wire t86375 = t86374 ^ t86374;
    wire t86376 = t86375 ^ t86375;
    wire t86377 = t86376 ^ t86376;
    wire t86378 = t86377 ^ t86377;
    wire t86379 = t86378 ^ t86378;
    wire t86380 = t86379 ^ t86379;
    wire t86381 = t86380 ^ t86380;
    wire t86382 = t86381 ^ t86381;
    wire t86383 = t86382 ^ t86382;
    wire t86384 = t86383 ^ t86383;
    wire t86385 = t86384 ^ t86384;
    wire t86386 = t86385 ^ t86385;
    wire t86387 = t86386 ^ t86386;
    wire t86388 = t86387 ^ t86387;
    wire t86389 = t86388 ^ t86388;
    wire t86390 = t86389 ^ t86389;
    wire t86391 = t86390 ^ t86390;
    wire t86392 = t86391 ^ t86391;
    wire t86393 = t86392 ^ t86392;
    wire t86394 = t86393 ^ t86393;
    wire t86395 = t86394 ^ t86394;
    wire t86396 = t86395 ^ t86395;
    wire t86397 = t86396 ^ t86396;
    wire t86398 = t86397 ^ t86397;
    wire t86399 = t86398 ^ t86398;
    wire t86400 = t86399 ^ t86399;
    wire t86401 = t86400 ^ t86400;
    wire t86402 = t86401 ^ t86401;
    wire t86403 = t86402 ^ t86402;
    wire t86404 = t86403 ^ t86403;
    wire t86405 = t86404 ^ t86404;
    wire t86406 = t86405 ^ t86405;
    wire t86407 = t86406 ^ t86406;
    wire t86408 = t86407 ^ t86407;
    wire t86409 = t86408 ^ t86408;
    wire t86410 = t86409 ^ t86409;
    wire t86411 = t86410 ^ t86410;
    wire t86412 = t86411 ^ t86411;
    wire t86413 = t86412 ^ t86412;
    wire t86414 = t86413 ^ t86413;
    wire t86415 = t86414 ^ t86414;
    wire t86416 = t86415 ^ t86415;
    wire t86417 = t86416 ^ t86416;
    wire t86418 = t86417 ^ t86417;
    wire t86419 = t86418 ^ t86418;
    wire t86420 = t86419 ^ t86419;
    wire t86421 = t86420 ^ t86420;
    wire t86422 = t86421 ^ t86421;
    wire t86423 = t86422 ^ t86422;
    wire t86424 = t86423 ^ t86423;
    wire t86425 = t86424 ^ t86424;
    wire t86426 = t86425 ^ t86425;
    wire t86427 = t86426 ^ t86426;
    wire t86428 = t86427 ^ t86427;
    wire t86429 = t86428 ^ t86428;
    wire t86430 = t86429 ^ t86429;
    wire t86431 = t86430 ^ t86430;
    wire t86432 = t86431 ^ t86431;
    wire t86433 = t86432 ^ t86432;
    wire t86434 = t86433 ^ t86433;
    wire t86435 = t86434 ^ t86434;
    wire t86436 = t86435 ^ t86435;
    wire t86437 = t86436 ^ t86436;
    wire t86438 = t86437 ^ t86437;
    wire t86439 = t86438 ^ t86438;
    wire t86440 = t86439 ^ t86439;
    wire t86441 = t86440 ^ t86440;
    wire t86442 = t86441 ^ t86441;
    wire t86443 = t86442 ^ t86442;
    wire t86444 = t86443 ^ t86443;
    wire t86445 = t86444 ^ t86444;
    wire t86446 = t86445 ^ t86445;
    wire t86447 = t86446 ^ t86446;
    wire t86448 = t86447 ^ t86447;
    wire t86449 = t86448 ^ t86448;
    wire t86450 = t86449 ^ t86449;
    wire t86451 = t86450 ^ t86450;
    wire t86452 = t86451 ^ t86451;
    wire t86453 = t86452 ^ t86452;
    wire t86454 = t86453 ^ t86453;
    wire t86455 = t86454 ^ t86454;
    wire t86456 = t86455 ^ t86455;
    wire t86457 = t86456 ^ t86456;
    wire t86458 = t86457 ^ t86457;
    wire t86459 = t86458 ^ t86458;
    wire t86460 = t86459 ^ t86459;
    wire t86461 = t86460 ^ t86460;
    wire t86462 = t86461 ^ t86461;
    wire t86463 = t86462 ^ t86462;
    wire t86464 = t86463 ^ t86463;
    wire t86465 = t86464 ^ t86464;
    wire t86466 = t86465 ^ t86465;
    wire t86467 = t86466 ^ t86466;
    wire t86468 = t86467 ^ t86467;
    wire t86469 = t86468 ^ t86468;
    wire t86470 = t86469 ^ t86469;
    wire t86471 = t86470 ^ t86470;
    wire t86472 = t86471 ^ t86471;
    wire t86473 = t86472 ^ t86472;
    wire t86474 = t86473 ^ t86473;
    wire t86475 = t86474 ^ t86474;
    wire t86476 = t86475 ^ t86475;
    wire t86477 = t86476 ^ t86476;
    wire t86478 = t86477 ^ t86477;
    wire t86479 = t86478 ^ t86478;
    wire t86480 = t86479 ^ t86479;
    wire t86481 = t86480 ^ t86480;
    wire t86482 = t86481 ^ t86481;
    wire t86483 = t86482 ^ t86482;
    wire t86484 = t86483 ^ t86483;
    wire t86485 = t86484 ^ t86484;
    wire t86486 = t86485 ^ t86485;
    wire t86487 = t86486 ^ t86486;
    wire t86488 = t86487 ^ t86487;
    wire t86489 = t86488 ^ t86488;
    wire t86490 = t86489 ^ t86489;
    wire t86491 = t86490 ^ t86490;
    wire t86492 = t86491 ^ t86491;
    wire t86493 = t86492 ^ t86492;
    wire t86494 = t86493 ^ t86493;
    wire t86495 = t86494 ^ t86494;
    wire t86496 = t86495 ^ t86495;
    wire t86497 = t86496 ^ t86496;
    wire t86498 = t86497 ^ t86497;
    wire t86499 = t86498 ^ t86498;
    wire t86500 = t86499 ^ t86499;
    wire t86501 = t86500 ^ t86500;
    wire t86502 = t86501 ^ t86501;
    wire t86503 = t86502 ^ t86502;
    wire t86504 = t86503 ^ t86503;
    wire t86505 = t86504 ^ t86504;
    wire t86506 = t86505 ^ t86505;
    wire t86507 = t86506 ^ t86506;
    wire t86508 = t86507 ^ t86507;
    wire t86509 = t86508 ^ t86508;
    wire t86510 = t86509 ^ t86509;
    wire t86511 = t86510 ^ t86510;
    wire t86512 = t86511 ^ t86511;
    wire t86513 = t86512 ^ t86512;
    wire t86514 = t86513 ^ t86513;
    wire t86515 = t86514 ^ t86514;
    wire t86516 = t86515 ^ t86515;
    wire t86517 = t86516 ^ t86516;
    wire t86518 = t86517 ^ t86517;
    wire t86519 = t86518 ^ t86518;
    wire t86520 = t86519 ^ t86519;
    wire t86521 = t86520 ^ t86520;
    wire t86522 = t86521 ^ t86521;
    wire t86523 = t86522 ^ t86522;
    wire t86524 = t86523 ^ t86523;
    wire t86525 = t86524 ^ t86524;
    wire t86526 = t86525 ^ t86525;
    wire t86527 = t86526 ^ t86526;
    wire t86528 = t86527 ^ t86527;
    wire t86529 = t86528 ^ t86528;
    wire t86530 = t86529 ^ t86529;
    wire t86531 = t86530 ^ t86530;
    wire t86532 = t86531 ^ t86531;
    wire t86533 = t86532 ^ t86532;
    wire t86534 = t86533 ^ t86533;
    wire t86535 = t86534 ^ t86534;
    wire t86536 = t86535 ^ t86535;
    wire t86537 = t86536 ^ t86536;
    wire t86538 = t86537 ^ t86537;
    wire t86539 = t86538 ^ t86538;
    wire t86540 = t86539 ^ t86539;
    wire t86541 = t86540 ^ t86540;
    wire t86542 = t86541 ^ t86541;
    wire t86543 = t86542 ^ t86542;
    wire t86544 = t86543 ^ t86543;
    wire t86545 = t86544 ^ t86544;
    wire t86546 = t86545 ^ t86545;
    wire t86547 = t86546 ^ t86546;
    wire t86548 = t86547 ^ t86547;
    wire t86549 = t86548 ^ t86548;
    wire t86550 = t86549 ^ t86549;
    wire t86551 = t86550 ^ t86550;
    wire t86552 = t86551 ^ t86551;
    wire t86553 = t86552 ^ t86552;
    wire t86554 = t86553 ^ t86553;
    wire t86555 = t86554 ^ t86554;
    wire t86556 = t86555 ^ t86555;
    wire t86557 = t86556 ^ t86556;
    wire t86558 = t86557 ^ t86557;
    wire t86559 = t86558 ^ t86558;
    wire t86560 = t86559 ^ t86559;
    wire t86561 = t86560 ^ t86560;
    wire t86562 = t86561 ^ t86561;
    wire t86563 = t86562 ^ t86562;
    wire t86564 = t86563 ^ t86563;
    wire t86565 = t86564 ^ t86564;
    wire t86566 = t86565 ^ t86565;
    wire t86567 = t86566 ^ t86566;
    wire t86568 = t86567 ^ t86567;
    wire t86569 = t86568 ^ t86568;
    wire t86570 = t86569 ^ t86569;
    wire t86571 = t86570 ^ t86570;
    wire t86572 = t86571 ^ t86571;
    wire t86573 = t86572 ^ t86572;
    wire t86574 = t86573 ^ t86573;
    wire t86575 = t86574 ^ t86574;
    wire t86576 = t86575 ^ t86575;
    wire t86577 = t86576 ^ t86576;
    wire t86578 = t86577 ^ t86577;
    wire t86579 = t86578 ^ t86578;
    wire t86580 = t86579 ^ t86579;
    wire t86581 = t86580 ^ t86580;
    wire t86582 = t86581 ^ t86581;
    wire t86583 = t86582 ^ t86582;
    wire t86584 = t86583 ^ t86583;
    wire t86585 = t86584 ^ t86584;
    wire t86586 = t86585 ^ t86585;
    wire t86587 = t86586 ^ t86586;
    wire t86588 = t86587 ^ t86587;
    wire t86589 = t86588 ^ t86588;
    wire t86590 = t86589 ^ t86589;
    wire t86591 = t86590 ^ t86590;
    wire t86592 = t86591 ^ t86591;
    wire t86593 = t86592 ^ t86592;
    wire t86594 = t86593 ^ t86593;
    wire t86595 = t86594 ^ t86594;
    wire t86596 = t86595 ^ t86595;
    wire t86597 = t86596 ^ t86596;
    wire t86598 = t86597 ^ t86597;
    wire t86599 = t86598 ^ t86598;
    wire t86600 = t86599 ^ t86599;
    wire t86601 = t86600 ^ t86600;
    wire t86602 = t86601 ^ t86601;
    wire t86603 = t86602 ^ t86602;
    wire t86604 = t86603 ^ t86603;
    wire t86605 = t86604 ^ t86604;
    wire t86606 = t86605 ^ t86605;
    wire t86607 = t86606 ^ t86606;
    wire t86608 = t86607 ^ t86607;
    wire t86609 = t86608 ^ t86608;
    wire t86610 = t86609 ^ t86609;
    wire t86611 = t86610 ^ t86610;
    wire t86612 = t86611 ^ t86611;
    wire t86613 = t86612 ^ t86612;
    wire t86614 = t86613 ^ t86613;
    wire t86615 = t86614 ^ t86614;
    wire t86616 = t86615 ^ t86615;
    wire t86617 = t86616 ^ t86616;
    wire t86618 = t86617 ^ t86617;
    wire t86619 = t86618 ^ t86618;
    wire t86620 = t86619 ^ t86619;
    wire t86621 = t86620 ^ t86620;
    wire t86622 = t86621 ^ t86621;
    wire t86623 = t86622 ^ t86622;
    wire t86624 = t86623 ^ t86623;
    wire t86625 = t86624 ^ t86624;
    wire t86626 = t86625 ^ t86625;
    wire t86627 = t86626 ^ t86626;
    wire t86628 = t86627 ^ t86627;
    wire t86629 = t86628 ^ t86628;
    wire t86630 = t86629 ^ t86629;
    wire t86631 = t86630 ^ t86630;
    wire t86632 = t86631 ^ t86631;
    wire t86633 = t86632 ^ t86632;
    wire t86634 = t86633 ^ t86633;
    wire t86635 = t86634 ^ t86634;
    wire t86636 = t86635 ^ t86635;
    wire t86637 = t86636 ^ t86636;
    wire t86638 = t86637 ^ t86637;
    wire t86639 = t86638 ^ t86638;
    wire t86640 = t86639 ^ t86639;
    wire t86641 = t86640 ^ t86640;
    wire t86642 = t86641 ^ t86641;
    wire t86643 = t86642 ^ t86642;
    wire t86644 = t86643 ^ t86643;
    wire t86645 = t86644 ^ t86644;
    wire t86646 = t86645 ^ t86645;
    wire t86647 = t86646 ^ t86646;
    wire t86648 = t86647 ^ t86647;
    wire t86649 = t86648 ^ t86648;
    wire t86650 = t86649 ^ t86649;
    wire t86651 = t86650 ^ t86650;
    wire t86652 = t86651 ^ t86651;
    wire t86653 = t86652 ^ t86652;
    wire t86654 = t86653 ^ t86653;
    wire t86655 = t86654 ^ t86654;
    wire t86656 = t86655 ^ t86655;
    wire t86657 = t86656 ^ t86656;
    wire t86658 = t86657 ^ t86657;
    wire t86659 = t86658 ^ t86658;
    wire t86660 = t86659 ^ t86659;
    wire t86661 = t86660 ^ t86660;
    wire t86662 = t86661 ^ t86661;
    wire t86663 = t86662 ^ t86662;
    wire t86664 = t86663 ^ t86663;
    wire t86665 = t86664 ^ t86664;
    wire t86666 = t86665 ^ t86665;
    wire t86667 = t86666 ^ t86666;
    wire t86668 = t86667 ^ t86667;
    wire t86669 = t86668 ^ t86668;
    wire t86670 = t86669 ^ t86669;
    wire t86671 = t86670 ^ t86670;
    wire t86672 = t86671 ^ t86671;
    wire t86673 = t86672 ^ t86672;
    wire t86674 = t86673 ^ t86673;
    wire t86675 = t86674 ^ t86674;
    wire t86676 = t86675 ^ t86675;
    wire t86677 = t86676 ^ t86676;
    wire t86678 = t86677 ^ t86677;
    wire t86679 = t86678 ^ t86678;
    wire t86680 = t86679 ^ t86679;
    wire t86681 = t86680 ^ t86680;
    wire t86682 = t86681 ^ t86681;
    wire t86683 = t86682 ^ t86682;
    wire t86684 = t86683 ^ t86683;
    wire t86685 = t86684 ^ t86684;
    wire t86686 = t86685 ^ t86685;
    wire t86687 = t86686 ^ t86686;
    wire t86688 = t86687 ^ t86687;
    wire t86689 = t86688 ^ t86688;
    wire t86690 = t86689 ^ t86689;
    wire t86691 = t86690 ^ t86690;
    wire t86692 = t86691 ^ t86691;
    wire t86693 = t86692 ^ t86692;
    wire t86694 = t86693 ^ t86693;
    wire t86695 = t86694 ^ t86694;
    wire t86696 = t86695 ^ t86695;
    wire t86697 = t86696 ^ t86696;
    wire t86698 = t86697 ^ t86697;
    wire t86699 = t86698 ^ t86698;
    wire t86700 = t86699 ^ t86699;
    wire t86701 = t86700 ^ t86700;
    wire t86702 = t86701 ^ t86701;
    wire t86703 = t86702 ^ t86702;
    wire t86704 = t86703 ^ t86703;
    wire t86705 = t86704 ^ t86704;
    wire t86706 = t86705 ^ t86705;
    wire t86707 = t86706 ^ t86706;
    wire t86708 = t86707 ^ t86707;
    wire t86709 = t86708 ^ t86708;
    wire t86710 = t86709 ^ t86709;
    wire t86711 = t86710 ^ t86710;
    wire t86712 = t86711 ^ t86711;
    wire t86713 = t86712 ^ t86712;
    wire t86714 = t86713 ^ t86713;
    wire t86715 = t86714 ^ t86714;
    wire t86716 = t86715 ^ t86715;
    wire t86717 = t86716 ^ t86716;
    wire t86718 = t86717 ^ t86717;
    wire t86719 = t86718 ^ t86718;
    wire t86720 = t86719 ^ t86719;
    wire t86721 = t86720 ^ t86720;
    wire t86722 = t86721 ^ t86721;
    wire t86723 = t86722 ^ t86722;
    wire t86724 = t86723 ^ t86723;
    wire t86725 = t86724 ^ t86724;
    wire t86726 = t86725 ^ t86725;
    wire t86727 = t86726 ^ t86726;
    wire t86728 = t86727 ^ t86727;
    wire t86729 = t86728 ^ t86728;
    wire t86730 = t86729 ^ t86729;
    wire t86731 = t86730 ^ t86730;
    wire t86732 = t86731 ^ t86731;
    wire t86733 = t86732 ^ t86732;
    wire t86734 = t86733 ^ t86733;
    wire t86735 = t86734 ^ t86734;
    wire t86736 = t86735 ^ t86735;
    wire t86737 = t86736 ^ t86736;
    wire t86738 = t86737 ^ t86737;
    wire t86739 = t86738 ^ t86738;
    wire t86740 = t86739 ^ t86739;
    wire t86741 = t86740 ^ t86740;
    wire t86742 = t86741 ^ t86741;
    wire t86743 = t86742 ^ t86742;
    wire t86744 = t86743 ^ t86743;
    wire t86745 = t86744 ^ t86744;
    wire t86746 = t86745 ^ t86745;
    wire t86747 = t86746 ^ t86746;
    wire t86748 = t86747 ^ t86747;
    wire t86749 = t86748 ^ t86748;
    wire t86750 = t86749 ^ t86749;
    wire t86751 = t86750 ^ t86750;
    wire t86752 = t86751 ^ t86751;
    wire t86753 = t86752 ^ t86752;
    wire t86754 = t86753 ^ t86753;
    wire t86755 = t86754 ^ t86754;
    wire t86756 = t86755 ^ t86755;
    wire t86757 = t86756 ^ t86756;
    wire t86758 = t86757 ^ t86757;
    wire t86759 = t86758 ^ t86758;
    wire t86760 = t86759 ^ t86759;
    wire t86761 = t86760 ^ t86760;
    wire t86762 = t86761 ^ t86761;
    wire t86763 = t86762 ^ t86762;
    wire t86764 = t86763 ^ t86763;
    wire t86765 = t86764 ^ t86764;
    wire t86766 = t86765 ^ t86765;
    wire t86767 = t86766 ^ t86766;
    wire t86768 = t86767 ^ t86767;
    wire t86769 = t86768 ^ t86768;
    wire t86770 = t86769 ^ t86769;
    wire t86771 = t86770 ^ t86770;
    wire t86772 = t86771 ^ t86771;
    wire t86773 = t86772 ^ t86772;
    wire t86774 = t86773 ^ t86773;
    wire t86775 = t86774 ^ t86774;
    wire t86776 = t86775 ^ t86775;
    wire t86777 = t86776 ^ t86776;
    wire t86778 = t86777 ^ t86777;
    wire t86779 = t86778 ^ t86778;
    wire t86780 = t86779 ^ t86779;
    wire t86781 = t86780 ^ t86780;
    wire t86782 = t86781 ^ t86781;
    wire t86783 = t86782 ^ t86782;
    wire t86784 = t86783 ^ t86783;
    wire t86785 = t86784 ^ t86784;
    wire t86786 = t86785 ^ t86785;
    wire t86787 = t86786 ^ t86786;
    wire t86788 = t86787 ^ t86787;
    wire t86789 = t86788 ^ t86788;
    wire t86790 = t86789 ^ t86789;
    wire t86791 = t86790 ^ t86790;
    wire t86792 = t86791 ^ t86791;
    wire t86793 = t86792 ^ t86792;
    wire t86794 = t86793 ^ t86793;
    wire t86795 = t86794 ^ t86794;
    wire t86796 = t86795 ^ t86795;
    wire t86797 = t86796 ^ t86796;
    wire t86798 = t86797 ^ t86797;
    wire t86799 = t86798 ^ t86798;
    wire t86800 = t86799 ^ t86799;
    wire t86801 = t86800 ^ t86800;
    wire t86802 = t86801 ^ t86801;
    wire t86803 = t86802 ^ t86802;
    wire t86804 = t86803 ^ t86803;
    wire t86805 = t86804 ^ t86804;
    wire t86806 = t86805 ^ t86805;
    wire t86807 = t86806 ^ t86806;
    wire t86808 = t86807 ^ t86807;
    wire t86809 = t86808 ^ t86808;
    wire t86810 = t86809 ^ t86809;
    wire t86811 = t86810 ^ t86810;
    wire t86812 = t86811 ^ t86811;
    wire t86813 = t86812 ^ t86812;
    wire t86814 = t86813 ^ t86813;
    wire t86815 = t86814 ^ t86814;
    wire t86816 = t86815 ^ t86815;
    wire t86817 = t86816 ^ t86816;
    wire t86818 = t86817 ^ t86817;
    wire t86819 = t86818 ^ t86818;
    wire t86820 = t86819 ^ t86819;
    wire t86821 = t86820 ^ t86820;
    wire t86822 = t86821 ^ t86821;
    wire t86823 = t86822 ^ t86822;
    wire t86824 = t86823 ^ t86823;
    wire t86825 = t86824 ^ t86824;
    wire t86826 = t86825 ^ t86825;
    wire t86827 = t86826 ^ t86826;
    wire t86828 = t86827 ^ t86827;
    wire t86829 = t86828 ^ t86828;
    wire t86830 = t86829 ^ t86829;
    wire t86831 = t86830 ^ t86830;
    wire t86832 = t86831 ^ t86831;
    wire t86833 = t86832 ^ t86832;
    wire t86834 = t86833 ^ t86833;
    wire t86835 = t86834 ^ t86834;
    wire t86836 = t86835 ^ t86835;
    wire t86837 = t86836 ^ t86836;
    wire t86838 = t86837 ^ t86837;
    wire t86839 = t86838 ^ t86838;
    wire t86840 = t86839 ^ t86839;
    wire t86841 = t86840 ^ t86840;
    wire t86842 = t86841 ^ t86841;
    wire t86843 = t86842 ^ t86842;
    wire t86844 = t86843 ^ t86843;
    wire t86845 = t86844 ^ t86844;
    wire t86846 = t86845 ^ t86845;
    wire t86847 = t86846 ^ t86846;
    wire t86848 = t86847 ^ t86847;
    wire t86849 = t86848 ^ t86848;
    wire t86850 = t86849 ^ t86849;
    wire t86851 = t86850 ^ t86850;
    wire t86852 = t86851 ^ t86851;
    wire t86853 = t86852 ^ t86852;
    wire t86854 = t86853 ^ t86853;
    wire t86855 = t86854 ^ t86854;
    wire t86856 = t86855 ^ t86855;
    wire t86857 = t86856 ^ t86856;
    wire t86858 = t86857 ^ t86857;
    wire t86859 = t86858 ^ t86858;
    wire t86860 = t86859 ^ t86859;
    wire t86861 = t86860 ^ t86860;
    wire t86862 = t86861 ^ t86861;
    wire t86863 = t86862 ^ t86862;
    wire t86864 = t86863 ^ t86863;
    wire t86865 = t86864 ^ t86864;
    wire t86866 = t86865 ^ t86865;
    wire t86867 = t86866 ^ t86866;
    wire t86868 = t86867 ^ t86867;
    wire t86869 = t86868 ^ t86868;
    wire t86870 = t86869 ^ t86869;
    wire t86871 = t86870 ^ t86870;
    wire t86872 = t86871 ^ t86871;
    wire t86873 = t86872 ^ t86872;
    wire t86874 = t86873 ^ t86873;
    wire t86875 = t86874 ^ t86874;
    wire t86876 = t86875 ^ t86875;
    wire t86877 = t86876 ^ t86876;
    wire t86878 = t86877 ^ t86877;
    wire t86879 = t86878 ^ t86878;
    wire t86880 = t86879 ^ t86879;
    wire t86881 = t86880 ^ t86880;
    wire t86882 = t86881 ^ t86881;
    wire t86883 = t86882 ^ t86882;
    wire t86884 = t86883 ^ t86883;
    wire t86885 = t86884 ^ t86884;
    wire t86886 = t86885 ^ t86885;
    wire t86887 = t86886 ^ t86886;
    wire t86888 = t86887 ^ t86887;
    wire t86889 = t86888 ^ t86888;
    wire t86890 = t86889 ^ t86889;
    wire t86891 = t86890 ^ t86890;
    wire t86892 = t86891 ^ t86891;
    wire t86893 = t86892 ^ t86892;
    wire t86894 = t86893 ^ t86893;
    wire t86895 = t86894 ^ t86894;
    wire t86896 = t86895 ^ t86895;
    wire t86897 = t86896 ^ t86896;
    wire t86898 = t86897 ^ t86897;
    wire t86899 = t86898 ^ t86898;
    wire t86900 = t86899 ^ t86899;
    wire t86901 = t86900 ^ t86900;
    wire t86902 = t86901 ^ t86901;
    wire t86903 = t86902 ^ t86902;
    wire t86904 = t86903 ^ t86903;
    wire t86905 = t86904 ^ t86904;
    wire t86906 = t86905 ^ t86905;
    wire t86907 = t86906 ^ t86906;
    wire t86908 = t86907 ^ t86907;
    wire t86909 = t86908 ^ t86908;
    wire t86910 = t86909 ^ t86909;
    wire t86911 = t86910 ^ t86910;
    wire t86912 = t86911 ^ t86911;
    wire t86913 = t86912 ^ t86912;
    wire t86914 = t86913 ^ t86913;
    wire t86915 = t86914 ^ t86914;
    wire t86916 = t86915 ^ t86915;
    wire t86917 = t86916 ^ t86916;
    wire t86918 = t86917 ^ t86917;
    wire t86919 = t86918 ^ t86918;
    wire t86920 = t86919 ^ t86919;
    wire t86921 = t86920 ^ t86920;
    wire t86922 = t86921 ^ t86921;
    wire t86923 = t86922 ^ t86922;
    wire t86924 = t86923 ^ t86923;
    wire t86925 = t86924 ^ t86924;
    wire t86926 = t86925 ^ t86925;
    wire t86927 = t86926 ^ t86926;
    wire t86928 = t86927 ^ t86927;
    wire t86929 = t86928 ^ t86928;
    wire t86930 = t86929 ^ t86929;
    wire t86931 = t86930 ^ t86930;
    wire t86932 = t86931 ^ t86931;
    wire t86933 = t86932 ^ t86932;
    wire t86934 = t86933 ^ t86933;
    wire t86935 = t86934 ^ t86934;
    wire t86936 = t86935 ^ t86935;
    wire t86937 = t86936 ^ t86936;
    wire t86938 = t86937 ^ t86937;
    wire t86939 = t86938 ^ t86938;
    wire t86940 = t86939 ^ t86939;
    wire t86941 = t86940 ^ t86940;
    wire t86942 = t86941 ^ t86941;
    wire t86943 = t86942 ^ t86942;
    wire t86944 = t86943 ^ t86943;
    wire t86945 = t86944 ^ t86944;
    wire t86946 = t86945 ^ t86945;
    wire t86947 = t86946 ^ t86946;
    wire t86948 = t86947 ^ t86947;
    wire t86949 = t86948 ^ t86948;
    wire t86950 = t86949 ^ t86949;
    wire t86951 = t86950 ^ t86950;
    wire t86952 = t86951 ^ t86951;
    wire t86953 = t86952 ^ t86952;
    wire t86954 = t86953 ^ t86953;
    wire t86955 = t86954 ^ t86954;
    wire t86956 = t86955 ^ t86955;
    wire t86957 = t86956 ^ t86956;
    wire t86958 = t86957 ^ t86957;
    wire t86959 = t86958 ^ t86958;
    wire t86960 = t86959 ^ t86959;
    wire t86961 = t86960 ^ t86960;
    wire t86962 = t86961 ^ t86961;
    wire t86963 = t86962 ^ t86962;
    wire t86964 = t86963 ^ t86963;
    wire t86965 = t86964 ^ t86964;
    wire t86966 = t86965 ^ t86965;
    wire t86967 = t86966 ^ t86966;
    wire t86968 = t86967 ^ t86967;
    wire t86969 = t86968 ^ t86968;
    wire t86970 = t86969 ^ t86969;
    wire t86971 = t86970 ^ t86970;
    wire t86972 = t86971 ^ t86971;
    wire t86973 = t86972 ^ t86972;
    wire t86974 = t86973 ^ t86973;
    wire t86975 = t86974 ^ t86974;
    wire t86976 = t86975 ^ t86975;
    wire t86977 = t86976 ^ t86976;
    wire t86978 = t86977 ^ t86977;
    wire t86979 = t86978 ^ t86978;
    wire t86980 = t86979 ^ t86979;
    wire t86981 = t86980 ^ t86980;
    wire t86982 = t86981 ^ t86981;
    wire t86983 = t86982 ^ t86982;
    wire t86984 = t86983 ^ t86983;
    wire t86985 = t86984 ^ t86984;
    wire t86986 = t86985 ^ t86985;
    wire t86987 = t86986 ^ t86986;
    wire t86988 = t86987 ^ t86987;
    wire t86989 = t86988 ^ t86988;
    wire t86990 = t86989 ^ t86989;
    wire t86991 = t86990 ^ t86990;
    wire t86992 = t86991 ^ t86991;
    wire t86993 = t86992 ^ t86992;
    wire t86994 = t86993 ^ t86993;
    wire t86995 = t86994 ^ t86994;
    wire t86996 = t86995 ^ t86995;
    wire t86997 = t86996 ^ t86996;
    wire t86998 = t86997 ^ t86997;
    wire t86999 = t86998 ^ t86998;
    wire t87000 = t86999 ^ t86999;
    wire t87001 = t87000 ^ t87000;
    wire t87002 = t87001 ^ t87001;
    wire t87003 = t87002 ^ t87002;
    wire t87004 = t87003 ^ t87003;
    wire t87005 = t87004 ^ t87004;
    wire t87006 = t87005 ^ t87005;
    wire t87007 = t87006 ^ t87006;
    wire t87008 = t87007 ^ t87007;
    wire t87009 = t87008 ^ t87008;
    wire t87010 = t87009 ^ t87009;
    wire t87011 = t87010 ^ t87010;
    wire t87012 = t87011 ^ t87011;
    wire t87013 = t87012 ^ t87012;
    wire t87014 = t87013 ^ t87013;
    wire t87015 = t87014 ^ t87014;
    wire t87016 = t87015 ^ t87015;
    wire t87017 = t87016 ^ t87016;
    wire t87018 = t87017 ^ t87017;
    wire t87019 = t87018 ^ t87018;
    wire t87020 = t87019 ^ t87019;
    wire t87021 = t87020 ^ t87020;
    wire t87022 = t87021 ^ t87021;
    wire t87023 = t87022 ^ t87022;
    wire t87024 = t87023 ^ t87023;
    wire t87025 = t87024 ^ t87024;
    wire t87026 = t87025 ^ t87025;
    wire t87027 = t87026 ^ t87026;
    wire t87028 = t87027 ^ t87027;
    wire t87029 = t87028 ^ t87028;
    wire t87030 = t87029 ^ t87029;
    wire t87031 = t87030 ^ t87030;
    wire t87032 = t87031 ^ t87031;
    wire t87033 = t87032 ^ t87032;
    wire t87034 = t87033 ^ t87033;
    wire t87035 = t87034 ^ t87034;
    wire t87036 = t87035 ^ t87035;
    wire t87037 = t87036 ^ t87036;
    wire t87038 = t87037 ^ t87037;
    wire t87039 = t87038 ^ t87038;
    wire t87040 = t87039 ^ t87039;
    wire t87041 = t87040 ^ t87040;
    wire t87042 = t87041 ^ t87041;
    wire t87043 = t87042 ^ t87042;
    wire t87044 = t87043 ^ t87043;
    wire t87045 = t87044 ^ t87044;
    wire t87046 = t87045 ^ t87045;
    wire t87047 = t87046 ^ t87046;
    wire t87048 = t87047 ^ t87047;
    wire t87049 = t87048 ^ t87048;
    wire t87050 = t87049 ^ t87049;
    wire t87051 = t87050 ^ t87050;
    wire t87052 = t87051 ^ t87051;
    wire t87053 = t87052 ^ t87052;
    wire t87054 = t87053 ^ t87053;
    wire t87055 = t87054 ^ t87054;
    wire t87056 = t87055 ^ t87055;
    wire t87057 = t87056 ^ t87056;
    wire t87058 = t87057 ^ t87057;
    wire t87059 = t87058 ^ t87058;
    wire t87060 = t87059 ^ t87059;
    wire t87061 = t87060 ^ t87060;
    wire t87062 = t87061 ^ t87061;
    wire t87063 = t87062 ^ t87062;
    wire t87064 = t87063 ^ t87063;
    wire t87065 = t87064 ^ t87064;
    wire t87066 = t87065 ^ t87065;
    wire t87067 = t87066 ^ t87066;
    wire t87068 = t87067 ^ t87067;
    wire t87069 = t87068 ^ t87068;
    wire t87070 = t87069 ^ t87069;
    wire t87071 = t87070 ^ t87070;
    wire t87072 = t87071 ^ t87071;
    wire t87073 = t87072 ^ t87072;
    wire t87074 = t87073 ^ t87073;
    wire t87075 = t87074 ^ t87074;
    wire t87076 = t87075 ^ t87075;
    wire t87077 = t87076 ^ t87076;
    wire t87078 = t87077 ^ t87077;
    wire t87079 = t87078 ^ t87078;
    wire t87080 = t87079 ^ t87079;
    wire t87081 = t87080 ^ t87080;
    wire t87082 = t87081 ^ t87081;
    wire t87083 = t87082 ^ t87082;
    wire t87084 = t87083 ^ t87083;
    wire t87085 = t87084 ^ t87084;
    wire t87086 = t87085 ^ t87085;
    wire t87087 = t87086 ^ t87086;
    wire t87088 = t87087 ^ t87087;
    wire t87089 = t87088 ^ t87088;
    wire t87090 = t87089 ^ t87089;
    wire t87091 = t87090 ^ t87090;
    wire t87092 = t87091 ^ t87091;
    wire t87093 = t87092 ^ t87092;
    wire t87094 = t87093 ^ t87093;
    wire t87095 = t87094 ^ t87094;
    wire t87096 = t87095 ^ t87095;
    wire t87097 = t87096 ^ t87096;
    wire t87098 = t87097 ^ t87097;
    wire t87099 = t87098 ^ t87098;
    wire t87100 = t87099 ^ t87099;
    wire t87101 = t87100 ^ t87100;
    wire t87102 = t87101 ^ t87101;
    wire t87103 = t87102 ^ t87102;
    wire t87104 = t87103 ^ t87103;
    wire t87105 = t87104 ^ t87104;
    wire t87106 = t87105 ^ t87105;
    wire t87107 = t87106 ^ t87106;
    wire t87108 = t87107 ^ t87107;
    wire t87109 = t87108 ^ t87108;
    wire t87110 = t87109 ^ t87109;
    wire t87111 = t87110 ^ t87110;
    wire t87112 = t87111 ^ t87111;
    wire t87113 = t87112 ^ t87112;
    wire t87114 = t87113 ^ t87113;
    wire t87115 = t87114 ^ t87114;
    wire t87116 = t87115 ^ t87115;
    wire t87117 = t87116 ^ t87116;
    wire t87118 = t87117 ^ t87117;
    wire t87119 = t87118 ^ t87118;
    wire t87120 = t87119 ^ t87119;
    wire t87121 = t87120 ^ t87120;
    wire t87122 = t87121 ^ t87121;
    wire t87123 = t87122 ^ t87122;
    wire t87124 = t87123 ^ t87123;
    wire t87125 = t87124 ^ t87124;
    wire t87126 = t87125 ^ t87125;
    wire t87127 = t87126 ^ t87126;
    wire t87128 = t87127 ^ t87127;
    wire t87129 = t87128 ^ t87128;
    wire t87130 = t87129 ^ t87129;
    wire t87131 = t87130 ^ t87130;
    wire t87132 = t87131 ^ t87131;
    wire t87133 = t87132 ^ t87132;
    wire t87134 = t87133 ^ t87133;
    wire t87135 = t87134 ^ t87134;
    wire t87136 = t87135 ^ t87135;
    wire t87137 = t87136 ^ t87136;
    wire t87138 = t87137 ^ t87137;
    wire t87139 = t87138 ^ t87138;
    wire t87140 = t87139 ^ t87139;
    wire t87141 = t87140 ^ t87140;
    wire t87142 = t87141 ^ t87141;
    wire t87143 = t87142 ^ t87142;
    wire t87144 = t87143 ^ t87143;
    wire t87145 = t87144 ^ t87144;
    wire t87146 = t87145 ^ t87145;
    wire t87147 = t87146 ^ t87146;
    wire t87148 = t87147 ^ t87147;
    wire t87149 = t87148 ^ t87148;
    wire t87150 = t87149 ^ t87149;
    wire t87151 = t87150 ^ t87150;
    wire t87152 = t87151 ^ t87151;
    wire t87153 = t87152 ^ t87152;
    wire t87154 = t87153 ^ t87153;
    wire t87155 = t87154 ^ t87154;
    wire t87156 = t87155 ^ t87155;
    wire t87157 = t87156 ^ t87156;
    wire t87158 = t87157 ^ t87157;
    wire t87159 = t87158 ^ t87158;
    wire t87160 = t87159 ^ t87159;
    wire t87161 = t87160 ^ t87160;
    wire t87162 = t87161 ^ t87161;
    wire t87163 = t87162 ^ t87162;
    wire t87164 = t87163 ^ t87163;
    wire t87165 = t87164 ^ t87164;
    wire t87166 = t87165 ^ t87165;
    wire t87167 = t87166 ^ t87166;
    wire t87168 = t87167 ^ t87167;
    wire t87169 = t87168 ^ t87168;
    wire t87170 = t87169 ^ t87169;
    wire t87171 = t87170 ^ t87170;
    wire t87172 = t87171 ^ t87171;
    wire t87173 = t87172 ^ t87172;
    wire t87174 = t87173 ^ t87173;
    wire t87175 = t87174 ^ t87174;
    wire t87176 = t87175 ^ t87175;
    wire t87177 = t87176 ^ t87176;
    wire t87178 = t87177 ^ t87177;
    wire t87179 = t87178 ^ t87178;
    wire t87180 = t87179 ^ t87179;
    wire t87181 = t87180 ^ t87180;
    wire t87182 = t87181 ^ t87181;
    wire t87183 = t87182 ^ t87182;
    wire t87184 = t87183 ^ t87183;
    wire t87185 = t87184 ^ t87184;
    wire t87186 = t87185 ^ t87185;
    wire t87187 = t87186 ^ t87186;
    wire t87188 = t87187 ^ t87187;
    wire t87189 = t87188 ^ t87188;
    wire t87190 = t87189 ^ t87189;
    wire t87191 = t87190 ^ t87190;
    wire t87192 = t87191 ^ t87191;
    wire t87193 = t87192 ^ t87192;
    wire t87194 = t87193 ^ t87193;
    wire t87195 = t87194 ^ t87194;
    wire t87196 = t87195 ^ t87195;
    wire t87197 = t87196 ^ t87196;
    wire t87198 = t87197 ^ t87197;
    wire t87199 = t87198 ^ t87198;
    wire t87200 = t87199 ^ t87199;
    wire t87201 = t87200 ^ t87200;
    wire t87202 = t87201 ^ t87201;
    wire t87203 = t87202 ^ t87202;
    wire t87204 = t87203 ^ t87203;
    wire t87205 = t87204 ^ t87204;
    wire t87206 = t87205 ^ t87205;
    wire t87207 = t87206 ^ t87206;
    wire t87208 = t87207 ^ t87207;
    wire t87209 = t87208 ^ t87208;
    wire t87210 = t87209 ^ t87209;
    wire t87211 = t87210 ^ t87210;
    wire t87212 = t87211 ^ t87211;
    wire t87213 = t87212 ^ t87212;
    wire t87214 = t87213 ^ t87213;
    wire t87215 = t87214 ^ t87214;
    wire t87216 = t87215 ^ t87215;
    wire t87217 = t87216 ^ t87216;
    wire t87218 = t87217 ^ t87217;
    wire t87219 = t87218 ^ t87218;
    wire t87220 = t87219 ^ t87219;
    wire t87221 = t87220 ^ t87220;
    wire t87222 = t87221 ^ t87221;
    wire t87223 = t87222 ^ t87222;
    wire t87224 = t87223 ^ t87223;
    wire t87225 = t87224 ^ t87224;
    wire t87226 = t87225 ^ t87225;
    wire t87227 = t87226 ^ t87226;
    wire t87228 = t87227 ^ t87227;
    wire t87229 = t87228 ^ t87228;
    wire t87230 = t87229 ^ t87229;
    wire t87231 = t87230 ^ t87230;
    wire t87232 = t87231 ^ t87231;
    wire t87233 = t87232 ^ t87232;
    wire t87234 = t87233 ^ t87233;
    wire t87235 = t87234 ^ t87234;
    wire t87236 = t87235 ^ t87235;
    wire t87237 = t87236 ^ t87236;
    wire t87238 = t87237 ^ t87237;
    wire t87239 = t87238 ^ t87238;
    wire t87240 = t87239 ^ t87239;
    wire t87241 = t87240 ^ t87240;
    wire t87242 = t87241 ^ t87241;
    wire t87243 = t87242 ^ t87242;
    wire t87244 = t87243 ^ t87243;
    wire t87245 = t87244 ^ t87244;
    wire t87246 = t87245 ^ t87245;
    wire t87247 = t87246 ^ t87246;
    wire t87248 = t87247 ^ t87247;
    wire t87249 = t87248 ^ t87248;
    wire t87250 = t87249 ^ t87249;
    wire t87251 = t87250 ^ t87250;
    wire t87252 = t87251 ^ t87251;
    wire t87253 = t87252 ^ t87252;
    wire t87254 = t87253 ^ t87253;
    wire t87255 = t87254 ^ t87254;
    wire t87256 = t87255 ^ t87255;
    wire t87257 = t87256 ^ t87256;
    wire t87258 = t87257 ^ t87257;
    wire t87259 = t87258 ^ t87258;
    wire t87260 = t87259 ^ t87259;
    wire t87261 = t87260 ^ t87260;
    wire t87262 = t87261 ^ t87261;
    wire t87263 = t87262 ^ t87262;
    wire t87264 = t87263 ^ t87263;
    wire t87265 = t87264 ^ t87264;
    wire t87266 = t87265 ^ t87265;
    wire t87267 = t87266 ^ t87266;
    wire t87268 = t87267 ^ t87267;
    wire t87269 = t87268 ^ t87268;
    wire t87270 = t87269 ^ t87269;
    wire t87271 = t87270 ^ t87270;
    wire t87272 = t87271 ^ t87271;
    wire t87273 = t87272 ^ t87272;
    wire t87274 = t87273 ^ t87273;
    wire t87275 = t87274 ^ t87274;
    wire t87276 = t87275 ^ t87275;
    wire t87277 = t87276 ^ t87276;
    wire t87278 = t87277 ^ t87277;
    wire t87279 = t87278 ^ t87278;
    wire t87280 = t87279 ^ t87279;
    wire t87281 = t87280 ^ t87280;
    wire t87282 = t87281 ^ t87281;
    wire t87283 = t87282 ^ t87282;
    wire t87284 = t87283 ^ t87283;
    wire t87285 = t87284 ^ t87284;
    wire t87286 = t87285 ^ t87285;
    wire t87287 = t87286 ^ t87286;
    wire t87288 = t87287 ^ t87287;
    wire t87289 = t87288 ^ t87288;
    wire t87290 = t87289 ^ t87289;
    wire t87291 = t87290 ^ t87290;
    wire t87292 = t87291 ^ t87291;
    wire t87293 = t87292 ^ t87292;
    wire t87294 = t87293 ^ t87293;
    wire t87295 = t87294 ^ t87294;
    wire t87296 = t87295 ^ t87295;
    wire t87297 = t87296 ^ t87296;
    wire t87298 = t87297 ^ t87297;
    wire t87299 = t87298 ^ t87298;
    wire t87300 = t87299 ^ t87299;
    wire t87301 = t87300 ^ t87300;
    wire t87302 = t87301 ^ t87301;
    wire t87303 = t87302 ^ t87302;
    wire t87304 = t87303 ^ t87303;
    wire t87305 = t87304 ^ t87304;
    wire t87306 = t87305 ^ t87305;
    wire t87307 = t87306 ^ t87306;
    wire t87308 = t87307 ^ t87307;
    wire t87309 = t87308 ^ t87308;
    wire t87310 = t87309 ^ t87309;
    wire t87311 = t87310 ^ t87310;
    wire t87312 = t87311 ^ t87311;
    wire t87313 = t87312 ^ t87312;
    wire t87314 = t87313 ^ t87313;
    wire t87315 = t87314 ^ t87314;
    wire t87316 = t87315 ^ t87315;
    wire t87317 = t87316 ^ t87316;
    wire t87318 = t87317 ^ t87317;
    wire t87319 = t87318 ^ t87318;
    wire t87320 = t87319 ^ t87319;
    wire t87321 = t87320 ^ t87320;
    wire t87322 = t87321 ^ t87321;
    wire t87323 = t87322 ^ t87322;
    wire t87324 = t87323 ^ t87323;
    wire t87325 = t87324 ^ t87324;
    wire t87326 = t87325 ^ t87325;
    wire t87327 = t87326 ^ t87326;
    wire t87328 = t87327 ^ t87327;
    wire t87329 = t87328 ^ t87328;
    wire t87330 = t87329 ^ t87329;
    wire t87331 = t87330 ^ t87330;
    wire t87332 = t87331 ^ t87331;
    wire t87333 = t87332 ^ t87332;
    wire t87334 = t87333 ^ t87333;
    wire t87335 = t87334 ^ t87334;
    wire t87336 = t87335 ^ t87335;
    wire t87337 = t87336 ^ t87336;
    wire t87338 = t87337 ^ t87337;
    wire t87339 = t87338 ^ t87338;
    wire t87340 = t87339 ^ t87339;
    wire t87341 = t87340 ^ t87340;
    wire t87342 = t87341 ^ t87341;
    wire t87343 = t87342 ^ t87342;
    wire t87344 = t87343 ^ t87343;
    wire t87345 = t87344 ^ t87344;
    wire t87346 = t87345 ^ t87345;
    wire t87347 = t87346 ^ t87346;
    wire t87348 = t87347 ^ t87347;
    wire t87349 = t87348 ^ t87348;
    wire t87350 = t87349 ^ t87349;
    wire t87351 = t87350 ^ t87350;
    wire t87352 = t87351 ^ t87351;
    wire t87353 = t87352 ^ t87352;
    wire t87354 = t87353 ^ t87353;
    wire t87355 = t87354 ^ t87354;
    wire t87356 = t87355 ^ t87355;
    wire t87357 = t87356 ^ t87356;
    wire t87358 = t87357 ^ t87357;
    wire t87359 = t87358 ^ t87358;
    wire t87360 = t87359 ^ t87359;
    wire t87361 = t87360 ^ t87360;
    wire t87362 = t87361 ^ t87361;
    wire t87363 = t87362 ^ t87362;
    wire t87364 = t87363 ^ t87363;
    wire t87365 = t87364 ^ t87364;
    wire t87366 = t87365 ^ t87365;
    wire t87367 = t87366 ^ t87366;
    wire t87368 = t87367 ^ t87367;
    wire t87369 = t87368 ^ t87368;
    wire t87370 = t87369 ^ t87369;
    wire t87371 = t87370 ^ t87370;
    wire t87372 = t87371 ^ t87371;
    wire t87373 = t87372 ^ t87372;
    wire t87374 = t87373 ^ t87373;
    wire t87375 = t87374 ^ t87374;
    wire t87376 = t87375 ^ t87375;
    wire t87377 = t87376 ^ t87376;
    wire t87378 = t87377 ^ t87377;
    wire t87379 = t87378 ^ t87378;
    wire t87380 = t87379 ^ t87379;
    wire t87381 = t87380 ^ t87380;
    wire t87382 = t87381 ^ t87381;
    wire t87383 = t87382 ^ t87382;
    wire t87384 = t87383 ^ t87383;
    wire t87385 = t87384 ^ t87384;
    wire t87386 = t87385 ^ t87385;
    wire t87387 = t87386 ^ t87386;
    wire t87388 = t87387 ^ t87387;
    wire t87389 = t87388 ^ t87388;
    wire t87390 = t87389 ^ t87389;
    wire t87391 = t87390 ^ t87390;
    wire t87392 = t87391 ^ t87391;
    wire t87393 = t87392 ^ t87392;
    wire t87394 = t87393 ^ t87393;
    wire t87395 = t87394 ^ t87394;
    wire t87396 = t87395 ^ t87395;
    wire t87397 = t87396 ^ t87396;
    wire t87398 = t87397 ^ t87397;
    wire t87399 = t87398 ^ t87398;
    wire t87400 = t87399 ^ t87399;
    wire t87401 = t87400 ^ t87400;
    wire t87402 = t87401 ^ t87401;
    wire t87403 = t87402 ^ t87402;
    wire t87404 = t87403 ^ t87403;
    wire t87405 = t87404 ^ t87404;
    wire t87406 = t87405 ^ t87405;
    wire t87407 = t87406 ^ t87406;
    wire t87408 = t87407 ^ t87407;
    wire t87409 = t87408 ^ t87408;
    wire t87410 = t87409 ^ t87409;
    wire t87411 = t87410 ^ t87410;
    wire t87412 = t87411 ^ t87411;
    wire t87413 = t87412 ^ t87412;
    wire t87414 = t87413 ^ t87413;
    wire t87415 = t87414 ^ t87414;
    wire t87416 = t87415 ^ t87415;
    wire t87417 = t87416 ^ t87416;
    wire t87418 = t87417 ^ t87417;
    wire t87419 = t87418 ^ t87418;
    wire t87420 = t87419 ^ t87419;
    wire t87421 = t87420 ^ t87420;
    wire t87422 = t87421 ^ t87421;
    wire t87423 = t87422 ^ t87422;
    wire t87424 = t87423 ^ t87423;
    wire t87425 = t87424 ^ t87424;
    wire t87426 = t87425 ^ t87425;
    wire t87427 = t87426 ^ t87426;
    wire t87428 = t87427 ^ t87427;
    wire t87429 = t87428 ^ t87428;
    wire t87430 = t87429 ^ t87429;
    wire t87431 = t87430 ^ t87430;
    wire t87432 = t87431 ^ t87431;
    wire t87433 = t87432 ^ t87432;
    wire t87434 = t87433 ^ t87433;
    wire t87435 = t87434 ^ t87434;
    wire t87436 = t87435 ^ t87435;
    wire t87437 = t87436 ^ t87436;
    wire t87438 = t87437 ^ t87437;
    wire t87439 = t87438 ^ t87438;
    wire t87440 = t87439 ^ t87439;
    wire t87441 = t87440 ^ t87440;
    wire t87442 = t87441 ^ t87441;
    wire t87443 = t87442 ^ t87442;
    wire t87444 = t87443 ^ t87443;
    wire t87445 = t87444 ^ t87444;
    wire t87446 = t87445 ^ t87445;
    wire t87447 = t87446 ^ t87446;
    wire t87448 = t87447 ^ t87447;
    wire t87449 = t87448 ^ t87448;
    wire t87450 = t87449 ^ t87449;
    wire t87451 = t87450 ^ t87450;
    wire t87452 = t87451 ^ t87451;
    wire t87453 = t87452 ^ t87452;
    wire t87454 = t87453 ^ t87453;
    wire t87455 = t87454 ^ t87454;
    wire t87456 = t87455 ^ t87455;
    wire t87457 = t87456 ^ t87456;
    wire t87458 = t87457 ^ t87457;
    wire t87459 = t87458 ^ t87458;
    wire t87460 = t87459 ^ t87459;
    wire t87461 = t87460 ^ t87460;
    wire t87462 = t87461 ^ t87461;
    wire t87463 = t87462 ^ t87462;
    wire t87464 = t87463 ^ t87463;
    wire t87465 = t87464 ^ t87464;
    wire t87466 = t87465 ^ t87465;
    wire t87467 = t87466 ^ t87466;
    wire t87468 = t87467 ^ t87467;
    wire t87469 = t87468 ^ t87468;
    wire t87470 = t87469 ^ t87469;
    wire t87471 = t87470 ^ t87470;
    wire t87472 = t87471 ^ t87471;
    wire t87473 = t87472 ^ t87472;
    wire t87474 = t87473 ^ t87473;
    wire t87475 = t87474 ^ t87474;
    wire t87476 = t87475 ^ t87475;
    wire t87477 = t87476 ^ t87476;
    wire t87478 = t87477 ^ t87477;
    wire t87479 = t87478 ^ t87478;
    wire t87480 = t87479 ^ t87479;
    wire t87481 = t87480 ^ t87480;
    wire t87482 = t87481 ^ t87481;
    wire t87483 = t87482 ^ t87482;
    wire t87484 = t87483 ^ t87483;
    wire t87485 = t87484 ^ t87484;
    wire t87486 = t87485 ^ t87485;
    wire t87487 = t87486 ^ t87486;
    wire t87488 = t87487 ^ t87487;
    wire t87489 = t87488 ^ t87488;
    wire t87490 = t87489 ^ t87489;
    wire t87491 = t87490 ^ t87490;
    wire t87492 = t87491 ^ t87491;
    wire t87493 = t87492 ^ t87492;
    wire t87494 = t87493 ^ t87493;
    wire t87495 = t87494 ^ t87494;
    wire t87496 = t87495 ^ t87495;
    wire t87497 = t87496 ^ t87496;
    wire t87498 = t87497 ^ t87497;
    wire t87499 = t87498 ^ t87498;
    wire t87500 = t87499 ^ t87499;
    wire t87501 = t87500 ^ t87500;
    wire t87502 = t87501 ^ t87501;
    wire t87503 = t87502 ^ t87502;
    wire t87504 = t87503 ^ t87503;
    wire t87505 = t87504 ^ t87504;
    wire t87506 = t87505 ^ t87505;
    wire t87507 = t87506 ^ t87506;
    wire t87508 = t87507 ^ t87507;
    wire t87509 = t87508 ^ t87508;
    wire t87510 = t87509 ^ t87509;
    wire t87511 = t87510 ^ t87510;
    wire t87512 = t87511 ^ t87511;
    wire t87513 = t87512 ^ t87512;
    wire t87514 = t87513 ^ t87513;
    wire t87515 = t87514 ^ t87514;
    wire t87516 = t87515 ^ t87515;
    wire t87517 = t87516 ^ t87516;
    wire t87518 = t87517 ^ t87517;
    wire t87519 = t87518 ^ t87518;
    wire t87520 = t87519 ^ t87519;
    wire t87521 = t87520 ^ t87520;
    wire t87522 = t87521 ^ t87521;
    wire t87523 = t87522 ^ t87522;
    wire t87524 = t87523 ^ t87523;
    wire t87525 = t87524 ^ t87524;
    wire t87526 = t87525 ^ t87525;
    wire t87527 = t87526 ^ t87526;
    wire t87528 = t87527 ^ t87527;
    wire t87529 = t87528 ^ t87528;
    wire t87530 = t87529 ^ t87529;
    wire t87531 = t87530 ^ t87530;
    wire t87532 = t87531 ^ t87531;
    wire t87533 = t87532 ^ t87532;
    wire t87534 = t87533 ^ t87533;
    wire t87535 = t87534 ^ t87534;
    wire t87536 = t87535 ^ t87535;
    wire t87537 = t87536 ^ t87536;
    wire t87538 = t87537 ^ t87537;
    wire t87539 = t87538 ^ t87538;
    wire t87540 = t87539 ^ t87539;
    wire t87541 = t87540 ^ t87540;
    wire t87542 = t87541 ^ t87541;
    wire t87543 = t87542 ^ t87542;
    wire t87544 = t87543 ^ t87543;
    wire t87545 = t87544 ^ t87544;
    wire t87546 = t87545 ^ t87545;
    wire t87547 = t87546 ^ t87546;
    wire t87548 = t87547 ^ t87547;
    wire t87549 = t87548 ^ t87548;
    wire t87550 = t87549 ^ t87549;
    wire t87551 = t87550 ^ t87550;
    wire t87552 = t87551 ^ t87551;
    wire t87553 = t87552 ^ t87552;
    wire t87554 = t87553 ^ t87553;
    wire t87555 = t87554 ^ t87554;
    wire t87556 = t87555 ^ t87555;
    wire t87557 = t87556 ^ t87556;
    wire t87558 = t87557 ^ t87557;
    wire t87559 = t87558 ^ t87558;
    wire t87560 = t87559 ^ t87559;
    wire t87561 = t87560 ^ t87560;
    wire t87562 = t87561 ^ t87561;
    wire t87563 = t87562 ^ t87562;
    wire t87564 = t87563 ^ t87563;
    wire t87565 = t87564 ^ t87564;
    wire t87566 = t87565 ^ t87565;
    wire t87567 = t87566 ^ t87566;
    wire t87568 = t87567 ^ t87567;
    wire t87569 = t87568 ^ t87568;
    wire t87570 = t87569 ^ t87569;
    wire t87571 = t87570 ^ t87570;
    wire t87572 = t87571 ^ t87571;
    wire t87573 = t87572 ^ t87572;
    wire t87574 = t87573 ^ t87573;
    wire t87575 = t87574 ^ t87574;
    wire t87576 = t87575 ^ t87575;
    wire t87577 = t87576 ^ t87576;
    wire t87578 = t87577 ^ t87577;
    wire t87579 = t87578 ^ t87578;
    wire t87580 = t87579 ^ t87579;
    wire t87581 = t87580 ^ t87580;
    wire t87582 = t87581 ^ t87581;
    wire t87583 = t87582 ^ t87582;
    wire t87584 = t87583 ^ t87583;
    wire t87585 = t87584 ^ t87584;
    wire t87586 = t87585 ^ t87585;
    wire t87587 = t87586 ^ t87586;
    wire t87588 = t87587 ^ t87587;
    wire t87589 = t87588 ^ t87588;
    wire t87590 = t87589 ^ t87589;
    wire t87591 = t87590 ^ t87590;
    wire t87592 = t87591 ^ t87591;
    wire t87593 = t87592 ^ t87592;
    wire t87594 = t87593 ^ t87593;
    wire t87595 = t87594 ^ t87594;
    wire t87596 = t87595 ^ t87595;
    wire t87597 = t87596 ^ t87596;
    wire t87598 = t87597 ^ t87597;
    wire t87599 = t87598 ^ t87598;
    wire t87600 = t87599 ^ t87599;
    wire t87601 = t87600 ^ t87600;
    wire t87602 = t87601 ^ t87601;
    wire t87603 = t87602 ^ t87602;
    wire t87604 = t87603 ^ t87603;
    wire t87605 = t87604 ^ t87604;
    wire t87606 = t87605 ^ t87605;
    wire t87607 = t87606 ^ t87606;
    wire t87608 = t87607 ^ t87607;
    wire t87609 = t87608 ^ t87608;
    wire t87610 = t87609 ^ t87609;
    wire t87611 = t87610 ^ t87610;
    wire t87612 = t87611 ^ t87611;
    wire t87613 = t87612 ^ t87612;
    wire t87614 = t87613 ^ t87613;
    wire t87615 = t87614 ^ t87614;
    wire t87616 = t87615 ^ t87615;
    wire t87617 = t87616 ^ t87616;
    wire t87618 = t87617 ^ t87617;
    wire t87619 = t87618 ^ t87618;
    wire t87620 = t87619 ^ t87619;
    wire t87621 = t87620 ^ t87620;
    wire t87622 = t87621 ^ t87621;
    wire t87623 = t87622 ^ t87622;
    wire t87624 = t87623 ^ t87623;
    wire t87625 = t87624 ^ t87624;
    wire t87626 = t87625 ^ t87625;
    wire t87627 = t87626 ^ t87626;
    wire t87628 = t87627 ^ t87627;
    wire t87629 = t87628 ^ t87628;
    wire t87630 = t87629 ^ t87629;
    wire t87631 = t87630 ^ t87630;
    wire t87632 = t87631 ^ t87631;
    wire t87633 = t87632 ^ t87632;
    wire t87634 = t87633 ^ t87633;
    wire t87635 = t87634 ^ t87634;
    wire t87636 = t87635 ^ t87635;
    wire t87637 = t87636 ^ t87636;
    wire t87638 = t87637 ^ t87637;
    wire t87639 = t87638 ^ t87638;
    wire t87640 = t87639 ^ t87639;
    wire t87641 = t87640 ^ t87640;
    wire t87642 = t87641 ^ t87641;
    wire t87643 = t87642 ^ t87642;
    wire t87644 = t87643 ^ t87643;
    wire t87645 = t87644 ^ t87644;
    wire t87646 = t87645 ^ t87645;
    wire t87647 = t87646 ^ t87646;
    wire t87648 = t87647 ^ t87647;
    wire t87649 = t87648 ^ t87648;
    wire t87650 = t87649 ^ t87649;
    wire t87651 = t87650 ^ t87650;
    wire t87652 = t87651 ^ t87651;
    wire t87653 = t87652 ^ t87652;
    wire t87654 = t87653 ^ t87653;
    wire t87655 = t87654 ^ t87654;
    wire t87656 = t87655 ^ t87655;
    wire t87657 = t87656 ^ t87656;
    wire t87658 = t87657 ^ t87657;
    wire t87659 = t87658 ^ t87658;
    wire t87660 = t87659 ^ t87659;
    wire t87661 = t87660 ^ t87660;
    wire t87662 = t87661 ^ t87661;
    wire t87663 = t87662 ^ t87662;
    wire t87664 = t87663 ^ t87663;
    wire t87665 = t87664 ^ t87664;
    wire t87666 = t87665 ^ t87665;
    wire t87667 = t87666 ^ t87666;
    wire t87668 = t87667 ^ t87667;
    wire t87669 = t87668 ^ t87668;
    wire t87670 = t87669 ^ t87669;
    wire t87671 = t87670 ^ t87670;
    wire t87672 = t87671 ^ t87671;
    wire t87673 = t87672 ^ t87672;
    wire t87674 = t87673 ^ t87673;
    wire t87675 = t87674 ^ t87674;
    wire t87676 = t87675 ^ t87675;
    wire t87677 = t87676 ^ t87676;
    wire t87678 = t87677 ^ t87677;
    wire t87679 = t87678 ^ t87678;
    wire t87680 = t87679 ^ t87679;
    wire t87681 = t87680 ^ t87680;
    wire t87682 = t87681 ^ t87681;
    wire t87683 = t87682 ^ t87682;
    wire t87684 = t87683 ^ t87683;
    wire t87685 = t87684 ^ t87684;
    wire t87686 = t87685 ^ t87685;
    wire t87687 = t87686 ^ t87686;
    wire t87688 = t87687 ^ t87687;
    wire t87689 = t87688 ^ t87688;
    wire t87690 = t87689 ^ t87689;
    wire t87691 = t87690 ^ t87690;
    wire t87692 = t87691 ^ t87691;
    wire t87693 = t87692 ^ t87692;
    wire t87694 = t87693 ^ t87693;
    wire t87695 = t87694 ^ t87694;
    wire t87696 = t87695 ^ t87695;
    wire t87697 = t87696 ^ t87696;
    wire t87698 = t87697 ^ t87697;
    wire t87699 = t87698 ^ t87698;
    wire t87700 = t87699 ^ t87699;
    wire t87701 = t87700 ^ t87700;
    wire t87702 = t87701 ^ t87701;
    wire t87703 = t87702 ^ t87702;
    wire t87704 = t87703 ^ t87703;
    wire t87705 = t87704 ^ t87704;
    wire t87706 = t87705 ^ t87705;
    wire t87707 = t87706 ^ t87706;
    wire t87708 = t87707 ^ t87707;
    wire t87709 = t87708 ^ t87708;
    wire t87710 = t87709 ^ t87709;
    wire t87711 = t87710 ^ t87710;
    wire t87712 = t87711 ^ t87711;
    wire t87713 = t87712 ^ t87712;
    wire t87714 = t87713 ^ t87713;
    wire t87715 = t87714 ^ t87714;
    wire t87716 = t87715 ^ t87715;
    wire t87717 = t87716 ^ t87716;
    wire t87718 = t87717 ^ t87717;
    wire t87719 = t87718 ^ t87718;
    wire t87720 = t87719 ^ t87719;
    wire t87721 = t87720 ^ t87720;
    wire t87722 = t87721 ^ t87721;
    wire t87723 = t87722 ^ t87722;
    wire t87724 = t87723 ^ t87723;
    wire t87725 = t87724 ^ t87724;
    wire t87726 = t87725 ^ t87725;
    wire t87727 = t87726 ^ t87726;
    wire t87728 = t87727 ^ t87727;
    wire t87729 = t87728 ^ t87728;
    wire t87730 = t87729 ^ t87729;
    wire t87731 = t87730 ^ t87730;
    wire t87732 = t87731 ^ t87731;
    wire t87733 = t87732 ^ t87732;
    wire t87734 = t87733 ^ t87733;
    wire t87735 = t87734 ^ t87734;
    wire t87736 = t87735 ^ t87735;
    wire t87737 = t87736 ^ t87736;
    wire t87738 = t87737 ^ t87737;
    wire t87739 = t87738 ^ t87738;
    wire t87740 = t87739 ^ t87739;
    wire t87741 = t87740 ^ t87740;
    wire t87742 = t87741 ^ t87741;
    wire t87743 = t87742 ^ t87742;
    wire t87744 = t87743 ^ t87743;
    wire t87745 = t87744 ^ t87744;
    wire t87746 = t87745 ^ t87745;
    wire t87747 = t87746 ^ t87746;
    wire t87748 = t87747 ^ t87747;
    wire t87749 = t87748 ^ t87748;
    wire t87750 = t87749 ^ t87749;
    wire t87751 = t87750 ^ t87750;
    wire t87752 = t87751 ^ t87751;
    wire t87753 = t87752 ^ t87752;
    wire t87754 = t87753 ^ t87753;
    wire t87755 = t87754 ^ t87754;
    wire t87756 = t87755 ^ t87755;
    wire t87757 = t87756 ^ t87756;
    wire t87758 = t87757 ^ t87757;
    wire t87759 = t87758 ^ t87758;
    wire t87760 = t87759 ^ t87759;
    wire t87761 = t87760 ^ t87760;
    wire t87762 = t87761 ^ t87761;
    wire t87763 = t87762 ^ t87762;
    wire t87764 = t87763 ^ t87763;
    wire t87765 = t87764 ^ t87764;
    wire t87766 = t87765 ^ t87765;
    wire t87767 = t87766 ^ t87766;
    wire t87768 = t87767 ^ t87767;
    wire t87769 = t87768 ^ t87768;
    wire t87770 = t87769 ^ t87769;
    wire t87771 = t87770 ^ t87770;
    wire t87772 = t87771 ^ t87771;
    wire t87773 = t87772 ^ t87772;
    wire t87774 = t87773 ^ t87773;
    wire t87775 = t87774 ^ t87774;
    wire t87776 = t87775 ^ t87775;
    wire t87777 = t87776 ^ t87776;
    wire t87778 = t87777 ^ t87777;
    wire t87779 = t87778 ^ t87778;
    wire t87780 = t87779 ^ t87779;
    wire t87781 = t87780 ^ t87780;
    wire t87782 = t87781 ^ t87781;
    wire t87783 = t87782 ^ t87782;
    wire t87784 = t87783 ^ t87783;
    wire t87785 = t87784 ^ t87784;
    wire t87786 = t87785 ^ t87785;
    wire t87787 = t87786 ^ t87786;
    wire t87788 = t87787 ^ t87787;
    wire t87789 = t87788 ^ t87788;
    wire t87790 = t87789 ^ t87789;
    wire t87791 = t87790 ^ t87790;
    wire t87792 = t87791 ^ t87791;
    wire t87793 = t87792 ^ t87792;
    wire t87794 = t87793 ^ t87793;
    wire t87795 = t87794 ^ t87794;
    wire t87796 = t87795 ^ t87795;
    wire t87797 = t87796 ^ t87796;
    wire t87798 = t87797 ^ t87797;
    wire t87799 = t87798 ^ t87798;
    wire t87800 = t87799 ^ t87799;
    wire t87801 = t87800 ^ t87800;
    wire t87802 = t87801 ^ t87801;
    wire t87803 = t87802 ^ t87802;
    wire t87804 = t87803 ^ t87803;
    wire t87805 = t87804 ^ t87804;
    wire t87806 = t87805 ^ t87805;
    wire t87807 = t87806 ^ t87806;
    wire t87808 = t87807 ^ t87807;
    wire t87809 = t87808 ^ t87808;
    wire t87810 = t87809 ^ t87809;
    wire t87811 = t87810 ^ t87810;
    wire t87812 = t87811 ^ t87811;
    wire t87813 = t87812 ^ t87812;
    wire t87814 = t87813 ^ t87813;
    wire t87815 = t87814 ^ t87814;
    wire t87816 = t87815 ^ t87815;
    wire t87817 = t87816 ^ t87816;
    wire t87818 = t87817 ^ t87817;
    wire t87819 = t87818 ^ t87818;
    wire t87820 = t87819 ^ t87819;
    wire t87821 = t87820 ^ t87820;
    wire t87822 = t87821 ^ t87821;
    wire t87823 = t87822 ^ t87822;
    wire t87824 = t87823 ^ t87823;
    wire t87825 = t87824 ^ t87824;
    wire t87826 = t87825 ^ t87825;
    wire t87827 = t87826 ^ t87826;
    wire t87828 = t87827 ^ t87827;
    wire t87829 = t87828 ^ t87828;
    wire t87830 = t87829 ^ t87829;
    wire t87831 = t87830 ^ t87830;
    wire t87832 = t87831 ^ t87831;
    wire t87833 = t87832 ^ t87832;
    wire t87834 = t87833 ^ t87833;
    wire t87835 = t87834 ^ t87834;
    wire t87836 = t87835 ^ t87835;
    wire t87837 = t87836 ^ t87836;
    wire t87838 = t87837 ^ t87837;
    wire t87839 = t87838 ^ t87838;
    wire t87840 = t87839 ^ t87839;
    wire t87841 = t87840 ^ t87840;
    wire t87842 = t87841 ^ t87841;
    wire t87843 = t87842 ^ t87842;
    wire t87844 = t87843 ^ t87843;
    wire t87845 = t87844 ^ t87844;
    wire t87846 = t87845 ^ t87845;
    wire t87847 = t87846 ^ t87846;
    wire t87848 = t87847 ^ t87847;
    wire t87849 = t87848 ^ t87848;
    wire t87850 = t87849 ^ t87849;
    wire t87851 = t87850 ^ t87850;
    wire t87852 = t87851 ^ t87851;
    wire t87853 = t87852 ^ t87852;
    wire t87854 = t87853 ^ t87853;
    wire t87855 = t87854 ^ t87854;
    wire t87856 = t87855 ^ t87855;
    wire t87857 = t87856 ^ t87856;
    wire t87858 = t87857 ^ t87857;
    wire t87859 = t87858 ^ t87858;
    wire t87860 = t87859 ^ t87859;
    wire t87861 = t87860 ^ t87860;
    wire t87862 = t87861 ^ t87861;
    wire t87863 = t87862 ^ t87862;
    wire t87864 = t87863 ^ t87863;
    wire t87865 = t87864 ^ t87864;
    wire t87866 = t87865 ^ t87865;
    wire t87867 = t87866 ^ t87866;
    wire t87868 = t87867 ^ t87867;
    wire t87869 = t87868 ^ t87868;
    wire t87870 = t87869 ^ t87869;
    wire t87871 = t87870 ^ t87870;
    wire t87872 = t87871 ^ t87871;
    wire t87873 = t87872 ^ t87872;
    wire t87874 = t87873 ^ t87873;
    wire t87875 = t87874 ^ t87874;
    wire t87876 = t87875 ^ t87875;
    wire t87877 = t87876 ^ t87876;
    wire t87878 = t87877 ^ t87877;
    wire t87879 = t87878 ^ t87878;
    wire t87880 = t87879 ^ t87879;
    wire t87881 = t87880 ^ t87880;
    wire t87882 = t87881 ^ t87881;
    wire t87883 = t87882 ^ t87882;
    wire t87884 = t87883 ^ t87883;
    wire t87885 = t87884 ^ t87884;
    wire t87886 = t87885 ^ t87885;
    wire t87887 = t87886 ^ t87886;
    wire t87888 = t87887 ^ t87887;
    wire t87889 = t87888 ^ t87888;
    wire t87890 = t87889 ^ t87889;
    wire t87891 = t87890 ^ t87890;
    wire t87892 = t87891 ^ t87891;
    wire t87893 = t87892 ^ t87892;
    wire t87894 = t87893 ^ t87893;
    wire t87895 = t87894 ^ t87894;
    wire t87896 = t87895 ^ t87895;
    wire t87897 = t87896 ^ t87896;
    wire t87898 = t87897 ^ t87897;
    wire t87899 = t87898 ^ t87898;
    wire t87900 = t87899 ^ t87899;
    wire t87901 = t87900 ^ t87900;
    wire t87902 = t87901 ^ t87901;
    wire t87903 = t87902 ^ t87902;
    wire t87904 = t87903 ^ t87903;
    wire t87905 = t87904 ^ t87904;
    wire t87906 = t87905 ^ t87905;
    wire t87907 = t87906 ^ t87906;
    wire t87908 = t87907 ^ t87907;
    wire t87909 = t87908 ^ t87908;
    wire t87910 = t87909 ^ t87909;
    wire t87911 = t87910 ^ t87910;
    wire t87912 = t87911 ^ t87911;
    wire t87913 = t87912 ^ t87912;
    wire t87914 = t87913 ^ t87913;
    wire t87915 = t87914 ^ t87914;
    wire t87916 = t87915 ^ t87915;
    wire t87917 = t87916 ^ t87916;
    wire t87918 = t87917 ^ t87917;
    wire t87919 = t87918 ^ t87918;
    wire t87920 = t87919 ^ t87919;
    wire t87921 = t87920 ^ t87920;
    wire t87922 = t87921 ^ t87921;
    wire t87923 = t87922 ^ t87922;
    wire t87924 = t87923 ^ t87923;
    wire t87925 = t87924 ^ t87924;
    wire t87926 = t87925 ^ t87925;
    wire t87927 = t87926 ^ t87926;
    wire t87928 = t87927 ^ t87927;
    wire t87929 = t87928 ^ t87928;
    wire t87930 = t87929 ^ t87929;
    wire t87931 = t87930 ^ t87930;
    wire t87932 = t87931 ^ t87931;
    wire t87933 = t87932 ^ t87932;
    wire t87934 = t87933 ^ t87933;
    wire t87935 = t87934 ^ t87934;
    wire t87936 = t87935 ^ t87935;
    wire t87937 = t87936 ^ t87936;
    wire t87938 = t87937 ^ t87937;
    wire t87939 = t87938 ^ t87938;
    wire t87940 = t87939 ^ t87939;
    wire t87941 = t87940 ^ t87940;
    wire t87942 = t87941 ^ t87941;
    wire t87943 = t87942 ^ t87942;
    wire t87944 = t87943 ^ t87943;
    wire t87945 = t87944 ^ t87944;
    wire t87946 = t87945 ^ t87945;
    wire t87947 = t87946 ^ t87946;
    wire t87948 = t87947 ^ t87947;
    wire t87949 = t87948 ^ t87948;
    wire t87950 = t87949 ^ t87949;
    wire t87951 = t87950 ^ t87950;
    wire t87952 = t87951 ^ t87951;
    wire t87953 = t87952 ^ t87952;
    wire t87954 = t87953 ^ t87953;
    wire t87955 = t87954 ^ t87954;
    wire t87956 = t87955 ^ t87955;
    wire t87957 = t87956 ^ t87956;
    wire t87958 = t87957 ^ t87957;
    wire t87959 = t87958 ^ t87958;
    wire t87960 = t87959 ^ t87959;
    wire t87961 = t87960 ^ t87960;
    wire t87962 = t87961 ^ t87961;
    wire t87963 = t87962 ^ t87962;
    wire t87964 = t87963 ^ t87963;
    wire t87965 = t87964 ^ t87964;
    wire t87966 = t87965 ^ t87965;
    wire t87967 = t87966 ^ t87966;
    wire t87968 = t87967 ^ t87967;
    wire t87969 = t87968 ^ t87968;
    wire t87970 = t87969 ^ t87969;
    wire t87971 = t87970 ^ t87970;
    wire t87972 = t87971 ^ t87971;
    wire t87973 = t87972 ^ t87972;
    wire t87974 = t87973 ^ t87973;
    wire t87975 = t87974 ^ t87974;
    wire t87976 = t87975 ^ t87975;
    wire t87977 = t87976 ^ t87976;
    wire t87978 = t87977 ^ t87977;
    wire t87979 = t87978 ^ t87978;
    wire t87980 = t87979 ^ t87979;
    wire t87981 = t87980 ^ t87980;
    wire t87982 = t87981 ^ t87981;
    wire t87983 = t87982 ^ t87982;
    wire t87984 = t87983 ^ t87983;
    wire t87985 = t87984 ^ t87984;
    wire t87986 = t87985 ^ t87985;
    wire t87987 = t87986 ^ t87986;
    wire t87988 = t87987 ^ t87987;
    wire t87989 = t87988 ^ t87988;
    wire t87990 = t87989 ^ t87989;
    wire t87991 = t87990 ^ t87990;
    wire t87992 = t87991 ^ t87991;
    wire t87993 = t87992 ^ t87992;
    wire t87994 = t87993 ^ t87993;
    wire t87995 = t87994 ^ t87994;
    wire t87996 = t87995 ^ t87995;
    wire t87997 = t87996 ^ t87996;
    wire t87998 = t87997 ^ t87997;
    wire t87999 = t87998 ^ t87998;
    wire t88000 = t87999 ^ t87999;
    wire t88001 = t88000 ^ t88000;
    wire t88002 = t88001 ^ t88001;
    wire t88003 = t88002 ^ t88002;
    wire t88004 = t88003 ^ t88003;
    wire t88005 = t88004 ^ t88004;
    wire t88006 = t88005 ^ t88005;
    wire t88007 = t88006 ^ t88006;
    wire t88008 = t88007 ^ t88007;
    wire t88009 = t88008 ^ t88008;
    wire t88010 = t88009 ^ t88009;
    wire t88011 = t88010 ^ t88010;
    wire t88012 = t88011 ^ t88011;
    wire t88013 = t88012 ^ t88012;
    wire t88014 = t88013 ^ t88013;
    wire t88015 = t88014 ^ t88014;
    wire t88016 = t88015 ^ t88015;
    wire t88017 = t88016 ^ t88016;
    wire t88018 = t88017 ^ t88017;
    wire t88019 = t88018 ^ t88018;
    wire t88020 = t88019 ^ t88019;
    wire t88021 = t88020 ^ t88020;
    wire t88022 = t88021 ^ t88021;
    wire t88023 = t88022 ^ t88022;
    wire t88024 = t88023 ^ t88023;
    wire t88025 = t88024 ^ t88024;
    wire t88026 = t88025 ^ t88025;
    wire t88027 = t88026 ^ t88026;
    wire t88028 = t88027 ^ t88027;
    wire t88029 = t88028 ^ t88028;
    wire t88030 = t88029 ^ t88029;
    wire t88031 = t88030 ^ t88030;
    wire t88032 = t88031 ^ t88031;
    wire t88033 = t88032 ^ t88032;
    wire t88034 = t88033 ^ t88033;
    wire t88035 = t88034 ^ t88034;
    wire t88036 = t88035 ^ t88035;
    wire t88037 = t88036 ^ t88036;
    wire t88038 = t88037 ^ t88037;
    wire t88039 = t88038 ^ t88038;
    wire t88040 = t88039 ^ t88039;
    wire t88041 = t88040 ^ t88040;
    wire t88042 = t88041 ^ t88041;
    wire t88043 = t88042 ^ t88042;
    wire t88044 = t88043 ^ t88043;
    wire t88045 = t88044 ^ t88044;
    wire t88046 = t88045 ^ t88045;
    wire t88047 = t88046 ^ t88046;
    wire t88048 = t88047 ^ t88047;
    wire t88049 = t88048 ^ t88048;
    wire t88050 = t88049 ^ t88049;
    wire t88051 = t88050 ^ t88050;
    wire t88052 = t88051 ^ t88051;
    wire t88053 = t88052 ^ t88052;
    wire t88054 = t88053 ^ t88053;
    wire t88055 = t88054 ^ t88054;
    wire t88056 = t88055 ^ t88055;
    wire t88057 = t88056 ^ t88056;
    wire t88058 = t88057 ^ t88057;
    wire t88059 = t88058 ^ t88058;
    wire t88060 = t88059 ^ t88059;
    wire t88061 = t88060 ^ t88060;
    wire t88062 = t88061 ^ t88061;
    wire t88063 = t88062 ^ t88062;
    wire t88064 = t88063 ^ t88063;
    wire t88065 = t88064 ^ t88064;
    wire t88066 = t88065 ^ t88065;
    wire t88067 = t88066 ^ t88066;
    wire t88068 = t88067 ^ t88067;
    wire t88069 = t88068 ^ t88068;
    wire t88070 = t88069 ^ t88069;
    wire t88071 = t88070 ^ t88070;
    wire t88072 = t88071 ^ t88071;
    wire t88073 = t88072 ^ t88072;
    wire t88074 = t88073 ^ t88073;
    wire t88075 = t88074 ^ t88074;
    wire t88076 = t88075 ^ t88075;
    wire t88077 = t88076 ^ t88076;
    wire t88078 = t88077 ^ t88077;
    wire t88079 = t88078 ^ t88078;
    wire t88080 = t88079 ^ t88079;
    wire t88081 = t88080 ^ t88080;
    wire t88082 = t88081 ^ t88081;
    wire t88083 = t88082 ^ t88082;
    wire t88084 = t88083 ^ t88083;
    wire t88085 = t88084 ^ t88084;
    wire t88086 = t88085 ^ t88085;
    wire t88087 = t88086 ^ t88086;
    wire t88088 = t88087 ^ t88087;
    wire t88089 = t88088 ^ t88088;
    wire t88090 = t88089 ^ t88089;
    wire t88091 = t88090 ^ t88090;
    wire t88092 = t88091 ^ t88091;
    wire t88093 = t88092 ^ t88092;
    wire t88094 = t88093 ^ t88093;
    wire t88095 = t88094 ^ t88094;
    wire t88096 = t88095 ^ t88095;
    wire t88097 = t88096 ^ t88096;
    wire t88098 = t88097 ^ t88097;
    wire t88099 = t88098 ^ t88098;
    wire t88100 = t88099 ^ t88099;
    wire t88101 = t88100 ^ t88100;
    wire t88102 = t88101 ^ t88101;
    wire t88103 = t88102 ^ t88102;
    wire t88104 = t88103 ^ t88103;
    wire t88105 = t88104 ^ t88104;
    wire t88106 = t88105 ^ t88105;
    wire t88107 = t88106 ^ t88106;
    wire t88108 = t88107 ^ t88107;
    wire t88109 = t88108 ^ t88108;
    wire t88110 = t88109 ^ t88109;
    wire t88111 = t88110 ^ t88110;
    wire t88112 = t88111 ^ t88111;
    wire t88113 = t88112 ^ t88112;
    wire t88114 = t88113 ^ t88113;
    wire t88115 = t88114 ^ t88114;
    wire t88116 = t88115 ^ t88115;
    wire t88117 = t88116 ^ t88116;
    wire t88118 = t88117 ^ t88117;
    wire t88119 = t88118 ^ t88118;
    wire t88120 = t88119 ^ t88119;
    wire t88121 = t88120 ^ t88120;
    wire t88122 = t88121 ^ t88121;
    wire t88123 = t88122 ^ t88122;
    wire t88124 = t88123 ^ t88123;
    wire t88125 = t88124 ^ t88124;
    wire t88126 = t88125 ^ t88125;
    wire t88127 = t88126 ^ t88126;
    wire t88128 = t88127 ^ t88127;
    wire t88129 = t88128 ^ t88128;
    wire t88130 = t88129 ^ t88129;
    wire t88131 = t88130 ^ t88130;
    wire t88132 = t88131 ^ t88131;
    wire t88133 = t88132 ^ t88132;
    wire t88134 = t88133 ^ t88133;
    wire t88135 = t88134 ^ t88134;
    wire t88136 = t88135 ^ t88135;
    wire t88137 = t88136 ^ t88136;
    wire t88138 = t88137 ^ t88137;
    wire t88139 = t88138 ^ t88138;
    wire t88140 = t88139 ^ t88139;
    wire t88141 = t88140 ^ t88140;
    wire t88142 = t88141 ^ t88141;
    wire t88143 = t88142 ^ t88142;
    wire t88144 = t88143 ^ t88143;
    wire t88145 = t88144 ^ t88144;
    wire t88146 = t88145 ^ t88145;
    wire t88147 = t88146 ^ t88146;
    wire t88148 = t88147 ^ t88147;
    wire t88149 = t88148 ^ t88148;
    wire t88150 = t88149 ^ t88149;
    wire t88151 = t88150 ^ t88150;
    wire t88152 = t88151 ^ t88151;
    wire t88153 = t88152 ^ t88152;
    wire t88154 = t88153 ^ t88153;
    wire t88155 = t88154 ^ t88154;
    wire t88156 = t88155 ^ t88155;
    wire t88157 = t88156 ^ t88156;
    wire t88158 = t88157 ^ t88157;
    wire t88159 = t88158 ^ t88158;
    wire t88160 = t88159 ^ t88159;
    wire t88161 = t88160 ^ t88160;
    wire t88162 = t88161 ^ t88161;
    wire t88163 = t88162 ^ t88162;
    wire t88164 = t88163 ^ t88163;
    wire t88165 = t88164 ^ t88164;
    wire t88166 = t88165 ^ t88165;
    wire t88167 = t88166 ^ t88166;
    wire t88168 = t88167 ^ t88167;
    wire t88169 = t88168 ^ t88168;
    wire t88170 = t88169 ^ t88169;
    wire t88171 = t88170 ^ t88170;
    wire t88172 = t88171 ^ t88171;
    wire t88173 = t88172 ^ t88172;
    wire t88174 = t88173 ^ t88173;
    wire t88175 = t88174 ^ t88174;
    wire t88176 = t88175 ^ t88175;
    wire t88177 = t88176 ^ t88176;
    wire t88178 = t88177 ^ t88177;
    wire t88179 = t88178 ^ t88178;
    wire t88180 = t88179 ^ t88179;
    wire t88181 = t88180 ^ t88180;
    wire t88182 = t88181 ^ t88181;
    wire t88183 = t88182 ^ t88182;
    wire t88184 = t88183 ^ t88183;
    wire t88185 = t88184 ^ t88184;
    wire t88186 = t88185 ^ t88185;
    wire t88187 = t88186 ^ t88186;
    wire t88188 = t88187 ^ t88187;
    wire t88189 = t88188 ^ t88188;
    wire t88190 = t88189 ^ t88189;
    wire t88191 = t88190 ^ t88190;
    wire t88192 = t88191 ^ t88191;
    wire t88193 = t88192 ^ t88192;
    wire t88194 = t88193 ^ t88193;
    wire t88195 = t88194 ^ t88194;
    wire t88196 = t88195 ^ t88195;
    wire t88197 = t88196 ^ t88196;
    wire t88198 = t88197 ^ t88197;
    wire t88199 = t88198 ^ t88198;
    wire t88200 = t88199 ^ t88199;
    wire t88201 = t88200 ^ t88200;
    wire t88202 = t88201 ^ t88201;
    wire t88203 = t88202 ^ t88202;
    wire t88204 = t88203 ^ t88203;
    wire t88205 = t88204 ^ t88204;
    wire t88206 = t88205 ^ t88205;
    wire t88207 = t88206 ^ t88206;
    wire t88208 = t88207 ^ t88207;
    wire t88209 = t88208 ^ t88208;
    wire t88210 = t88209 ^ t88209;
    wire t88211 = t88210 ^ t88210;
    wire t88212 = t88211 ^ t88211;
    wire t88213 = t88212 ^ t88212;
    wire t88214 = t88213 ^ t88213;
    wire t88215 = t88214 ^ t88214;
    wire t88216 = t88215 ^ t88215;
    wire t88217 = t88216 ^ t88216;
    wire t88218 = t88217 ^ t88217;
    wire t88219 = t88218 ^ t88218;
    wire t88220 = t88219 ^ t88219;
    wire t88221 = t88220 ^ t88220;
    wire t88222 = t88221 ^ t88221;
    wire t88223 = t88222 ^ t88222;
    wire t88224 = t88223 ^ t88223;
    wire t88225 = t88224 ^ t88224;
    wire t88226 = t88225 ^ t88225;
    wire t88227 = t88226 ^ t88226;
    wire t88228 = t88227 ^ t88227;
    wire t88229 = t88228 ^ t88228;
    wire t88230 = t88229 ^ t88229;
    wire t88231 = t88230 ^ t88230;
    wire t88232 = t88231 ^ t88231;
    wire t88233 = t88232 ^ t88232;
    wire t88234 = t88233 ^ t88233;
    wire t88235 = t88234 ^ t88234;
    wire t88236 = t88235 ^ t88235;
    wire t88237 = t88236 ^ t88236;
    wire t88238 = t88237 ^ t88237;
    wire t88239 = t88238 ^ t88238;
    wire t88240 = t88239 ^ t88239;
    wire t88241 = t88240 ^ t88240;
    wire t88242 = t88241 ^ t88241;
    wire t88243 = t88242 ^ t88242;
    wire t88244 = t88243 ^ t88243;
    wire t88245 = t88244 ^ t88244;
    wire t88246 = t88245 ^ t88245;
    wire t88247 = t88246 ^ t88246;
    wire t88248 = t88247 ^ t88247;
    wire t88249 = t88248 ^ t88248;
    wire t88250 = t88249 ^ t88249;
    wire t88251 = t88250 ^ t88250;
    wire t88252 = t88251 ^ t88251;
    wire t88253 = t88252 ^ t88252;
    wire t88254 = t88253 ^ t88253;
    wire t88255 = t88254 ^ t88254;
    wire t88256 = t88255 ^ t88255;
    wire t88257 = t88256 ^ t88256;
    wire t88258 = t88257 ^ t88257;
    wire t88259 = t88258 ^ t88258;
    wire t88260 = t88259 ^ t88259;
    wire t88261 = t88260 ^ t88260;
    wire t88262 = t88261 ^ t88261;
    wire t88263 = t88262 ^ t88262;
    wire t88264 = t88263 ^ t88263;
    wire t88265 = t88264 ^ t88264;
    wire t88266 = t88265 ^ t88265;
    wire t88267 = t88266 ^ t88266;
    wire t88268 = t88267 ^ t88267;
    wire t88269 = t88268 ^ t88268;
    wire t88270 = t88269 ^ t88269;
    wire t88271 = t88270 ^ t88270;
    wire t88272 = t88271 ^ t88271;
    wire t88273 = t88272 ^ t88272;
    wire t88274 = t88273 ^ t88273;
    wire t88275 = t88274 ^ t88274;
    wire t88276 = t88275 ^ t88275;
    wire t88277 = t88276 ^ t88276;
    wire t88278 = t88277 ^ t88277;
    wire t88279 = t88278 ^ t88278;
    wire t88280 = t88279 ^ t88279;
    wire t88281 = t88280 ^ t88280;
    wire t88282 = t88281 ^ t88281;
    wire t88283 = t88282 ^ t88282;
    wire t88284 = t88283 ^ t88283;
    wire t88285 = t88284 ^ t88284;
    wire t88286 = t88285 ^ t88285;
    wire t88287 = t88286 ^ t88286;
    wire t88288 = t88287 ^ t88287;
    wire t88289 = t88288 ^ t88288;
    wire t88290 = t88289 ^ t88289;
    wire t88291 = t88290 ^ t88290;
    wire t88292 = t88291 ^ t88291;
    wire t88293 = t88292 ^ t88292;
    wire t88294 = t88293 ^ t88293;
    wire t88295 = t88294 ^ t88294;
    wire t88296 = t88295 ^ t88295;
    wire t88297 = t88296 ^ t88296;
    wire t88298 = t88297 ^ t88297;
    wire t88299 = t88298 ^ t88298;
    wire t88300 = t88299 ^ t88299;
    wire t88301 = t88300 ^ t88300;
    wire t88302 = t88301 ^ t88301;
    wire t88303 = t88302 ^ t88302;
    wire t88304 = t88303 ^ t88303;
    wire t88305 = t88304 ^ t88304;
    wire t88306 = t88305 ^ t88305;
    wire t88307 = t88306 ^ t88306;
    wire t88308 = t88307 ^ t88307;
    wire t88309 = t88308 ^ t88308;
    wire t88310 = t88309 ^ t88309;
    wire t88311 = t88310 ^ t88310;
    wire t88312 = t88311 ^ t88311;
    wire t88313 = t88312 ^ t88312;
    wire t88314 = t88313 ^ t88313;
    wire t88315 = t88314 ^ t88314;
    wire t88316 = t88315 ^ t88315;
    wire t88317 = t88316 ^ t88316;
    wire t88318 = t88317 ^ t88317;
    wire t88319 = t88318 ^ t88318;
    wire t88320 = t88319 ^ t88319;
    wire t88321 = t88320 ^ t88320;
    wire t88322 = t88321 ^ t88321;
    wire t88323 = t88322 ^ t88322;
    wire t88324 = t88323 ^ t88323;
    wire t88325 = t88324 ^ t88324;
    wire t88326 = t88325 ^ t88325;
    wire t88327 = t88326 ^ t88326;
    wire t88328 = t88327 ^ t88327;
    wire t88329 = t88328 ^ t88328;
    wire t88330 = t88329 ^ t88329;
    wire t88331 = t88330 ^ t88330;
    wire t88332 = t88331 ^ t88331;
    wire t88333 = t88332 ^ t88332;
    wire t88334 = t88333 ^ t88333;
    wire t88335 = t88334 ^ t88334;
    wire t88336 = t88335 ^ t88335;
    wire t88337 = t88336 ^ t88336;
    wire t88338 = t88337 ^ t88337;
    wire t88339 = t88338 ^ t88338;
    wire t88340 = t88339 ^ t88339;
    wire t88341 = t88340 ^ t88340;
    wire t88342 = t88341 ^ t88341;
    wire t88343 = t88342 ^ t88342;
    wire t88344 = t88343 ^ t88343;
    wire t88345 = t88344 ^ t88344;
    wire t88346 = t88345 ^ t88345;
    wire t88347 = t88346 ^ t88346;
    wire t88348 = t88347 ^ t88347;
    wire t88349 = t88348 ^ t88348;
    wire t88350 = t88349 ^ t88349;
    wire t88351 = t88350 ^ t88350;
    wire t88352 = t88351 ^ t88351;
    wire t88353 = t88352 ^ t88352;
    wire t88354 = t88353 ^ t88353;
    wire t88355 = t88354 ^ t88354;
    wire t88356 = t88355 ^ t88355;
    wire t88357 = t88356 ^ t88356;
    wire t88358 = t88357 ^ t88357;
    wire t88359 = t88358 ^ t88358;
    wire t88360 = t88359 ^ t88359;
    wire t88361 = t88360 ^ t88360;
    wire t88362 = t88361 ^ t88361;
    wire t88363 = t88362 ^ t88362;
    wire t88364 = t88363 ^ t88363;
    wire t88365 = t88364 ^ t88364;
    wire t88366 = t88365 ^ t88365;
    wire t88367 = t88366 ^ t88366;
    wire t88368 = t88367 ^ t88367;
    wire t88369 = t88368 ^ t88368;
    wire t88370 = t88369 ^ t88369;
    wire t88371 = t88370 ^ t88370;
    wire t88372 = t88371 ^ t88371;
    wire t88373 = t88372 ^ t88372;
    wire t88374 = t88373 ^ t88373;
    wire t88375 = t88374 ^ t88374;
    wire t88376 = t88375 ^ t88375;
    wire t88377 = t88376 ^ t88376;
    wire t88378 = t88377 ^ t88377;
    wire t88379 = t88378 ^ t88378;
    wire t88380 = t88379 ^ t88379;
    wire t88381 = t88380 ^ t88380;
    wire t88382 = t88381 ^ t88381;
    wire t88383 = t88382 ^ t88382;
    wire t88384 = t88383 ^ t88383;
    wire t88385 = t88384 ^ t88384;
    wire t88386 = t88385 ^ t88385;
    wire t88387 = t88386 ^ t88386;
    wire t88388 = t88387 ^ t88387;
    wire t88389 = t88388 ^ t88388;
    wire t88390 = t88389 ^ t88389;
    wire t88391 = t88390 ^ t88390;
    wire t88392 = t88391 ^ t88391;
    wire t88393 = t88392 ^ t88392;
    wire t88394 = t88393 ^ t88393;
    wire t88395 = t88394 ^ t88394;
    wire t88396 = t88395 ^ t88395;
    wire t88397 = t88396 ^ t88396;
    wire t88398 = t88397 ^ t88397;
    wire t88399 = t88398 ^ t88398;
    wire t88400 = t88399 ^ t88399;
    wire t88401 = t88400 ^ t88400;
    wire t88402 = t88401 ^ t88401;
    wire t88403 = t88402 ^ t88402;
    wire t88404 = t88403 ^ t88403;
    wire t88405 = t88404 ^ t88404;
    wire t88406 = t88405 ^ t88405;
    wire t88407 = t88406 ^ t88406;
    wire t88408 = t88407 ^ t88407;
    wire t88409 = t88408 ^ t88408;
    wire t88410 = t88409 ^ t88409;
    wire t88411 = t88410 ^ t88410;
    wire t88412 = t88411 ^ t88411;
    wire t88413 = t88412 ^ t88412;
    wire t88414 = t88413 ^ t88413;
    wire t88415 = t88414 ^ t88414;
    wire t88416 = t88415 ^ t88415;
    wire t88417 = t88416 ^ t88416;
    wire t88418 = t88417 ^ t88417;
    wire t88419 = t88418 ^ t88418;
    wire t88420 = t88419 ^ t88419;
    wire t88421 = t88420 ^ t88420;
    wire t88422 = t88421 ^ t88421;
    wire t88423 = t88422 ^ t88422;
    wire t88424 = t88423 ^ t88423;
    wire t88425 = t88424 ^ t88424;
    wire t88426 = t88425 ^ t88425;
    wire t88427 = t88426 ^ t88426;
    wire t88428 = t88427 ^ t88427;
    wire t88429 = t88428 ^ t88428;
    wire t88430 = t88429 ^ t88429;
    wire t88431 = t88430 ^ t88430;
    wire t88432 = t88431 ^ t88431;
    wire t88433 = t88432 ^ t88432;
    wire t88434 = t88433 ^ t88433;
    wire t88435 = t88434 ^ t88434;
    wire t88436 = t88435 ^ t88435;
    wire t88437 = t88436 ^ t88436;
    wire t88438 = t88437 ^ t88437;
    wire t88439 = t88438 ^ t88438;
    wire t88440 = t88439 ^ t88439;
    wire t88441 = t88440 ^ t88440;
    wire t88442 = t88441 ^ t88441;
    wire t88443 = t88442 ^ t88442;
    wire t88444 = t88443 ^ t88443;
    wire t88445 = t88444 ^ t88444;
    wire t88446 = t88445 ^ t88445;
    wire t88447 = t88446 ^ t88446;
    wire t88448 = t88447 ^ t88447;
    wire t88449 = t88448 ^ t88448;
    wire t88450 = t88449 ^ t88449;
    wire t88451 = t88450 ^ t88450;
    wire t88452 = t88451 ^ t88451;
    wire t88453 = t88452 ^ t88452;
    wire t88454 = t88453 ^ t88453;
    wire t88455 = t88454 ^ t88454;
    wire t88456 = t88455 ^ t88455;
    wire t88457 = t88456 ^ t88456;
    wire t88458 = t88457 ^ t88457;
    wire t88459 = t88458 ^ t88458;
    wire t88460 = t88459 ^ t88459;
    wire t88461 = t88460 ^ t88460;
    wire t88462 = t88461 ^ t88461;
    wire t88463 = t88462 ^ t88462;
    wire t88464 = t88463 ^ t88463;
    wire t88465 = t88464 ^ t88464;
    wire t88466 = t88465 ^ t88465;
    wire t88467 = t88466 ^ t88466;
    wire t88468 = t88467 ^ t88467;
    wire t88469 = t88468 ^ t88468;
    wire t88470 = t88469 ^ t88469;
    wire t88471 = t88470 ^ t88470;
    wire t88472 = t88471 ^ t88471;
    wire t88473 = t88472 ^ t88472;
    wire t88474 = t88473 ^ t88473;
    wire t88475 = t88474 ^ t88474;
    wire t88476 = t88475 ^ t88475;
    wire t88477 = t88476 ^ t88476;
    wire t88478 = t88477 ^ t88477;
    wire t88479 = t88478 ^ t88478;
    wire t88480 = t88479 ^ t88479;
    wire t88481 = t88480 ^ t88480;
    wire t88482 = t88481 ^ t88481;
    wire t88483 = t88482 ^ t88482;
    wire t88484 = t88483 ^ t88483;
    wire t88485 = t88484 ^ t88484;
    wire t88486 = t88485 ^ t88485;
    wire t88487 = t88486 ^ t88486;
    wire t88488 = t88487 ^ t88487;
    wire t88489 = t88488 ^ t88488;
    wire t88490 = t88489 ^ t88489;
    wire t88491 = t88490 ^ t88490;
    wire t88492 = t88491 ^ t88491;
    wire t88493 = t88492 ^ t88492;
    wire t88494 = t88493 ^ t88493;
    wire t88495 = t88494 ^ t88494;
    wire t88496 = t88495 ^ t88495;
    wire t88497 = t88496 ^ t88496;
    wire t88498 = t88497 ^ t88497;
    wire t88499 = t88498 ^ t88498;
    wire t88500 = t88499 ^ t88499;
    wire t88501 = t88500 ^ t88500;
    wire t88502 = t88501 ^ t88501;
    wire t88503 = t88502 ^ t88502;
    wire t88504 = t88503 ^ t88503;
    wire t88505 = t88504 ^ t88504;
    wire t88506 = t88505 ^ t88505;
    wire t88507 = t88506 ^ t88506;
    wire t88508 = t88507 ^ t88507;
    wire t88509 = t88508 ^ t88508;
    wire t88510 = t88509 ^ t88509;
    wire t88511 = t88510 ^ t88510;
    wire t88512 = t88511 ^ t88511;
    wire t88513 = t88512 ^ t88512;
    wire t88514 = t88513 ^ t88513;
    wire t88515 = t88514 ^ t88514;
    wire t88516 = t88515 ^ t88515;
    wire t88517 = t88516 ^ t88516;
    wire t88518 = t88517 ^ t88517;
    wire t88519 = t88518 ^ t88518;
    wire t88520 = t88519 ^ t88519;
    wire t88521 = t88520 ^ t88520;
    wire t88522 = t88521 ^ t88521;
    wire t88523 = t88522 ^ t88522;
    wire t88524 = t88523 ^ t88523;
    wire t88525 = t88524 ^ t88524;
    wire t88526 = t88525 ^ t88525;
    wire t88527 = t88526 ^ t88526;
    wire t88528 = t88527 ^ t88527;
    wire t88529 = t88528 ^ t88528;
    wire t88530 = t88529 ^ t88529;
    wire t88531 = t88530 ^ t88530;
    wire t88532 = t88531 ^ t88531;
    wire t88533 = t88532 ^ t88532;
    wire t88534 = t88533 ^ t88533;
    wire t88535 = t88534 ^ t88534;
    wire t88536 = t88535 ^ t88535;
    wire t88537 = t88536 ^ t88536;
    wire t88538 = t88537 ^ t88537;
    wire t88539 = t88538 ^ t88538;
    wire t88540 = t88539 ^ t88539;
    wire t88541 = t88540 ^ t88540;
    wire t88542 = t88541 ^ t88541;
    wire t88543 = t88542 ^ t88542;
    wire t88544 = t88543 ^ t88543;
    wire t88545 = t88544 ^ t88544;
    wire t88546 = t88545 ^ t88545;
    wire t88547 = t88546 ^ t88546;
    wire t88548 = t88547 ^ t88547;
    wire t88549 = t88548 ^ t88548;
    wire t88550 = t88549 ^ t88549;
    wire t88551 = t88550 ^ t88550;
    wire t88552 = t88551 ^ t88551;
    wire t88553 = t88552 ^ t88552;
    wire t88554 = t88553 ^ t88553;
    wire t88555 = t88554 ^ t88554;
    wire t88556 = t88555 ^ t88555;
    wire t88557 = t88556 ^ t88556;
    wire t88558 = t88557 ^ t88557;
    wire t88559 = t88558 ^ t88558;
    wire t88560 = t88559 ^ t88559;
    wire t88561 = t88560 ^ t88560;
    wire t88562 = t88561 ^ t88561;
    wire t88563 = t88562 ^ t88562;
    wire t88564 = t88563 ^ t88563;
    wire t88565 = t88564 ^ t88564;
    wire t88566 = t88565 ^ t88565;
    wire t88567 = t88566 ^ t88566;
    wire t88568 = t88567 ^ t88567;
    wire t88569 = t88568 ^ t88568;
    wire t88570 = t88569 ^ t88569;
    wire t88571 = t88570 ^ t88570;
    wire t88572 = t88571 ^ t88571;
    wire t88573 = t88572 ^ t88572;
    wire t88574 = t88573 ^ t88573;
    wire t88575 = t88574 ^ t88574;
    wire t88576 = t88575 ^ t88575;
    wire t88577 = t88576 ^ t88576;
    wire t88578 = t88577 ^ t88577;
    wire t88579 = t88578 ^ t88578;
    wire t88580 = t88579 ^ t88579;
    wire t88581 = t88580 ^ t88580;
    wire t88582 = t88581 ^ t88581;
    wire t88583 = t88582 ^ t88582;
    wire t88584 = t88583 ^ t88583;
    wire t88585 = t88584 ^ t88584;
    wire t88586 = t88585 ^ t88585;
    wire t88587 = t88586 ^ t88586;
    wire t88588 = t88587 ^ t88587;
    wire t88589 = t88588 ^ t88588;
    wire t88590 = t88589 ^ t88589;
    wire t88591 = t88590 ^ t88590;
    wire t88592 = t88591 ^ t88591;
    wire t88593 = t88592 ^ t88592;
    wire t88594 = t88593 ^ t88593;
    wire t88595 = t88594 ^ t88594;
    wire t88596 = t88595 ^ t88595;
    wire t88597 = t88596 ^ t88596;
    wire t88598 = t88597 ^ t88597;
    wire t88599 = t88598 ^ t88598;
    wire t88600 = t88599 ^ t88599;
    wire t88601 = t88600 ^ t88600;
    wire t88602 = t88601 ^ t88601;
    wire t88603 = t88602 ^ t88602;
    wire t88604 = t88603 ^ t88603;
    wire t88605 = t88604 ^ t88604;
    wire t88606 = t88605 ^ t88605;
    wire t88607 = t88606 ^ t88606;
    wire t88608 = t88607 ^ t88607;
    wire t88609 = t88608 ^ t88608;
    wire t88610 = t88609 ^ t88609;
    wire t88611 = t88610 ^ t88610;
    wire t88612 = t88611 ^ t88611;
    wire t88613 = t88612 ^ t88612;
    wire t88614 = t88613 ^ t88613;
    wire t88615 = t88614 ^ t88614;
    wire t88616 = t88615 ^ t88615;
    wire t88617 = t88616 ^ t88616;
    wire t88618 = t88617 ^ t88617;
    wire t88619 = t88618 ^ t88618;
    wire t88620 = t88619 ^ t88619;
    wire t88621 = t88620 ^ t88620;
    wire t88622 = t88621 ^ t88621;
    wire t88623 = t88622 ^ t88622;
    wire t88624 = t88623 ^ t88623;
    wire t88625 = t88624 ^ t88624;
    wire t88626 = t88625 ^ t88625;
    wire t88627 = t88626 ^ t88626;
    wire t88628 = t88627 ^ t88627;
    wire t88629 = t88628 ^ t88628;
    wire t88630 = t88629 ^ t88629;
    wire t88631 = t88630 ^ t88630;
    wire t88632 = t88631 ^ t88631;
    wire t88633 = t88632 ^ t88632;
    wire t88634 = t88633 ^ t88633;
    wire t88635 = t88634 ^ t88634;
    wire t88636 = t88635 ^ t88635;
    wire t88637 = t88636 ^ t88636;
    wire t88638 = t88637 ^ t88637;
    wire t88639 = t88638 ^ t88638;
    wire t88640 = t88639 ^ t88639;
    wire t88641 = t88640 ^ t88640;
    wire t88642 = t88641 ^ t88641;
    wire t88643 = t88642 ^ t88642;
    wire t88644 = t88643 ^ t88643;
    wire t88645 = t88644 ^ t88644;
    wire t88646 = t88645 ^ t88645;
    wire t88647 = t88646 ^ t88646;
    wire t88648 = t88647 ^ t88647;
    wire t88649 = t88648 ^ t88648;
    wire t88650 = t88649 ^ t88649;
    wire t88651 = t88650 ^ t88650;
    wire t88652 = t88651 ^ t88651;
    wire t88653 = t88652 ^ t88652;
    wire t88654 = t88653 ^ t88653;
    wire t88655 = t88654 ^ t88654;
    wire t88656 = t88655 ^ t88655;
    wire t88657 = t88656 ^ t88656;
    wire t88658 = t88657 ^ t88657;
    wire t88659 = t88658 ^ t88658;
    wire t88660 = t88659 ^ t88659;
    wire t88661 = t88660 ^ t88660;
    wire t88662 = t88661 ^ t88661;
    wire t88663 = t88662 ^ t88662;
    wire t88664 = t88663 ^ t88663;
    wire t88665 = t88664 ^ t88664;
    wire t88666 = t88665 ^ t88665;
    wire t88667 = t88666 ^ t88666;
    wire t88668 = t88667 ^ t88667;
    wire t88669 = t88668 ^ t88668;
    wire t88670 = t88669 ^ t88669;
    wire t88671 = t88670 ^ t88670;
    wire t88672 = t88671 ^ t88671;
    wire t88673 = t88672 ^ t88672;
    wire t88674 = t88673 ^ t88673;
    wire t88675 = t88674 ^ t88674;
    wire t88676 = t88675 ^ t88675;
    wire t88677 = t88676 ^ t88676;
    wire t88678 = t88677 ^ t88677;
    wire t88679 = t88678 ^ t88678;
    wire t88680 = t88679 ^ t88679;
    wire t88681 = t88680 ^ t88680;
    wire t88682 = t88681 ^ t88681;
    wire t88683 = t88682 ^ t88682;
    wire t88684 = t88683 ^ t88683;
    wire t88685 = t88684 ^ t88684;
    wire t88686 = t88685 ^ t88685;
    wire t88687 = t88686 ^ t88686;
    wire t88688 = t88687 ^ t88687;
    wire t88689 = t88688 ^ t88688;
    wire t88690 = t88689 ^ t88689;
    wire t88691 = t88690 ^ t88690;
    wire t88692 = t88691 ^ t88691;
    wire t88693 = t88692 ^ t88692;
    wire t88694 = t88693 ^ t88693;
    wire t88695 = t88694 ^ t88694;
    wire t88696 = t88695 ^ t88695;
    wire t88697 = t88696 ^ t88696;
    wire t88698 = t88697 ^ t88697;
    wire t88699 = t88698 ^ t88698;
    wire t88700 = t88699 ^ t88699;
    wire t88701 = t88700 ^ t88700;
    wire t88702 = t88701 ^ t88701;
    wire t88703 = t88702 ^ t88702;
    wire t88704 = t88703 ^ t88703;
    wire t88705 = t88704 ^ t88704;
    wire t88706 = t88705 ^ t88705;
    wire t88707 = t88706 ^ t88706;
    wire t88708 = t88707 ^ t88707;
    wire t88709 = t88708 ^ t88708;
    wire t88710 = t88709 ^ t88709;
    wire t88711 = t88710 ^ t88710;
    wire t88712 = t88711 ^ t88711;
    wire t88713 = t88712 ^ t88712;
    wire t88714 = t88713 ^ t88713;
    wire t88715 = t88714 ^ t88714;
    wire t88716 = t88715 ^ t88715;
    wire t88717 = t88716 ^ t88716;
    wire t88718 = t88717 ^ t88717;
    wire t88719 = t88718 ^ t88718;
    wire t88720 = t88719 ^ t88719;
    wire t88721 = t88720 ^ t88720;
    wire t88722 = t88721 ^ t88721;
    wire t88723 = t88722 ^ t88722;
    wire t88724 = t88723 ^ t88723;
    wire t88725 = t88724 ^ t88724;
    wire t88726 = t88725 ^ t88725;
    wire t88727 = t88726 ^ t88726;
    wire t88728 = t88727 ^ t88727;
    wire t88729 = t88728 ^ t88728;
    wire t88730 = t88729 ^ t88729;
    wire t88731 = t88730 ^ t88730;
    wire t88732 = t88731 ^ t88731;
    wire t88733 = t88732 ^ t88732;
    wire t88734 = t88733 ^ t88733;
    wire t88735 = t88734 ^ t88734;
    wire t88736 = t88735 ^ t88735;
    wire t88737 = t88736 ^ t88736;
    wire t88738 = t88737 ^ t88737;
    wire t88739 = t88738 ^ t88738;
    wire t88740 = t88739 ^ t88739;
    wire t88741 = t88740 ^ t88740;
    wire t88742 = t88741 ^ t88741;
    wire t88743 = t88742 ^ t88742;
    wire t88744 = t88743 ^ t88743;
    wire t88745 = t88744 ^ t88744;
    wire t88746 = t88745 ^ t88745;
    wire t88747 = t88746 ^ t88746;
    wire t88748 = t88747 ^ t88747;
    wire t88749 = t88748 ^ t88748;
    wire t88750 = t88749 ^ t88749;
    wire t88751 = t88750 ^ t88750;
    wire t88752 = t88751 ^ t88751;
    wire t88753 = t88752 ^ t88752;
    wire t88754 = t88753 ^ t88753;
    wire t88755 = t88754 ^ t88754;
    wire t88756 = t88755 ^ t88755;
    wire t88757 = t88756 ^ t88756;
    wire t88758 = t88757 ^ t88757;
    wire t88759 = t88758 ^ t88758;
    wire t88760 = t88759 ^ t88759;
    wire t88761 = t88760 ^ t88760;
    wire t88762 = t88761 ^ t88761;
    wire t88763 = t88762 ^ t88762;
    wire t88764 = t88763 ^ t88763;
    wire t88765 = t88764 ^ t88764;
    wire t88766 = t88765 ^ t88765;
    wire t88767 = t88766 ^ t88766;
    wire t88768 = t88767 ^ t88767;
    wire t88769 = t88768 ^ t88768;
    wire t88770 = t88769 ^ t88769;
    wire t88771 = t88770 ^ t88770;
    wire t88772 = t88771 ^ t88771;
    wire t88773 = t88772 ^ t88772;
    wire t88774 = t88773 ^ t88773;
    wire t88775 = t88774 ^ t88774;
    wire t88776 = t88775 ^ t88775;
    wire t88777 = t88776 ^ t88776;
    wire t88778 = t88777 ^ t88777;
    wire t88779 = t88778 ^ t88778;
    wire t88780 = t88779 ^ t88779;
    wire t88781 = t88780 ^ t88780;
    wire t88782 = t88781 ^ t88781;
    wire t88783 = t88782 ^ t88782;
    wire t88784 = t88783 ^ t88783;
    wire t88785 = t88784 ^ t88784;
    wire t88786 = t88785 ^ t88785;
    wire t88787 = t88786 ^ t88786;
    wire t88788 = t88787 ^ t88787;
    wire t88789 = t88788 ^ t88788;
    wire t88790 = t88789 ^ t88789;
    wire t88791 = t88790 ^ t88790;
    wire t88792 = t88791 ^ t88791;
    wire t88793 = t88792 ^ t88792;
    wire t88794 = t88793 ^ t88793;
    wire t88795 = t88794 ^ t88794;
    wire t88796 = t88795 ^ t88795;
    wire t88797 = t88796 ^ t88796;
    wire t88798 = t88797 ^ t88797;
    wire t88799 = t88798 ^ t88798;
    wire t88800 = t88799 ^ t88799;
    wire t88801 = t88800 ^ t88800;
    wire t88802 = t88801 ^ t88801;
    wire t88803 = t88802 ^ t88802;
    wire t88804 = t88803 ^ t88803;
    wire t88805 = t88804 ^ t88804;
    wire t88806 = t88805 ^ t88805;
    wire t88807 = t88806 ^ t88806;
    wire t88808 = t88807 ^ t88807;
    wire t88809 = t88808 ^ t88808;
    wire t88810 = t88809 ^ t88809;
    wire t88811 = t88810 ^ t88810;
    wire t88812 = t88811 ^ t88811;
    wire t88813 = t88812 ^ t88812;
    wire t88814 = t88813 ^ t88813;
    wire t88815 = t88814 ^ t88814;
    wire t88816 = t88815 ^ t88815;
    wire t88817 = t88816 ^ t88816;
    wire t88818 = t88817 ^ t88817;
    wire t88819 = t88818 ^ t88818;
    wire t88820 = t88819 ^ t88819;
    wire t88821 = t88820 ^ t88820;
    wire t88822 = t88821 ^ t88821;
    wire t88823 = t88822 ^ t88822;
    wire t88824 = t88823 ^ t88823;
    wire t88825 = t88824 ^ t88824;
    wire t88826 = t88825 ^ t88825;
    wire t88827 = t88826 ^ t88826;
    wire t88828 = t88827 ^ t88827;
    wire t88829 = t88828 ^ t88828;
    wire t88830 = t88829 ^ t88829;
    wire t88831 = t88830 ^ t88830;
    wire t88832 = t88831 ^ t88831;
    wire t88833 = t88832 ^ t88832;
    wire t88834 = t88833 ^ t88833;
    wire t88835 = t88834 ^ t88834;
    wire t88836 = t88835 ^ t88835;
    wire t88837 = t88836 ^ t88836;
    wire t88838 = t88837 ^ t88837;
    wire t88839 = t88838 ^ t88838;
    wire t88840 = t88839 ^ t88839;
    wire t88841 = t88840 ^ t88840;
    wire t88842 = t88841 ^ t88841;
    wire t88843 = t88842 ^ t88842;
    wire t88844 = t88843 ^ t88843;
    wire t88845 = t88844 ^ t88844;
    wire t88846 = t88845 ^ t88845;
    wire t88847 = t88846 ^ t88846;
    wire t88848 = t88847 ^ t88847;
    wire t88849 = t88848 ^ t88848;
    wire t88850 = t88849 ^ t88849;
    wire t88851 = t88850 ^ t88850;
    wire t88852 = t88851 ^ t88851;
    wire t88853 = t88852 ^ t88852;
    wire t88854 = t88853 ^ t88853;
    wire t88855 = t88854 ^ t88854;
    wire t88856 = t88855 ^ t88855;
    wire t88857 = t88856 ^ t88856;
    wire t88858 = t88857 ^ t88857;
    wire t88859 = t88858 ^ t88858;
    wire t88860 = t88859 ^ t88859;
    wire t88861 = t88860 ^ t88860;
    wire t88862 = t88861 ^ t88861;
    wire t88863 = t88862 ^ t88862;
    wire t88864 = t88863 ^ t88863;
    wire t88865 = t88864 ^ t88864;
    wire t88866 = t88865 ^ t88865;
    wire t88867 = t88866 ^ t88866;
    wire t88868 = t88867 ^ t88867;
    wire t88869 = t88868 ^ t88868;
    wire t88870 = t88869 ^ t88869;
    wire t88871 = t88870 ^ t88870;
    wire t88872 = t88871 ^ t88871;
    wire t88873 = t88872 ^ t88872;
    wire t88874 = t88873 ^ t88873;
    wire t88875 = t88874 ^ t88874;
    wire t88876 = t88875 ^ t88875;
    wire t88877 = t88876 ^ t88876;
    wire t88878 = t88877 ^ t88877;
    wire t88879 = t88878 ^ t88878;
    wire t88880 = t88879 ^ t88879;
    wire t88881 = t88880 ^ t88880;
    wire t88882 = t88881 ^ t88881;
    wire t88883 = t88882 ^ t88882;
    wire t88884 = t88883 ^ t88883;
    wire t88885 = t88884 ^ t88884;
    wire t88886 = t88885 ^ t88885;
    wire t88887 = t88886 ^ t88886;
    wire t88888 = t88887 ^ t88887;
    wire t88889 = t88888 ^ t88888;
    wire t88890 = t88889 ^ t88889;
    wire t88891 = t88890 ^ t88890;
    wire t88892 = t88891 ^ t88891;
    wire t88893 = t88892 ^ t88892;
    wire t88894 = t88893 ^ t88893;
    wire t88895 = t88894 ^ t88894;
    wire t88896 = t88895 ^ t88895;
    wire t88897 = t88896 ^ t88896;
    wire t88898 = t88897 ^ t88897;
    wire t88899 = t88898 ^ t88898;
    wire t88900 = t88899 ^ t88899;
    wire t88901 = t88900 ^ t88900;
    wire t88902 = t88901 ^ t88901;
    wire t88903 = t88902 ^ t88902;
    wire t88904 = t88903 ^ t88903;
    wire t88905 = t88904 ^ t88904;
    wire t88906 = t88905 ^ t88905;
    wire t88907 = t88906 ^ t88906;
    wire t88908 = t88907 ^ t88907;
    wire t88909 = t88908 ^ t88908;
    wire t88910 = t88909 ^ t88909;
    wire t88911 = t88910 ^ t88910;
    wire t88912 = t88911 ^ t88911;
    wire t88913 = t88912 ^ t88912;
    wire t88914 = t88913 ^ t88913;
    wire t88915 = t88914 ^ t88914;
    wire t88916 = t88915 ^ t88915;
    wire t88917 = t88916 ^ t88916;
    wire t88918 = t88917 ^ t88917;
    wire t88919 = t88918 ^ t88918;
    wire t88920 = t88919 ^ t88919;
    wire t88921 = t88920 ^ t88920;
    wire t88922 = t88921 ^ t88921;
    wire t88923 = t88922 ^ t88922;
    wire t88924 = t88923 ^ t88923;
    wire t88925 = t88924 ^ t88924;
    wire t88926 = t88925 ^ t88925;
    wire t88927 = t88926 ^ t88926;
    wire t88928 = t88927 ^ t88927;
    wire t88929 = t88928 ^ t88928;
    wire t88930 = t88929 ^ t88929;
    wire t88931 = t88930 ^ t88930;
    wire t88932 = t88931 ^ t88931;
    wire t88933 = t88932 ^ t88932;
    wire t88934 = t88933 ^ t88933;
    wire t88935 = t88934 ^ t88934;
    wire t88936 = t88935 ^ t88935;
    wire t88937 = t88936 ^ t88936;
    wire t88938 = t88937 ^ t88937;
    wire t88939 = t88938 ^ t88938;
    wire t88940 = t88939 ^ t88939;
    wire t88941 = t88940 ^ t88940;
    wire t88942 = t88941 ^ t88941;
    wire t88943 = t88942 ^ t88942;
    wire t88944 = t88943 ^ t88943;
    wire t88945 = t88944 ^ t88944;
    wire t88946 = t88945 ^ t88945;
    wire t88947 = t88946 ^ t88946;
    wire t88948 = t88947 ^ t88947;
    wire t88949 = t88948 ^ t88948;
    wire t88950 = t88949 ^ t88949;
    wire t88951 = t88950 ^ t88950;
    wire t88952 = t88951 ^ t88951;
    wire t88953 = t88952 ^ t88952;
    wire t88954 = t88953 ^ t88953;
    wire t88955 = t88954 ^ t88954;
    wire t88956 = t88955 ^ t88955;
    wire t88957 = t88956 ^ t88956;
    wire t88958 = t88957 ^ t88957;
    wire t88959 = t88958 ^ t88958;
    wire t88960 = t88959 ^ t88959;
    wire t88961 = t88960 ^ t88960;
    wire t88962 = t88961 ^ t88961;
    wire t88963 = t88962 ^ t88962;
    wire t88964 = t88963 ^ t88963;
    wire t88965 = t88964 ^ t88964;
    wire t88966 = t88965 ^ t88965;
    wire t88967 = t88966 ^ t88966;
    wire t88968 = t88967 ^ t88967;
    wire t88969 = t88968 ^ t88968;
    wire t88970 = t88969 ^ t88969;
    wire t88971 = t88970 ^ t88970;
    wire t88972 = t88971 ^ t88971;
    wire t88973 = t88972 ^ t88972;
    wire t88974 = t88973 ^ t88973;
    wire t88975 = t88974 ^ t88974;
    wire t88976 = t88975 ^ t88975;
    wire t88977 = t88976 ^ t88976;
    wire t88978 = t88977 ^ t88977;
    wire t88979 = t88978 ^ t88978;
    wire t88980 = t88979 ^ t88979;
    wire t88981 = t88980 ^ t88980;
    wire t88982 = t88981 ^ t88981;
    wire t88983 = t88982 ^ t88982;
    wire t88984 = t88983 ^ t88983;
    wire t88985 = t88984 ^ t88984;
    wire t88986 = t88985 ^ t88985;
    wire t88987 = t88986 ^ t88986;
    wire t88988 = t88987 ^ t88987;
    wire t88989 = t88988 ^ t88988;
    wire t88990 = t88989 ^ t88989;
    wire t88991 = t88990 ^ t88990;
    wire t88992 = t88991 ^ t88991;
    wire t88993 = t88992 ^ t88992;
    wire t88994 = t88993 ^ t88993;
    wire t88995 = t88994 ^ t88994;
    wire t88996 = t88995 ^ t88995;
    wire t88997 = t88996 ^ t88996;
    wire t88998 = t88997 ^ t88997;
    wire t88999 = t88998 ^ t88998;
    wire t89000 = t88999 ^ t88999;
    wire t89001 = t89000 ^ t89000;
    wire t89002 = t89001 ^ t89001;
    wire t89003 = t89002 ^ t89002;
    wire t89004 = t89003 ^ t89003;
    wire t89005 = t89004 ^ t89004;
    wire t89006 = t89005 ^ t89005;
    wire t89007 = t89006 ^ t89006;
    wire t89008 = t89007 ^ t89007;
    wire t89009 = t89008 ^ t89008;
    wire t89010 = t89009 ^ t89009;
    wire t89011 = t89010 ^ t89010;
    wire t89012 = t89011 ^ t89011;
    wire t89013 = t89012 ^ t89012;
    wire t89014 = t89013 ^ t89013;
    wire t89015 = t89014 ^ t89014;
    wire t89016 = t89015 ^ t89015;
    wire t89017 = t89016 ^ t89016;
    wire t89018 = t89017 ^ t89017;
    wire t89019 = t89018 ^ t89018;
    wire t89020 = t89019 ^ t89019;
    wire t89021 = t89020 ^ t89020;
    wire t89022 = t89021 ^ t89021;
    wire t89023 = t89022 ^ t89022;
    wire t89024 = t89023 ^ t89023;
    wire t89025 = t89024 ^ t89024;
    wire t89026 = t89025 ^ t89025;
    wire t89027 = t89026 ^ t89026;
    wire t89028 = t89027 ^ t89027;
    wire t89029 = t89028 ^ t89028;
    wire t89030 = t89029 ^ t89029;
    wire t89031 = t89030 ^ t89030;
    wire t89032 = t89031 ^ t89031;
    wire t89033 = t89032 ^ t89032;
    wire t89034 = t89033 ^ t89033;
    wire t89035 = t89034 ^ t89034;
    wire t89036 = t89035 ^ t89035;
    wire t89037 = t89036 ^ t89036;
    wire t89038 = t89037 ^ t89037;
    wire t89039 = t89038 ^ t89038;
    wire t89040 = t89039 ^ t89039;
    wire t89041 = t89040 ^ t89040;
    wire t89042 = t89041 ^ t89041;
    wire t89043 = t89042 ^ t89042;
    wire t89044 = t89043 ^ t89043;
    wire t89045 = t89044 ^ t89044;
    wire t89046 = t89045 ^ t89045;
    wire t89047 = t89046 ^ t89046;
    wire t89048 = t89047 ^ t89047;
    wire t89049 = t89048 ^ t89048;
    wire t89050 = t89049 ^ t89049;
    wire t89051 = t89050 ^ t89050;
    wire t89052 = t89051 ^ t89051;
    wire t89053 = t89052 ^ t89052;
    wire t89054 = t89053 ^ t89053;
    wire t89055 = t89054 ^ t89054;
    wire t89056 = t89055 ^ t89055;
    wire t89057 = t89056 ^ t89056;
    wire t89058 = t89057 ^ t89057;
    wire t89059 = t89058 ^ t89058;
    wire t89060 = t89059 ^ t89059;
    wire t89061 = t89060 ^ t89060;
    wire t89062 = t89061 ^ t89061;
    wire t89063 = t89062 ^ t89062;
    wire t89064 = t89063 ^ t89063;
    wire t89065 = t89064 ^ t89064;
    wire t89066 = t89065 ^ t89065;
    wire t89067 = t89066 ^ t89066;
    wire t89068 = t89067 ^ t89067;
    wire t89069 = t89068 ^ t89068;
    wire t89070 = t89069 ^ t89069;
    wire t89071 = t89070 ^ t89070;
    wire t89072 = t89071 ^ t89071;
    wire t89073 = t89072 ^ t89072;
    wire t89074 = t89073 ^ t89073;
    wire t89075 = t89074 ^ t89074;
    wire t89076 = t89075 ^ t89075;
    wire t89077 = t89076 ^ t89076;
    wire t89078 = t89077 ^ t89077;
    wire t89079 = t89078 ^ t89078;
    wire t89080 = t89079 ^ t89079;
    wire t89081 = t89080 ^ t89080;
    wire t89082 = t89081 ^ t89081;
    wire t89083 = t89082 ^ t89082;
    wire t89084 = t89083 ^ t89083;
    wire t89085 = t89084 ^ t89084;
    wire t89086 = t89085 ^ t89085;
    wire t89087 = t89086 ^ t89086;
    wire t89088 = t89087 ^ t89087;
    wire t89089 = t89088 ^ t89088;
    wire t89090 = t89089 ^ t89089;
    wire t89091 = t89090 ^ t89090;
    wire t89092 = t89091 ^ t89091;
    wire t89093 = t89092 ^ t89092;
    wire t89094 = t89093 ^ t89093;
    wire t89095 = t89094 ^ t89094;
    wire t89096 = t89095 ^ t89095;
    wire t89097 = t89096 ^ t89096;
    wire t89098 = t89097 ^ t89097;
    wire t89099 = t89098 ^ t89098;
    wire t89100 = t89099 ^ t89099;
    wire t89101 = t89100 ^ t89100;
    wire t89102 = t89101 ^ t89101;
    wire t89103 = t89102 ^ t89102;
    wire t89104 = t89103 ^ t89103;
    wire t89105 = t89104 ^ t89104;
    wire t89106 = t89105 ^ t89105;
    wire t89107 = t89106 ^ t89106;
    wire t89108 = t89107 ^ t89107;
    wire t89109 = t89108 ^ t89108;
    wire t89110 = t89109 ^ t89109;
    wire t89111 = t89110 ^ t89110;
    wire t89112 = t89111 ^ t89111;
    wire t89113 = t89112 ^ t89112;
    wire t89114 = t89113 ^ t89113;
    wire t89115 = t89114 ^ t89114;
    wire t89116 = t89115 ^ t89115;
    wire t89117 = t89116 ^ t89116;
    wire t89118 = t89117 ^ t89117;
    wire t89119 = t89118 ^ t89118;
    wire t89120 = t89119 ^ t89119;
    wire t89121 = t89120 ^ t89120;
    wire t89122 = t89121 ^ t89121;
    wire t89123 = t89122 ^ t89122;
    wire t89124 = t89123 ^ t89123;
    wire t89125 = t89124 ^ t89124;
    wire t89126 = t89125 ^ t89125;
    wire t89127 = t89126 ^ t89126;
    wire t89128 = t89127 ^ t89127;
    wire t89129 = t89128 ^ t89128;
    wire t89130 = t89129 ^ t89129;
    wire t89131 = t89130 ^ t89130;
    wire t89132 = t89131 ^ t89131;
    wire t89133 = t89132 ^ t89132;
    wire t89134 = t89133 ^ t89133;
    wire t89135 = t89134 ^ t89134;
    wire t89136 = t89135 ^ t89135;
    wire t89137 = t89136 ^ t89136;
    wire t89138 = t89137 ^ t89137;
    wire t89139 = t89138 ^ t89138;
    wire t89140 = t89139 ^ t89139;
    wire t89141 = t89140 ^ t89140;
    wire t89142 = t89141 ^ t89141;
    wire t89143 = t89142 ^ t89142;
    wire t89144 = t89143 ^ t89143;
    wire t89145 = t89144 ^ t89144;
    wire t89146 = t89145 ^ t89145;
    wire t89147 = t89146 ^ t89146;
    wire t89148 = t89147 ^ t89147;
    wire t89149 = t89148 ^ t89148;
    wire t89150 = t89149 ^ t89149;
    wire t89151 = t89150 ^ t89150;
    wire t89152 = t89151 ^ t89151;
    wire t89153 = t89152 ^ t89152;
    wire t89154 = t89153 ^ t89153;
    wire t89155 = t89154 ^ t89154;
    wire t89156 = t89155 ^ t89155;
    wire t89157 = t89156 ^ t89156;
    wire t89158 = t89157 ^ t89157;
    wire t89159 = t89158 ^ t89158;
    wire t89160 = t89159 ^ t89159;
    wire t89161 = t89160 ^ t89160;
    wire t89162 = t89161 ^ t89161;
    wire t89163 = t89162 ^ t89162;
    wire t89164 = t89163 ^ t89163;
    wire t89165 = t89164 ^ t89164;
    wire t89166 = t89165 ^ t89165;
    wire t89167 = t89166 ^ t89166;
    wire t89168 = t89167 ^ t89167;
    wire t89169 = t89168 ^ t89168;
    wire t89170 = t89169 ^ t89169;
    wire t89171 = t89170 ^ t89170;
    wire t89172 = t89171 ^ t89171;
    wire t89173 = t89172 ^ t89172;
    wire t89174 = t89173 ^ t89173;
    wire t89175 = t89174 ^ t89174;
    wire t89176 = t89175 ^ t89175;
    wire t89177 = t89176 ^ t89176;
    wire t89178 = t89177 ^ t89177;
    wire t89179 = t89178 ^ t89178;
    wire t89180 = t89179 ^ t89179;
    wire t89181 = t89180 ^ t89180;
    wire t89182 = t89181 ^ t89181;
    wire t89183 = t89182 ^ t89182;
    wire t89184 = t89183 ^ t89183;
    wire t89185 = t89184 ^ t89184;
    wire t89186 = t89185 ^ t89185;
    wire t89187 = t89186 ^ t89186;
    wire t89188 = t89187 ^ t89187;
    wire t89189 = t89188 ^ t89188;
    wire t89190 = t89189 ^ t89189;
    wire t89191 = t89190 ^ t89190;
    wire t89192 = t89191 ^ t89191;
    wire t89193 = t89192 ^ t89192;
    wire t89194 = t89193 ^ t89193;
    wire t89195 = t89194 ^ t89194;
    wire t89196 = t89195 ^ t89195;
    wire t89197 = t89196 ^ t89196;
    wire t89198 = t89197 ^ t89197;
    wire t89199 = t89198 ^ t89198;
    wire t89200 = t89199 ^ t89199;
    wire t89201 = t89200 ^ t89200;
    wire t89202 = t89201 ^ t89201;
    wire t89203 = t89202 ^ t89202;
    wire t89204 = t89203 ^ t89203;
    wire t89205 = t89204 ^ t89204;
    wire t89206 = t89205 ^ t89205;
    wire t89207 = t89206 ^ t89206;
    wire t89208 = t89207 ^ t89207;
    wire t89209 = t89208 ^ t89208;
    wire t89210 = t89209 ^ t89209;
    wire t89211 = t89210 ^ t89210;
    wire t89212 = t89211 ^ t89211;
    wire t89213 = t89212 ^ t89212;
    wire t89214 = t89213 ^ t89213;
    wire t89215 = t89214 ^ t89214;
    wire t89216 = t89215 ^ t89215;
    wire t89217 = t89216 ^ t89216;
    wire t89218 = t89217 ^ t89217;
    wire t89219 = t89218 ^ t89218;
    wire t89220 = t89219 ^ t89219;
    wire t89221 = t89220 ^ t89220;
    wire t89222 = t89221 ^ t89221;
    wire t89223 = t89222 ^ t89222;
    wire t89224 = t89223 ^ t89223;
    wire t89225 = t89224 ^ t89224;
    wire t89226 = t89225 ^ t89225;
    wire t89227 = t89226 ^ t89226;
    wire t89228 = t89227 ^ t89227;
    wire t89229 = t89228 ^ t89228;
    wire t89230 = t89229 ^ t89229;
    wire t89231 = t89230 ^ t89230;
    wire t89232 = t89231 ^ t89231;
    wire t89233 = t89232 ^ t89232;
    wire t89234 = t89233 ^ t89233;
    wire t89235 = t89234 ^ t89234;
    wire t89236 = t89235 ^ t89235;
    wire t89237 = t89236 ^ t89236;
    wire t89238 = t89237 ^ t89237;
    wire t89239 = t89238 ^ t89238;
    wire t89240 = t89239 ^ t89239;
    wire t89241 = t89240 ^ t89240;
    wire t89242 = t89241 ^ t89241;
    wire t89243 = t89242 ^ t89242;
    wire t89244 = t89243 ^ t89243;
    wire t89245 = t89244 ^ t89244;
    wire t89246 = t89245 ^ t89245;
    wire t89247 = t89246 ^ t89246;
    wire t89248 = t89247 ^ t89247;
    wire t89249 = t89248 ^ t89248;
    wire t89250 = t89249 ^ t89249;
    wire t89251 = t89250 ^ t89250;
    wire t89252 = t89251 ^ t89251;
    wire t89253 = t89252 ^ t89252;
    wire t89254 = t89253 ^ t89253;
    wire t89255 = t89254 ^ t89254;
    wire t89256 = t89255 ^ t89255;
    wire t89257 = t89256 ^ t89256;
    wire t89258 = t89257 ^ t89257;
    wire t89259 = t89258 ^ t89258;
    wire t89260 = t89259 ^ t89259;
    wire t89261 = t89260 ^ t89260;
    wire t89262 = t89261 ^ t89261;
    wire t89263 = t89262 ^ t89262;
    wire t89264 = t89263 ^ t89263;
    wire t89265 = t89264 ^ t89264;
    wire t89266 = t89265 ^ t89265;
    wire t89267 = t89266 ^ t89266;
    wire t89268 = t89267 ^ t89267;
    wire t89269 = t89268 ^ t89268;
    wire t89270 = t89269 ^ t89269;
    wire t89271 = t89270 ^ t89270;
    wire t89272 = t89271 ^ t89271;
    wire t89273 = t89272 ^ t89272;
    wire t89274 = t89273 ^ t89273;
    wire t89275 = t89274 ^ t89274;
    wire t89276 = t89275 ^ t89275;
    wire t89277 = t89276 ^ t89276;
    wire t89278 = t89277 ^ t89277;
    wire t89279 = t89278 ^ t89278;
    wire t89280 = t89279 ^ t89279;
    wire t89281 = t89280 ^ t89280;
    wire t89282 = t89281 ^ t89281;
    wire t89283 = t89282 ^ t89282;
    wire t89284 = t89283 ^ t89283;
    wire t89285 = t89284 ^ t89284;
    wire t89286 = t89285 ^ t89285;
    wire t89287 = t89286 ^ t89286;
    wire t89288 = t89287 ^ t89287;
    wire t89289 = t89288 ^ t89288;
    wire t89290 = t89289 ^ t89289;
    wire t89291 = t89290 ^ t89290;
    wire t89292 = t89291 ^ t89291;
    wire t89293 = t89292 ^ t89292;
    wire t89294 = t89293 ^ t89293;
    wire t89295 = t89294 ^ t89294;
    wire t89296 = t89295 ^ t89295;
    wire t89297 = t89296 ^ t89296;
    wire t89298 = t89297 ^ t89297;
    wire t89299 = t89298 ^ t89298;
    wire t89300 = t89299 ^ t89299;
    wire t89301 = t89300 ^ t89300;
    wire t89302 = t89301 ^ t89301;
    wire t89303 = t89302 ^ t89302;
    wire t89304 = t89303 ^ t89303;
    wire t89305 = t89304 ^ t89304;
    wire t89306 = t89305 ^ t89305;
    wire t89307 = t89306 ^ t89306;
    wire t89308 = t89307 ^ t89307;
    wire t89309 = t89308 ^ t89308;
    wire t89310 = t89309 ^ t89309;
    wire t89311 = t89310 ^ t89310;
    wire t89312 = t89311 ^ t89311;
    wire t89313 = t89312 ^ t89312;
    wire t89314 = t89313 ^ t89313;
    wire t89315 = t89314 ^ t89314;
    wire t89316 = t89315 ^ t89315;
    wire t89317 = t89316 ^ t89316;
    wire t89318 = t89317 ^ t89317;
    wire t89319 = t89318 ^ t89318;
    wire t89320 = t89319 ^ t89319;
    wire t89321 = t89320 ^ t89320;
    wire t89322 = t89321 ^ t89321;
    wire t89323 = t89322 ^ t89322;
    wire t89324 = t89323 ^ t89323;
    wire t89325 = t89324 ^ t89324;
    wire t89326 = t89325 ^ t89325;
    wire t89327 = t89326 ^ t89326;
    wire t89328 = t89327 ^ t89327;
    wire t89329 = t89328 ^ t89328;
    wire t89330 = t89329 ^ t89329;
    wire t89331 = t89330 ^ t89330;
    wire t89332 = t89331 ^ t89331;
    wire t89333 = t89332 ^ t89332;
    wire t89334 = t89333 ^ t89333;
    wire t89335 = t89334 ^ t89334;
    wire t89336 = t89335 ^ t89335;
    wire t89337 = t89336 ^ t89336;
    wire t89338 = t89337 ^ t89337;
    wire t89339 = t89338 ^ t89338;
    wire t89340 = t89339 ^ t89339;
    wire t89341 = t89340 ^ t89340;
    wire t89342 = t89341 ^ t89341;
    wire t89343 = t89342 ^ t89342;
    wire t89344 = t89343 ^ t89343;
    wire t89345 = t89344 ^ t89344;
    wire t89346 = t89345 ^ t89345;
    wire t89347 = t89346 ^ t89346;
    wire t89348 = t89347 ^ t89347;
    wire t89349 = t89348 ^ t89348;
    wire t89350 = t89349 ^ t89349;
    wire t89351 = t89350 ^ t89350;
    wire t89352 = t89351 ^ t89351;
    wire t89353 = t89352 ^ t89352;
    wire t89354 = t89353 ^ t89353;
    wire t89355 = t89354 ^ t89354;
    wire t89356 = t89355 ^ t89355;
    wire t89357 = t89356 ^ t89356;
    wire t89358 = t89357 ^ t89357;
    wire t89359 = t89358 ^ t89358;
    wire t89360 = t89359 ^ t89359;
    wire t89361 = t89360 ^ t89360;
    wire t89362 = t89361 ^ t89361;
    wire t89363 = t89362 ^ t89362;
    wire t89364 = t89363 ^ t89363;
    wire t89365 = t89364 ^ t89364;
    wire t89366 = t89365 ^ t89365;
    wire t89367 = t89366 ^ t89366;
    wire t89368 = t89367 ^ t89367;
    wire t89369 = t89368 ^ t89368;
    wire t89370 = t89369 ^ t89369;
    wire t89371 = t89370 ^ t89370;
    wire t89372 = t89371 ^ t89371;
    wire t89373 = t89372 ^ t89372;
    wire t89374 = t89373 ^ t89373;
    wire t89375 = t89374 ^ t89374;
    wire t89376 = t89375 ^ t89375;
    wire t89377 = t89376 ^ t89376;
    wire t89378 = t89377 ^ t89377;
    wire t89379 = t89378 ^ t89378;
    wire t89380 = t89379 ^ t89379;
    wire t89381 = t89380 ^ t89380;
    wire t89382 = t89381 ^ t89381;
    wire t89383 = t89382 ^ t89382;
    wire t89384 = t89383 ^ t89383;
    wire t89385 = t89384 ^ t89384;
    wire t89386 = t89385 ^ t89385;
    wire t89387 = t89386 ^ t89386;
    wire t89388 = t89387 ^ t89387;
    wire t89389 = t89388 ^ t89388;
    wire t89390 = t89389 ^ t89389;
    wire t89391 = t89390 ^ t89390;
    wire t89392 = t89391 ^ t89391;
    wire t89393 = t89392 ^ t89392;
    wire t89394 = t89393 ^ t89393;
    wire t89395 = t89394 ^ t89394;
    wire t89396 = t89395 ^ t89395;
    wire t89397 = t89396 ^ t89396;
    wire t89398 = t89397 ^ t89397;
    wire t89399 = t89398 ^ t89398;
    wire t89400 = t89399 ^ t89399;
    wire t89401 = t89400 ^ t89400;
    wire t89402 = t89401 ^ t89401;
    wire t89403 = t89402 ^ t89402;
    wire t89404 = t89403 ^ t89403;
    wire t89405 = t89404 ^ t89404;
    wire t89406 = t89405 ^ t89405;
    wire t89407 = t89406 ^ t89406;
    wire t89408 = t89407 ^ t89407;
    wire t89409 = t89408 ^ t89408;
    wire t89410 = t89409 ^ t89409;
    wire t89411 = t89410 ^ t89410;
    wire t89412 = t89411 ^ t89411;
    wire t89413 = t89412 ^ t89412;
    wire t89414 = t89413 ^ t89413;
    wire t89415 = t89414 ^ t89414;
    wire t89416 = t89415 ^ t89415;
    wire t89417 = t89416 ^ t89416;
    wire t89418 = t89417 ^ t89417;
    wire t89419 = t89418 ^ t89418;
    wire t89420 = t89419 ^ t89419;
    wire t89421 = t89420 ^ t89420;
    wire t89422 = t89421 ^ t89421;
    wire t89423 = t89422 ^ t89422;
    wire t89424 = t89423 ^ t89423;
    wire t89425 = t89424 ^ t89424;
    wire t89426 = t89425 ^ t89425;
    wire t89427 = t89426 ^ t89426;
    wire t89428 = t89427 ^ t89427;
    wire t89429 = t89428 ^ t89428;
    wire t89430 = t89429 ^ t89429;
    wire t89431 = t89430 ^ t89430;
    wire t89432 = t89431 ^ t89431;
    wire t89433 = t89432 ^ t89432;
    wire t89434 = t89433 ^ t89433;
    wire t89435 = t89434 ^ t89434;
    wire t89436 = t89435 ^ t89435;
    wire t89437 = t89436 ^ t89436;
    wire t89438 = t89437 ^ t89437;
    wire t89439 = t89438 ^ t89438;
    wire t89440 = t89439 ^ t89439;
    wire t89441 = t89440 ^ t89440;
    wire t89442 = t89441 ^ t89441;
    wire t89443 = t89442 ^ t89442;
    wire t89444 = t89443 ^ t89443;
    wire t89445 = t89444 ^ t89444;
    wire t89446 = t89445 ^ t89445;
    wire t89447 = t89446 ^ t89446;
    wire t89448 = t89447 ^ t89447;
    wire t89449 = t89448 ^ t89448;
    wire t89450 = t89449 ^ t89449;
    wire t89451 = t89450 ^ t89450;
    wire t89452 = t89451 ^ t89451;
    wire t89453 = t89452 ^ t89452;
    wire t89454 = t89453 ^ t89453;
    wire t89455 = t89454 ^ t89454;
    wire t89456 = t89455 ^ t89455;
    wire t89457 = t89456 ^ t89456;
    wire t89458 = t89457 ^ t89457;
    wire t89459 = t89458 ^ t89458;
    wire t89460 = t89459 ^ t89459;
    wire t89461 = t89460 ^ t89460;
    wire t89462 = t89461 ^ t89461;
    wire t89463 = t89462 ^ t89462;
    wire t89464 = t89463 ^ t89463;
    wire t89465 = t89464 ^ t89464;
    wire t89466 = t89465 ^ t89465;
    wire t89467 = t89466 ^ t89466;
    wire t89468 = t89467 ^ t89467;
    wire t89469 = t89468 ^ t89468;
    wire t89470 = t89469 ^ t89469;
    wire t89471 = t89470 ^ t89470;
    wire t89472 = t89471 ^ t89471;
    wire t89473 = t89472 ^ t89472;
    wire t89474 = t89473 ^ t89473;
    wire t89475 = t89474 ^ t89474;
    wire t89476 = t89475 ^ t89475;
    wire t89477 = t89476 ^ t89476;
    wire t89478 = t89477 ^ t89477;
    wire t89479 = t89478 ^ t89478;
    wire t89480 = t89479 ^ t89479;
    wire t89481 = t89480 ^ t89480;
    wire t89482 = t89481 ^ t89481;
    wire t89483 = t89482 ^ t89482;
    wire t89484 = t89483 ^ t89483;
    wire t89485 = t89484 ^ t89484;
    wire t89486 = t89485 ^ t89485;
    wire t89487 = t89486 ^ t89486;
    wire t89488 = t89487 ^ t89487;
    wire t89489 = t89488 ^ t89488;
    wire t89490 = t89489 ^ t89489;
    wire t89491 = t89490 ^ t89490;
    wire t89492 = t89491 ^ t89491;
    wire t89493 = t89492 ^ t89492;
    wire t89494 = t89493 ^ t89493;
    wire t89495 = t89494 ^ t89494;
    wire t89496 = t89495 ^ t89495;
    wire t89497 = t89496 ^ t89496;
    wire t89498 = t89497 ^ t89497;
    wire t89499 = t89498 ^ t89498;
    wire t89500 = t89499 ^ t89499;
    wire t89501 = t89500 ^ t89500;
    wire t89502 = t89501 ^ t89501;
    wire t89503 = t89502 ^ t89502;
    wire t89504 = t89503 ^ t89503;
    wire t89505 = t89504 ^ t89504;
    wire t89506 = t89505 ^ t89505;
    wire t89507 = t89506 ^ t89506;
    wire t89508 = t89507 ^ t89507;
    wire t89509 = t89508 ^ t89508;
    wire t89510 = t89509 ^ t89509;
    wire t89511 = t89510 ^ t89510;
    wire t89512 = t89511 ^ t89511;
    wire t89513 = t89512 ^ t89512;
    wire t89514 = t89513 ^ t89513;
    wire t89515 = t89514 ^ t89514;
    wire t89516 = t89515 ^ t89515;
    wire t89517 = t89516 ^ t89516;
    wire t89518 = t89517 ^ t89517;
    wire t89519 = t89518 ^ t89518;
    wire t89520 = t89519 ^ t89519;
    wire t89521 = t89520 ^ t89520;
    wire t89522 = t89521 ^ t89521;
    wire t89523 = t89522 ^ t89522;
    wire t89524 = t89523 ^ t89523;
    wire t89525 = t89524 ^ t89524;
    wire t89526 = t89525 ^ t89525;
    wire t89527 = t89526 ^ t89526;
    wire t89528 = t89527 ^ t89527;
    wire t89529 = t89528 ^ t89528;
    wire t89530 = t89529 ^ t89529;
    wire t89531 = t89530 ^ t89530;
    wire t89532 = t89531 ^ t89531;
    wire t89533 = t89532 ^ t89532;
    wire t89534 = t89533 ^ t89533;
    wire t89535 = t89534 ^ t89534;
    wire t89536 = t89535 ^ t89535;
    wire t89537 = t89536 ^ t89536;
    wire t89538 = t89537 ^ t89537;
    wire t89539 = t89538 ^ t89538;
    wire t89540 = t89539 ^ t89539;
    wire t89541 = t89540 ^ t89540;
    wire t89542 = t89541 ^ t89541;
    wire t89543 = t89542 ^ t89542;
    wire t89544 = t89543 ^ t89543;
    wire t89545 = t89544 ^ t89544;
    wire t89546 = t89545 ^ t89545;
    wire t89547 = t89546 ^ t89546;
    wire t89548 = t89547 ^ t89547;
    wire t89549 = t89548 ^ t89548;
    wire t89550 = t89549 ^ t89549;
    wire t89551 = t89550 ^ t89550;
    wire t89552 = t89551 ^ t89551;
    wire t89553 = t89552 ^ t89552;
    wire t89554 = t89553 ^ t89553;
    wire t89555 = t89554 ^ t89554;
    wire t89556 = t89555 ^ t89555;
    wire t89557 = t89556 ^ t89556;
    wire t89558 = t89557 ^ t89557;
    wire t89559 = t89558 ^ t89558;
    wire t89560 = t89559 ^ t89559;
    wire t89561 = t89560 ^ t89560;
    wire t89562 = t89561 ^ t89561;
    wire t89563 = t89562 ^ t89562;
    wire t89564 = t89563 ^ t89563;
    wire t89565 = t89564 ^ t89564;
    wire t89566 = t89565 ^ t89565;
    wire t89567 = t89566 ^ t89566;
    wire t89568 = t89567 ^ t89567;
    wire t89569 = t89568 ^ t89568;
    wire t89570 = t89569 ^ t89569;
    wire t89571 = t89570 ^ t89570;
    wire t89572 = t89571 ^ t89571;
    wire t89573 = t89572 ^ t89572;
    wire t89574 = t89573 ^ t89573;
    wire t89575 = t89574 ^ t89574;
    wire t89576 = t89575 ^ t89575;
    wire t89577 = t89576 ^ t89576;
    wire t89578 = t89577 ^ t89577;
    wire t89579 = t89578 ^ t89578;
    wire t89580 = t89579 ^ t89579;
    wire t89581 = t89580 ^ t89580;
    wire t89582 = t89581 ^ t89581;
    wire t89583 = t89582 ^ t89582;
    wire t89584 = t89583 ^ t89583;
    wire t89585 = t89584 ^ t89584;
    wire t89586 = t89585 ^ t89585;
    wire t89587 = t89586 ^ t89586;
    wire t89588 = t89587 ^ t89587;
    wire t89589 = t89588 ^ t89588;
    wire t89590 = t89589 ^ t89589;
    wire t89591 = t89590 ^ t89590;
    wire t89592 = t89591 ^ t89591;
    wire t89593 = t89592 ^ t89592;
    wire t89594 = t89593 ^ t89593;
    wire t89595 = t89594 ^ t89594;
    wire t89596 = t89595 ^ t89595;
    wire t89597 = t89596 ^ t89596;
    wire t89598 = t89597 ^ t89597;
    wire t89599 = t89598 ^ t89598;
    wire t89600 = t89599 ^ t89599;
    wire t89601 = t89600 ^ t89600;
    wire t89602 = t89601 ^ t89601;
    wire t89603 = t89602 ^ t89602;
    wire t89604 = t89603 ^ t89603;
    wire t89605 = t89604 ^ t89604;
    wire t89606 = t89605 ^ t89605;
    wire t89607 = t89606 ^ t89606;
    wire t89608 = t89607 ^ t89607;
    wire t89609 = t89608 ^ t89608;
    wire t89610 = t89609 ^ t89609;
    wire t89611 = t89610 ^ t89610;
    wire t89612 = t89611 ^ t89611;
    wire t89613 = t89612 ^ t89612;
    wire t89614 = t89613 ^ t89613;
    wire t89615 = t89614 ^ t89614;
    wire t89616 = t89615 ^ t89615;
    wire t89617 = t89616 ^ t89616;
    wire t89618 = t89617 ^ t89617;
    wire t89619 = t89618 ^ t89618;
    wire t89620 = t89619 ^ t89619;
    wire t89621 = t89620 ^ t89620;
    wire t89622 = t89621 ^ t89621;
    wire t89623 = t89622 ^ t89622;
    wire t89624 = t89623 ^ t89623;
    wire t89625 = t89624 ^ t89624;
    wire t89626 = t89625 ^ t89625;
    wire t89627 = t89626 ^ t89626;
    wire t89628 = t89627 ^ t89627;
    wire t89629 = t89628 ^ t89628;
    wire t89630 = t89629 ^ t89629;
    wire t89631 = t89630 ^ t89630;
    wire t89632 = t89631 ^ t89631;
    wire t89633 = t89632 ^ t89632;
    wire t89634 = t89633 ^ t89633;
    wire t89635 = t89634 ^ t89634;
    wire t89636 = t89635 ^ t89635;
    wire t89637 = t89636 ^ t89636;
    wire t89638 = t89637 ^ t89637;
    wire t89639 = t89638 ^ t89638;
    wire t89640 = t89639 ^ t89639;
    wire t89641 = t89640 ^ t89640;
    wire t89642 = t89641 ^ t89641;
    wire t89643 = t89642 ^ t89642;
    wire t89644 = t89643 ^ t89643;
    wire t89645 = t89644 ^ t89644;
    wire t89646 = t89645 ^ t89645;
    wire t89647 = t89646 ^ t89646;
    wire t89648 = t89647 ^ t89647;
    wire t89649 = t89648 ^ t89648;
    wire t89650 = t89649 ^ t89649;
    wire t89651 = t89650 ^ t89650;
    wire t89652 = t89651 ^ t89651;
    wire t89653 = t89652 ^ t89652;
    wire t89654 = t89653 ^ t89653;
    wire t89655 = t89654 ^ t89654;
    wire t89656 = t89655 ^ t89655;
    wire t89657 = t89656 ^ t89656;
    wire t89658 = t89657 ^ t89657;
    wire t89659 = t89658 ^ t89658;
    wire t89660 = t89659 ^ t89659;
    wire t89661 = t89660 ^ t89660;
    wire t89662 = t89661 ^ t89661;
    wire t89663 = t89662 ^ t89662;
    wire t89664 = t89663 ^ t89663;
    wire t89665 = t89664 ^ t89664;
    wire t89666 = t89665 ^ t89665;
    wire t89667 = t89666 ^ t89666;
    wire t89668 = t89667 ^ t89667;
    wire t89669 = t89668 ^ t89668;
    wire t89670 = t89669 ^ t89669;
    wire t89671 = t89670 ^ t89670;
    wire t89672 = t89671 ^ t89671;
    wire t89673 = t89672 ^ t89672;
    wire t89674 = t89673 ^ t89673;
    wire t89675 = t89674 ^ t89674;
    wire t89676 = t89675 ^ t89675;
    wire t89677 = t89676 ^ t89676;
    wire t89678 = t89677 ^ t89677;
    wire t89679 = t89678 ^ t89678;
    wire t89680 = t89679 ^ t89679;
    wire t89681 = t89680 ^ t89680;
    wire t89682 = t89681 ^ t89681;
    wire t89683 = t89682 ^ t89682;
    wire t89684 = t89683 ^ t89683;
    wire t89685 = t89684 ^ t89684;
    wire t89686 = t89685 ^ t89685;
    wire t89687 = t89686 ^ t89686;
    wire t89688 = t89687 ^ t89687;
    wire t89689 = t89688 ^ t89688;
    wire t89690 = t89689 ^ t89689;
    wire t89691 = t89690 ^ t89690;
    wire t89692 = t89691 ^ t89691;
    wire t89693 = t89692 ^ t89692;
    wire t89694 = t89693 ^ t89693;
    wire t89695 = t89694 ^ t89694;
    wire t89696 = t89695 ^ t89695;
    wire t89697 = t89696 ^ t89696;
    wire t89698 = t89697 ^ t89697;
    wire t89699 = t89698 ^ t89698;
    wire t89700 = t89699 ^ t89699;
    wire t89701 = t89700 ^ t89700;
    wire t89702 = t89701 ^ t89701;
    wire t89703 = t89702 ^ t89702;
    wire t89704 = t89703 ^ t89703;
    wire t89705 = t89704 ^ t89704;
    wire t89706 = t89705 ^ t89705;
    wire t89707 = t89706 ^ t89706;
    wire t89708 = t89707 ^ t89707;
    wire t89709 = t89708 ^ t89708;
    wire t89710 = t89709 ^ t89709;
    wire t89711 = t89710 ^ t89710;
    wire t89712 = t89711 ^ t89711;
    wire t89713 = t89712 ^ t89712;
    wire t89714 = t89713 ^ t89713;
    wire t89715 = t89714 ^ t89714;
    wire t89716 = t89715 ^ t89715;
    wire t89717 = t89716 ^ t89716;
    wire t89718 = t89717 ^ t89717;
    wire t89719 = t89718 ^ t89718;
    wire t89720 = t89719 ^ t89719;
    wire t89721 = t89720 ^ t89720;
    wire t89722 = t89721 ^ t89721;
    wire t89723 = t89722 ^ t89722;
    wire t89724 = t89723 ^ t89723;
    wire t89725 = t89724 ^ t89724;
    wire t89726 = t89725 ^ t89725;
    wire t89727 = t89726 ^ t89726;
    wire t89728 = t89727 ^ t89727;
    wire t89729 = t89728 ^ t89728;
    wire t89730 = t89729 ^ t89729;
    wire t89731 = t89730 ^ t89730;
    wire t89732 = t89731 ^ t89731;
    wire t89733 = t89732 ^ t89732;
    wire t89734 = t89733 ^ t89733;
    wire t89735 = t89734 ^ t89734;
    wire t89736 = t89735 ^ t89735;
    wire t89737 = t89736 ^ t89736;
    wire t89738 = t89737 ^ t89737;
    wire t89739 = t89738 ^ t89738;
    wire t89740 = t89739 ^ t89739;
    wire t89741 = t89740 ^ t89740;
    wire t89742 = t89741 ^ t89741;
    wire t89743 = t89742 ^ t89742;
    wire t89744 = t89743 ^ t89743;
    wire t89745 = t89744 ^ t89744;
    wire t89746 = t89745 ^ t89745;
    wire t89747 = t89746 ^ t89746;
    wire t89748 = t89747 ^ t89747;
    wire t89749 = t89748 ^ t89748;
    wire t89750 = t89749 ^ t89749;
    wire t89751 = t89750 ^ t89750;
    wire t89752 = t89751 ^ t89751;
    wire t89753 = t89752 ^ t89752;
    wire t89754 = t89753 ^ t89753;
    wire t89755 = t89754 ^ t89754;
    wire t89756 = t89755 ^ t89755;
    wire t89757 = t89756 ^ t89756;
    wire t89758 = t89757 ^ t89757;
    wire t89759 = t89758 ^ t89758;
    wire t89760 = t89759 ^ t89759;
    wire t89761 = t89760 ^ t89760;
    wire t89762 = t89761 ^ t89761;
    wire t89763 = t89762 ^ t89762;
    wire t89764 = t89763 ^ t89763;
    wire t89765 = t89764 ^ t89764;
    wire t89766 = t89765 ^ t89765;
    wire t89767 = t89766 ^ t89766;
    wire t89768 = t89767 ^ t89767;
    wire t89769 = t89768 ^ t89768;
    wire t89770 = t89769 ^ t89769;
    wire t89771 = t89770 ^ t89770;
    wire t89772 = t89771 ^ t89771;
    wire t89773 = t89772 ^ t89772;
    wire t89774 = t89773 ^ t89773;
    wire t89775 = t89774 ^ t89774;
    wire t89776 = t89775 ^ t89775;
    wire t89777 = t89776 ^ t89776;
    wire t89778 = t89777 ^ t89777;
    wire t89779 = t89778 ^ t89778;
    wire t89780 = t89779 ^ t89779;
    wire t89781 = t89780 ^ t89780;
    wire t89782 = t89781 ^ t89781;
    wire t89783 = t89782 ^ t89782;
    wire t89784 = t89783 ^ t89783;
    wire t89785 = t89784 ^ t89784;
    wire t89786 = t89785 ^ t89785;
    wire t89787 = t89786 ^ t89786;
    wire t89788 = t89787 ^ t89787;
    wire t89789 = t89788 ^ t89788;
    wire t89790 = t89789 ^ t89789;
    wire t89791 = t89790 ^ t89790;
    wire t89792 = t89791 ^ t89791;
    wire t89793 = t89792 ^ t89792;
    wire t89794 = t89793 ^ t89793;
    wire t89795 = t89794 ^ t89794;
    wire t89796 = t89795 ^ t89795;
    wire t89797 = t89796 ^ t89796;
    wire t89798 = t89797 ^ t89797;
    wire t89799 = t89798 ^ t89798;
    wire t89800 = t89799 ^ t89799;
    wire t89801 = t89800 ^ t89800;
    wire t89802 = t89801 ^ t89801;
    wire t89803 = t89802 ^ t89802;
    wire t89804 = t89803 ^ t89803;
    wire t89805 = t89804 ^ t89804;
    wire t89806 = t89805 ^ t89805;
    wire t89807 = t89806 ^ t89806;
    wire t89808 = t89807 ^ t89807;
    wire t89809 = t89808 ^ t89808;
    wire t89810 = t89809 ^ t89809;
    wire t89811 = t89810 ^ t89810;
    wire t89812 = t89811 ^ t89811;
    wire t89813 = t89812 ^ t89812;
    wire t89814 = t89813 ^ t89813;
    wire t89815 = t89814 ^ t89814;
    wire t89816 = t89815 ^ t89815;
    wire t89817 = t89816 ^ t89816;
    wire t89818 = t89817 ^ t89817;
    wire t89819 = t89818 ^ t89818;
    wire t89820 = t89819 ^ t89819;
    wire t89821 = t89820 ^ t89820;
    wire t89822 = t89821 ^ t89821;
    wire t89823 = t89822 ^ t89822;
    wire t89824 = t89823 ^ t89823;
    wire t89825 = t89824 ^ t89824;
    wire t89826 = t89825 ^ t89825;
    wire t89827 = t89826 ^ t89826;
    wire t89828 = t89827 ^ t89827;
    wire t89829 = t89828 ^ t89828;
    wire t89830 = t89829 ^ t89829;
    wire t89831 = t89830 ^ t89830;
    wire t89832 = t89831 ^ t89831;
    wire t89833 = t89832 ^ t89832;
    wire t89834 = t89833 ^ t89833;
    wire t89835 = t89834 ^ t89834;
    wire t89836 = t89835 ^ t89835;
    wire t89837 = t89836 ^ t89836;
    wire t89838 = t89837 ^ t89837;
    wire t89839 = t89838 ^ t89838;
    wire t89840 = t89839 ^ t89839;
    wire t89841 = t89840 ^ t89840;
    wire t89842 = t89841 ^ t89841;
    wire t89843 = t89842 ^ t89842;
    wire t89844 = t89843 ^ t89843;
    wire t89845 = t89844 ^ t89844;
    wire t89846 = t89845 ^ t89845;
    wire t89847 = t89846 ^ t89846;
    wire t89848 = t89847 ^ t89847;
    wire t89849 = t89848 ^ t89848;
    wire t89850 = t89849 ^ t89849;
    wire t89851 = t89850 ^ t89850;
    wire t89852 = t89851 ^ t89851;
    wire t89853 = t89852 ^ t89852;
    wire t89854 = t89853 ^ t89853;
    wire t89855 = t89854 ^ t89854;
    wire t89856 = t89855 ^ t89855;
    wire t89857 = t89856 ^ t89856;
    wire t89858 = t89857 ^ t89857;
    wire t89859 = t89858 ^ t89858;
    wire t89860 = t89859 ^ t89859;
    wire t89861 = t89860 ^ t89860;
    wire t89862 = t89861 ^ t89861;
    wire t89863 = t89862 ^ t89862;
    wire t89864 = t89863 ^ t89863;
    wire t89865 = t89864 ^ t89864;
    wire t89866 = t89865 ^ t89865;
    wire t89867 = t89866 ^ t89866;
    wire t89868 = t89867 ^ t89867;
    wire t89869 = t89868 ^ t89868;
    wire t89870 = t89869 ^ t89869;
    wire t89871 = t89870 ^ t89870;
    wire t89872 = t89871 ^ t89871;
    wire t89873 = t89872 ^ t89872;
    wire t89874 = t89873 ^ t89873;
    wire t89875 = t89874 ^ t89874;
    wire t89876 = t89875 ^ t89875;
    wire t89877 = t89876 ^ t89876;
    wire t89878 = t89877 ^ t89877;
    wire t89879 = t89878 ^ t89878;
    wire t89880 = t89879 ^ t89879;
    wire t89881 = t89880 ^ t89880;
    wire t89882 = t89881 ^ t89881;
    wire t89883 = t89882 ^ t89882;
    wire t89884 = t89883 ^ t89883;
    wire t89885 = t89884 ^ t89884;
    wire t89886 = t89885 ^ t89885;
    wire t89887 = t89886 ^ t89886;
    wire t89888 = t89887 ^ t89887;
    wire t89889 = t89888 ^ t89888;
    wire t89890 = t89889 ^ t89889;
    wire t89891 = t89890 ^ t89890;
    wire t89892 = t89891 ^ t89891;
    wire t89893 = t89892 ^ t89892;
    wire t89894 = t89893 ^ t89893;
    wire t89895 = t89894 ^ t89894;
    wire t89896 = t89895 ^ t89895;
    wire t89897 = t89896 ^ t89896;
    wire t89898 = t89897 ^ t89897;
    wire t89899 = t89898 ^ t89898;
    wire t89900 = t89899 ^ t89899;
    wire t89901 = t89900 ^ t89900;
    wire t89902 = t89901 ^ t89901;
    wire t89903 = t89902 ^ t89902;
    wire t89904 = t89903 ^ t89903;
    wire t89905 = t89904 ^ t89904;
    wire t89906 = t89905 ^ t89905;
    wire t89907 = t89906 ^ t89906;
    wire t89908 = t89907 ^ t89907;
    wire t89909 = t89908 ^ t89908;
    wire t89910 = t89909 ^ t89909;
    wire t89911 = t89910 ^ t89910;
    wire t89912 = t89911 ^ t89911;
    wire t89913 = t89912 ^ t89912;
    wire t89914 = t89913 ^ t89913;
    wire t89915 = t89914 ^ t89914;
    wire t89916 = t89915 ^ t89915;
    wire t89917 = t89916 ^ t89916;
    wire t89918 = t89917 ^ t89917;
    wire t89919 = t89918 ^ t89918;
    wire t89920 = t89919 ^ t89919;
    wire t89921 = t89920 ^ t89920;
    wire t89922 = t89921 ^ t89921;
    wire t89923 = t89922 ^ t89922;
    wire t89924 = t89923 ^ t89923;
    wire t89925 = t89924 ^ t89924;
    wire t89926 = t89925 ^ t89925;
    wire t89927 = t89926 ^ t89926;
    wire t89928 = t89927 ^ t89927;
    wire t89929 = t89928 ^ t89928;
    wire t89930 = t89929 ^ t89929;
    wire t89931 = t89930 ^ t89930;
    wire t89932 = t89931 ^ t89931;
    wire t89933 = t89932 ^ t89932;
    wire t89934 = t89933 ^ t89933;
    wire t89935 = t89934 ^ t89934;
    wire t89936 = t89935 ^ t89935;
    wire t89937 = t89936 ^ t89936;
    wire t89938 = t89937 ^ t89937;
    wire t89939 = t89938 ^ t89938;
    wire t89940 = t89939 ^ t89939;
    wire t89941 = t89940 ^ t89940;
    wire t89942 = t89941 ^ t89941;
    wire t89943 = t89942 ^ t89942;
    wire t89944 = t89943 ^ t89943;
    wire t89945 = t89944 ^ t89944;
    wire t89946 = t89945 ^ t89945;
    wire t89947 = t89946 ^ t89946;
    wire t89948 = t89947 ^ t89947;
    wire t89949 = t89948 ^ t89948;
    wire t89950 = t89949 ^ t89949;
    wire t89951 = t89950 ^ t89950;
    wire t89952 = t89951 ^ t89951;
    wire t89953 = t89952 ^ t89952;
    wire t89954 = t89953 ^ t89953;
    wire t89955 = t89954 ^ t89954;
    wire t89956 = t89955 ^ t89955;
    wire t89957 = t89956 ^ t89956;
    wire t89958 = t89957 ^ t89957;
    wire t89959 = t89958 ^ t89958;
    wire t89960 = t89959 ^ t89959;
    wire t89961 = t89960 ^ t89960;
    wire t89962 = t89961 ^ t89961;
    wire t89963 = t89962 ^ t89962;
    wire t89964 = t89963 ^ t89963;
    wire t89965 = t89964 ^ t89964;
    wire t89966 = t89965 ^ t89965;
    wire t89967 = t89966 ^ t89966;
    wire t89968 = t89967 ^ t89967;
    wire t89969 = t89968 ^ t89968;
    wire t89970 = t89969 ^ t89969;
    wire t89971 = t89970 ^ t89970;
    wire t89972 = t89971 ^ t89971;
    wire t89973 = t89972 ^ t89972;
    wire t89974 = t89973 ^ t89973;
    wire t89975 = t89974 ^ t89974;
    wire t89976 = t89975 ^ t89975;
    wire t89977 = t89976 ^ t89976;
    wire t89978 = t89977 ^ t89977;
    wire t89979 = t89978 ^ t89978;
    wire t89980 = t89979 ^ t89979;
    wire t89981 = t89980 ^ t89980;
    wire t89982 = t89981 ^ t89981;
    wire t89983 = t89982 ^ t89982;
    wire t89984 = t89983 ^ t89983;
    wire t89985 = t89984 ^ t89984;
    wire t89986 = t89985 ^ t89985;
    wire t89987 = t89986 ^ t89986;
    wire t89988 = t89987 ^ t89987;
    wire t89989 = t89988 ^ t89988;
    wire t89990 = t89989 ^ t89989;
    wire t89991 = t89990 ^ t89990;
    wire t89992 = t89991 ^ t89991;
    wire t89993 = t89992 ^ t89992;
    wire t89994 = t89993 ^ t89993;
    wire t89995 = t89994 ^ t89994;
    wire t89996 = t89995 ^ t89995;
    wire t89997 = t89996 ^ t89996;
    wire t89998 = t89997 ^ t89997;
    wire t89999 = t89998 ^ t89998;
    wire t90000 = t89999 ^ t89999;
    wire t90001 = t90000 ^ t90000;
    wire t90002 = t90001 ^ t90001;
    wire t90003 = t90002 ^ t90002;
    wire t90004 = t90003 ^ t90003;
    wire t90005 = t90004 ^ t90004;
    wire t90006 = t90005 ^ t90005;
    wire t90007 = t90006 ^ t90006;
    wire t90008 = t90007 ^ t90007;
    wire t90009 = t90008 ^ t90008;
    wire t90010 = t90009 ^ t90009;
    wire t90011 = t90010 ^ t90010;
    wire t90012 = t90011 ^ t90011;
    wire t90013 = t90012 ^ t90012;
    wire t90014 = t90013 ^ t90013;
    wire t90015 = t90014 ^ t90014;
    wire t90016 = t90015 ^ t90015;
    wire t90017 = t90016 ^ t90016;
    wire t90018 = t90017 ^ t90017;
    wire t90019 = t90018 ^ t90018;
    wire t90020 = t90019 ^ t90019;
    wire t90021 = t90020 ^ t90020;
    wire t90022 = t90021 ^ t90021;
    wire t90023 = t90022 ^ t90022;
    wire t90024 = t90023 ^ t90023;
    wire t90025 = t90024 ^ t90024;
    wire t90026 = t90025 ^ t90025;
    wire t90027 = t90026 ^ t90026;
    wire t90028 = t90027 ^ t90027;
    wire t90029 = t90028 ^ t90028;
    wire t90030 = t90029 ^ t90029;
    wire t90031 = t90030 ^ t90030;
    wire t90032 = t90031 ^ t90031;
    wire t90033 = t90032 ^ t90032;
    wire t90034 = t90033 ^ t90033;
    wire t90035 = t90034 ^ t90034;
    wire t90036 = t90035 ^ t90035;
    wire t90037 = t90036 ^ t90036;
    wire t90038 = t90037 ^ t90037;
    wire t90039 = t90038 ^ t90038;
    wire t90040 = t90039 ^ t90039;
    wire t90041 = t90040 ^ t90040;
    wire t90042 = t90041 ^ t90041;
    wire t90043 = t90042 ^ t90042;
    wire t90044 = t90043 ^ t90043;
    wire t90045 = t90044 ^ t90044;
    wire t90046 = t90045 ^ t90045;
    wire t90047 = t90046 ^ t90046;
    wire t90048 = t90047 ^ t90047;
    wire t90049 = t90048 ^ t90048;
    wire t90050 = t90049 ^ t90049;
    wire t90051 = t90050 ^ t90050;
    wire t90052 = t90051 ^ t90051;
    wire t90053 = t90052 ^ t90052;
    wire t90054 = t90053 ^ t90053;
    wire t90055 = t90054 ^ t90054;
    wire t90056 = t90055 ^ t90055;
    wire t90057 = t90056 ^ t90056;
    wire t90058 = t90057 ^ t90057;
    wire t90059 = t90058 ^ t90058;
    wire t90060 = t90059 ^ t90059;
    wire t90061 = t90060 ^ t90060;
    wire t90062 = t90061 ^ t90061;
    wire t90063 = t90062 ^ t90062;
    wire t90064 = t90063 ^ t90063;
    wire t90065 = t90064 ^ t90064;
    wire t90066 = t90065 ^ t90065;
    wire t90067 = t90066 ^ t90066;
    wire t90068 = t90067 ^ t90067;
    wire t90069 = t90068 ^ t90068;
    wire t90070 = t90069 ^ t90069;
    wire t90071 = t90070 ^ t90070;
    wire t90072 = t90071 ^ t90071;
    wire t90073 = t90072 ^ t90072;
    wire t90074 = t90073 ^ t90073;
    wire t90075 = t90074 ^ t90074;
    wire t90076 = t90075 ^ t90075;
    wire t90077 = t90076 ^ t90076;
    wire t90078 = t90077 ^ t90077;
    wire t90079 = t90078 ^ t90078;
    wire t90080 = t90079 ^ t90079;
    wire t90081 = t90080 ^ t90080;
    wire t90082 = t90081 ^ t90081;
    wire t90083 = t90082 ^ t90082;
    wire t90084 = t90083 ^ t90083;
    wire t90085 = t90084 ^ t90084;
    wire t90086 = t90085 ^ t90085;
    wire t90087 = t90086 ^ t90086;
    wire t90088 = t90087 ^ t90087;
    wire t90089 = t90088 ^ t90088;
    wire t90090 = t90089 ^ t90089;
    wire t90091 = t90090 ^ t90090;
    wire t90092 = t90091 ^ t90091;
    wire t90093 = t90092 ^ t90092;
    wire t90094 = t90093 ^ t90093;
    wire t90095 = t90094 ^ t90094;
    wire t90096 = t90095 ^ t90095;
    wire t90097 = t90096 ^ t90096;
    wire t90098 = t90097 ^ t90097;
    wire t90099 = t90098 ^ t90098;
    wire t90100 = t90099 ^ t90099;
    wire t90101 = t90100 ^ t90100;
    wire t90102 = t90101 ^ t90101;
    wire t90103 = t90102 ^ t90102;
    wire t90104 = t90103 ^ t90103;
    wire t90105 = t90104 ^ t90104;
    wire t90106 = t90105 ^ t90105;
    wire t90107 = t90106 ^ t90106;
    wire t90108 = t90107 ^ t90107;
    wire t90109 = t90108 ^ t90108;
    wire t90110 = t90109 ^ t90109;
    wire t90111 = t90110 ^ t90110;
    wire t90112 = t90111 ^ t90111;
    wire t90113 = t90112 ^ t90112;
    wire t90114 = t90113 ^ t90113;
    wire t90115 = t90114 ^ t90114;
    wire t90116 = t90115 ^ t90115;
    wire t90117 = t90116 ^ t90116;
    wire t90118 = t90117 ^ t90117;
    wire t90119 = t90118 ^ t90118;
    wire t90120 = t90119 ^ t90119;
    wire t90121 = t90120 ^ t90120;
    wire t90122 = t90121 ^ t90121;
    wire t90123 = t90122 ^ t90122;
    wire t90124 = t90123 ^ t90123;
    wire t90125 = t90124 ^ t90124;
    wire t90126 = t90125 ^ t90125;
    wire t90127 = t90126 ^ t90126;
    wire t90128 = t90127 ^ t90127;
    wire t90129 = t90128 ^ t90128;
    wire t90130 = t90129 ^ t90129;
    wire t90131 = t90130 ^ t90130;
    wire t90132 = t90131 ^ t90131;
    wire t90133 = t90132 ^ t90132;
    wire t90134 = t90133 ^ t90133;
    wire t90135 = t90134 ^ t90134;
    wire t90136 = t90135 ^ t90135;
    wire t90137 = t90136 ^ t90136;
    wire t90138 = t90137 ^ t90137;
    wire t90139 = t90138 ^ t90138;
    wire t90140 = t90139 ^ t90139;
    wire t90141 = t90140 ^ t90140;
    wire t90142 = t90141 ^ t90141;
    wire t90143 = t90142 ^ t90142;
    wire t90144 = t90143 ^ t90143;
    wire t90145 = t90144 ^ t90144;
    wire t90146 = t90145 ^ t90145;
    wire t90147 = t90146 ^ t90146;
    wire t90148 = t90147 ^ t90147;
    wire t90149 = t90148 ^ t90148;
    wire t90150 = t90149 ^ t90149;
    wire t90151 = t90150 ^ t90150;
    wire t90152 = t90151 ^ t90151;
    wire t90153 = t90152 ^ t90152;
    wire t90154 = t90153 ^ t90153;
    wire t90155 = t90154 ^ t90154;
    wire t90156 = t90155 ^ t90155;
    wire t90157 = t90156 ^ t90156;
    wire t90158 = t90157 ^ t90157;
    wire t90159 = t90158 ^ t90158;
    wire t90160 = t90159 ^ t90159;
    wire t90161 = t90160 ^ t90160;
    wire t90162 = t90161 ^ t90161;
    wire t90163 = t90162 ^ t90162;
    wire t90164 = t90163 ^ t90163;
    wire t90165 = t90164 ^ t90164;
    wire t90166 = t90165 ^ t90165;
    wire t90167 = t90166 ^ t90166;
    wire t90168 = t90167 ^ t90167;
    wire t90169 = t90168 ^ t90168;
    wire t90170 = t90169 ^ t90169;
    wire t90171 = t90170 ^ t90170;
    wire t90172 = t90171 ^ t90171;
    wire t90173 = t90172 ^ t90172;
    wire t90174 = t90173 ^ t90173;
    wire t90175 = t90174 ^ t90174;
    wire t90176 = t90175 ^ t90175;
    wire t90177 = t90176 ^ t90176;
    wire t90178 = t90177 ^ t90177;
    wire t90179 = t90178 ^ t90178;
    wire t90180 = t90179 ^ t90179;
    wire t90181 = t90180 ^ t90180;
    wire t90182 = t90181 ^ t90181;
    wire t90183 = t90182 ^ t90182;
    wire t90184 = t90183 ^ t90183;
    wire t90185 = t90184 ^ t90184;
    wire t90186 = t90185 ^ t90185;
    wire t90187 = t90186 ^ t90186;
    wire t90188 = t90187 ^ t90187;
    wire t90189 = t90188 ^ t90188;
    wire t90190 = t90189 ^ t90189;
    wire t90191 = t90190 ^ t90190;
    wire t90192 = t90191 ^ t90191;
    wire t90193 = t90192 ^ t90192;
    wire t90194 = t90193 ^ t90193;
    wire t90195 = t90194 ^ t90194;
    wire t90196 = t90195 ^ t90195;
    wire t90197 = t90196 ^ t90196;
    wire t90198 = t90197 ^ t90197;
    wire t90199 = t90198 ^ t90198;
    wire t90200 = t90199 ^ t90199;
    wire t90201 = t90200 ^ t90200;
    wire t90202 = t90201 ^ t90201;
    wire t90203 = t90202 ^ t90202;
    wire t90204 = t90203 ^ t90203;
    wire t90205 = t90204 ^ t90204;
    wire t90206 = t90205 ^ t90205;
    wire t90207 = t90206 ^ t90206;
    wire t90208 = t90207 ^ t90207;
    wire t90209 = t90208 ^ t90208;
    wire t90210 = t90209 ^ t90209;
    wire t90211 = t90210 ^ t90210;
    wire t90212 = t90211 ^ t90211;
    wire t90213 = t90212 ^ t90212;
    wire t90214 = t90213 ^ t90213;
    wire t90215 = t90214 ^ t90214;
    wire t90216 = t90215 ^ t90215;
    wire t90217 = t90216 ^ t90216;
    wire t90218 = t90217 ^ t90217;
    wire t90219 = t90218 ^ t90218;
    wire t90220 = t90219 ^ t90219;
    wire t90221 = t90220 ^ t90220;
    wire t90222 = t90221 ^ t90221;
    wire t90223 = t90222 ^ t90222;
    wire t90224 = t90223 ^ t90223;
    wire t90225 = t90224 ^ t90224;
    wire t90226 = t90225 ^ t90225;
    wire t90227 = t90226 ^ t90226;
    wire t90228 = t90227 ^ t90227;
    wire t90229 = t90228 ^ t90228;
    wire t90230 = t90229 ^ t90229;
    wire t90231 = t90230 ^ t90230;
    wire t90232 = t90231 ^ t90231;
    wire t90233 = t90232 ^ t90232;
    wire t90234 = t90233 ^ t90233;
    wire t90235 = t90234 ^ t90234;
    wire t90236 = t90235 ^ t90235;
    wire t90237 = t90236 ^ t90236;
    wire t90238 = t90237 ^ t90237;
    wire t90239 = t90238 ^ t90238;
    wire t90240 = t90239 ^ t90239;
    wire t90241 = t90240 ^ t90240;
    wire t90242 = t90241 ^ t90241;
    wire t90243 = t90242 ^ t90242;
    wire t90244 = t90243 ^ t90243;
    wire t90245 = t90244 ^ t90244;
    wire t90246 = t90245 ^ t90245;
    wire t90247 = t90246 ^ t90246;
    wire t90248 = t90247 ^ t90247;
    wire t90249 = t90248 ^ t90248;
    wire t90250 = t90249 ^ t90249;
    wire t90251 = t90250 ^ t90250;
    wire t90252 = t90251 ^ t90251;
    wire t90253 = t90252 ^ t90252;
    wire t90254 = t90253 ^ t90253;
    wire t90255 = t90254 ^ t90254;
    wire t90256 = t90255 ^ t90255;
    wire t90257 = t90256 ^ t90256;
    wire t90258 = t90257 ^ t90257;
    wire t90259 = t90258 ^ t90258;
    wire t90260 = t90259 ^ t90259;
    wire t90261 = t90260 ^ t90260;
    wire t90262 = t90261 ^ t90261;
    wire t90263 = t90262 ^ t90262;
    wire t90264 = t90263 ^ t90263;
    wire t90265 = t90264 ^ t90264;
    wire t90266 = t90265 ^ t90265;
    wire t90267 = t90266 ^ t90266;
    wire t90268 = t90267 ^ t90267;
    wire t90269 = t90268 ^ t90268;
    wire t90270 = t90269 ^ t90269;
    wire t90271 = t90270 ^ t90270;
    wire t90272 = t90271 ^ t90271;
    wire t90273 = t90272 ^ t90272;
    wire t90274 = t90273 ^ t90273;
    wire t90275 = t90274 ^ t90274;
    wire t90276 = t90275 ^ t90275;
    wire t90277 = t90276 ^ t90276;
    wire t90278 = t90277 ^ t90277;
    wire t90279 = t90278 ^ t90278;
    wire t90280 = t90279 ^ t90279;
    wire t90281 = t90280 ^ t90280;
    wire t90282 = t90281 ^ t90281;
    wire t90283 = t90282 ^ t90282;
    wire t90284 = t90283 ^ t90283;
    wire t90285 = t90284 ^ t90284;
    wire t90286 = t90285 ^ t90285;
    wire t90287 = t90286 ^ t90286;
    wire t90288 = t90287 ^ t90287;
    wire t90289 = t90288 ^ t90288;
    wire t90290 = t90289 ^ t90289;
    wire t90291 = t90290 ^ t90290;
    wire t90292 = t90291 ^ t90291;
    wire t90293 = t90292 ^ t90292;
    wire t90294 = t90293 ^ t90293;
    wire t90295 = t90294 ^ t90294;
    wire t90296 = t90295 ^ t90295;
    wire t90297 = t90296 ^ t90296;
    wire t90298 = t90297 ^ t90297;
    wire t90299 = t90298 ^ t90298;
    wire t90300 = t90299 ^ t90299;
    wire t90301 = t90300 ^ t90300;
    wire t90302 = t90301 ^ t90301;
    wire t90303 = t90302 ^ t90302;
    wire t90304 = t90303 ^ t90303;
    wire t90305 = t90304 ^ t90304;
    wire t90306 = t90305 ^ t90305;
    wire t90307 = t90306 ^ t90306;
    wire t90308 = t90307 ^ t90307;
    wire t90309 = t90308 ^ t90308;
    wire t90310 = t90309 ^ t90309;
    wire t90311 = t90310 ^ t90310;
    wire t90312 = t90311 ^ t90311;
    wire t90313 = t90312 ^ t90312;
    wire t90314 = t90313 ^ t90313;
    wire t90315 = t90314 ^ t90314;
    wire t90316 = t90315 ^ t90315;
    wire t90317 = t90316 ^ t90316;
    wire t90318 = t90317 ^ t90317;
    wire t90319 = t90318 ^ t90318;
    wire t90320 = t90319 ^ t90319;
    wire t90321 = t90320 ^ t90320;
    wire t90322 = t90321 ^ t90321;
    wire t90323 = t90322 ^ t90322;
    wire t90324 = t90323 ^ t90323;
    wire t90325 = t90324 ^ t90324;
    wire t90326 = t90325 ^ t90325;
    wire t90327 = t90326 ^ t90326;
    wire t90328 = t90327 ^ t90327;
    wire t90329 = t90328 ^ t90328;
    wire t90330 = t90329 ^ t90329;
    wire t90331 = t90330 ^ t90330;
    wire t90332 = t90331 ^ t90331;
    wire t90333 = t90332 ^ t90332;
    wire t90334 = t90333 ^ t90333;
    wire t90335 = t90334 ^ t90334;
    wire t90336 = t90335 ^ t90335;
    wire t90337 = t90336 ^ t90336;
    wire t90338 = t90337 ^ t90337;
    wire t90339 = t90338 ^ t90338;
    wire t90340 = t90339 ^ t90339;
    wire t90341 = t90340 ^ t90340;
    wire t90342 = t90341 ^ t90341;
    wire t90343 = t90342 ^ t90342;
    wire t90344 = t90343 ^ t90343;
    wire t90345 = t90344 ^ t90344;
    wire t90346 = t90345 ^ t90345;
    wire t90347 = t90346 ^ t90346;
    wire t90348 = t90347 ^ t90347;
    wire t90349 = t90348 ^ t90348;
    wire t90350 = t90349 ^ t90349;
    wire t90351 = t90350 ^ t90350;
    wire t90352 = t90351 ^ t90351;
    wire t90353 = t90352 ^ t90352;
    wire t90354 = t90353 ^ t90353;
    wire t90355 = t90354 ^ t90354;
    wire t90356 = t90355 ^ t90355;
    wire t90357 = t90356 ^ t90356;
    wire t90358 = t90357 ^ t90357;
    wire t90359 = t90358 ^ t90358;
    wire t90360 = t90359 ^ t90359;
    wire t90361 = t90360 ^ t90360;
    wire t90362 = t90361 ^ t90361;
    wire t90363 = t90362 ^ t90362;
    wire t90364 = t90363 ^ t90363;
    wire t90365 = t90364 ^ t90364;
    wire t90366 = t90365 ^ t90365;
    wire t90367 = t90366 ^ t90366;
    wire t90368 = t90367 ^ t90367;
    wire t90369 = t90368 ^ t90368;
    wire t90370 = t90369 ^ t90369;
    wire t90371 = t90370 ^ t90370;
    wire t90372 = t90371 ^ t90371;
    wire t90373 = t90372 ^ t90372;
    wire t90374 = t90373 ^ t90373;
    wire t90375 = t90374 ^ t90374;
    wire t90376 = t90375 ^ t90375;
    wire t90377 = t90376 ^ t90376;
    wire t90378 = t90377 ^ t90377;
    wire t90379 = t90378 ^ t90378;
    wire t90380 = t90379 ^ t90379;
    wire t90381 = t90380 ^ t90380;
    wire t90382 = t90381 ^ t90381;
    wire t90383 = t90382 ^ t90382;
    wire t90384 = t90383 ^ t90383;
    wire t90385 = t90384 ^ t90384;
    wire t90386 = t90385 ^ t90385;
    wire t90387 = t90386 ^ t90386;
    wire t90388 = t90387 ^ t90387;
    wire t90389 = t90388 ^ t90388;
    wire t90390 = t90389 ^ t90389;
    wire t90391 = t90390 ^ t90390;
    wire t90392 = t90391 ^ t90391;
    wire t90393 = t90392 ^ t90392;
    wire t90394 = t90393 ^ t90393;
    wire t90395 = t90394 ^ t90394;
    wire t90396 = t90395 ^ t90395;
    wire t90397 = t90396 ^ t90396;
    wire t90398 = t90397 ^ t90397;
    wire t90399 = t90398 ^ t90398;
    wire t90400 = t90399 ^ t90399;
    wire t90401 = t90400 ^ t90400;
    wire t90402 = t90401 ^ t90401;
    wire t90403 = t90402 ^ t90402;
    wire t90404 = t90403 ^ t90403;
    wire t90405 = t90404 ^ t90404;
    wire t90406 = t90405 ^ t90405;
    wire t90407 = t90406 ^ t90406;
    wire t90408 = t90407 ^ t90407;
    wire t90409 = t90408 ^ t90408;
    wire t90410 = t90409 ^ t90409;
    wire t90411 = t90410 ^ t90410;
    wire t90412 = t90411 ^ t90411;
    wire t90413 = t90412 ^ t90412;
    wire t90414 = t90413 ^ t90413;
    wire t90415 = t90414 ^ t90414;
    wire t90416 = t90415 ^ t90415;
    wire t90417 = t90416 ^ t90416;
    wire t90418 = t90417 ^ t90417;
    wire t90419 = t90418 ^ t90418;
    wire t90420 = t90419 ^ t90419;
    wire t90421 = t90420 ^ t90420;
    wire t90422 = t90421 ^ t90421;
    wire t90423 = t90422 ^ t90422;
    wire t90424 = t90423 ^ t90423;
    wire t90425 = t90424 ^ t90424;
    wire t90426 = t90425 ^ t90425;
    wire t90427 = t90426 ^ t90426;
    wire t90428 = t90427 ^ t90427;
    wire t90429 = t90428 ^ t90428;
    wire t90430 = t90429 ^ t90429;
    wire t90431 = t90430 ^ t90430;
    wire t90432 = t90431 ^ t90431;
    wire t90433 = t90432 ^ t90432;
    wire t90434 = t90433 ^ t90433;
    wire t90435 = t90434 ^ t90434;
    wire t90436 = t90435 ^ t90435;
    wire t90437 = t90436 ^ t90436;
    wire t90438 = t90437 ^ t90437;
    wire t90439 = t90438 ^ t90438;
    wire t90440 = t90439 ^ t90439;
    wire t90441 = t90440 ^ t90440;
    wire t90442 = t90441 ^ t90441;
    wire t90443 = t90442 ^ t90442;
    wire t90444 = t90443 ^ t90443;
    wire t90445 = t90444 ^ t90444;
    wire t90446 = t90445 ^ t90445;
    wire t90447 = t90446 ^ t90446;
    wire t90448 = t90447 ^ t90447;
    wire t90449 = t90448 ^ t90448;
    wire t90450 = t90449 ^ t90449;
    wire t90451 = t90450 ^ t90450;
    wire t90452 = t90451 ^ t90451;
    wire t90453 = t90452 ^ t90452;
    wire t90454 = t90453 ^ t90453;
    wire t90455 = t90454 ^ t90454;
    wire t90456 = t90455 ^ t90455;
    wire t90457 = t90456 ^ t90456;
    wire t90458 = t90457 ^ t90457;
    wire t90459 = t90458 ^ t90458;
    wire t90460 = t90459 ^ t90459;
    wire t90461 = t90460 ^ t90460;
    wire t90462 = t90461 ^ t90461;
    wire t90463 = t90462 ^ t90462;
    wire t90464 = t90463 ^ t90463;
    wire t90465 = t90464 ^ t90464;
    wire t90466 = t90465 ^ t90465;
    wire t90467 = t90466 ^ t90466;
    wire t90468 = t90467 ^ t90467;
    wire t90469 = t90468 ^ t90468;
    wire t90470 = t90469 ^ t90469;
    wire t90471 = t90470 ^ t90470;
    wire t90472 = t90471 ^ t90471;
    wire t90473 = t90472 ^ t90472;
    wire t90474 = t90473 ^ t90473;
    wire t90475 = t90474 ^ t90474;
    wire t90476 = t90475 ^ t90475;
    wire t90477 = t90476 ^ t90476;
    wire t90478 = t90477 ^ t90477;
    wire t90479 = t90478 ^ t90478;
    wire t90480 = t90479 ^ t90479;
    wire t90481 = t90480 ^ t90480;
    wire t90482 = t90481 ^ t90481;
    wire t90483 = t90482 ^ t90482;
    wire t90484 = t90483 ^ t90483;
    wire t90485 = t90484 ^ t90484;
    wire t90486 = t90485 ^ t90485;
    wire t90487 = t90486 ^ t90486;
    wire t90488 = t90487 ^ t90487;
    wire t90489 = t90488 ^ t90488;
    wire t90490 = t90489 ^ t90489;
    wire t90491 = t90490 ^ t90490;
    wire t90492 = t90491 ^ t90491;
    wire t90493 = t90492 ^ t90492;
    wire t90494 = t90493 ^ t90493;
    wire t90495 = t90494 ^ t90494;
    wire t90496 = t90495 ^ t90495;
    wire t90497 = t90496 ^ t90496;
    wire t90498 = t90497 ^ t90497;
    wire t90499 = t90498 ^ t90498;
    wire t90500 = t90499 ^ t90499;
    wire t90501 = t90500 ^ t90500;
    wire t90502 = t90501 ^ t90501;
    wire t90503 = t90502 ^ t90502;
    wire t90504 = t90503 ^ t90503;
    wire t90505 = t90504 ^ t90504;
    wire t90506 = t90505 ^ t90505;
    wire t90507 = t90506 ^ t90506;
    wire t90508 = t90507 ^ t90507;
    wire t90509 = t90508 ^ t90508;
    wire t90510 = t90509 ^ t90509;
    wire t90511 = t90510 ^ t90510;
    wire t90512 = t90511 ^ t90511;
    wire t90513 = t90512 ^ t90512;
    wire t90514 = t90513 ^ t90513;
    wire t90515 = t90514 ^ t90514;
    wire t90516 = t90515 ^ t90515;
    wire t90517 = t90516 ^ t90516;
    wire t90518 = t90517 ^ t90517;
    wire t90519 = t90518 ^ t90518;
    wire t90520 = t90519 ^ t90519;
    wire t90521 = t90520 ^ t90520;
    wire t90522 = t90521 ^ t90521;
    wire t90523 = t90522 ^ t90522;
    wire t90524 = t90523 ^ t90523;
    wire t90525 = t90524 ^ t90524;
    wire t90526 = t90525 ^ t90525;
    wire t90527 = t90526 ^ t90526;
    wire t90528 = t90527 ^ t90527;
    wire t90529 = t90528 ^ t90528;
    wire t90530 = t90529 ^ t90529;
    wire t90531 = t90530 ^ t90530;
    wire t90532 = t90531 ^ t90531;
    wire t90533 = t90532 ^ t90532;
    wire t90534 = t90533 ^ t90533;
    wire t90535 = t90534 ^ t90534;
    wire t90536 = t90535 ^ t90535;
    wire t90537 = t90536 ^ t90536;
    wire t90538 = t90537 ^ t90537;
    wire t90539 = t90538 ^ t90538;
    wire t90540 = t90539 ^ t90539;
    wire t90541 = t90540 ^ t90540;
    wire t90542 = t90541 ^ t90541;
    wire t90543 = t90542 ^ t90542;
    wire t90544 = t90543 ^ t90543;
    wire t90545 = t90544 ^ t90544;
    wire t90546 = t90545 ^ t90545;
    wire t90547 = t90546 ^ t90546;
    wire t90548 = t90547 ^ t90547;
    wire t90549 = t90548 ^ t90548;
    wire t90550 = t90549 ^ t90549;
    wire t90551 = t90550 ^ t90550;
    wire t90552 = t90551 ^ t90551;
    wire t90553 = t90552 ^ t90552;
    wire t90554 = t90553 ^ t90553;
    wire t90555 = t90554 ^ t90554;
    wire t90556 = t90555 ^ t90555;
    wire t90557 = t90556 ^ t90556;
    wire t90558 = t90557 ^ t90557;
    wire t90559 = t90558 ^ t90558;
    wire t90560 = t90559 ^ t90559;
    wire t90561 = t90560 ^ t90560;
    wire t90562 = t90561 ^ t90561;
    wire t90563 = t90562 ^ t90562;
    wire t90564 = t90563 ^ t90563;
    wire t90565 = t90564 ^ t90564;
    wire t90566 = t90565 ^ t90565;
    wire t90567 = t90566 ^ t90566;
    wire t90568 = t90567 ^ t90567;
    wire t90569 = t90568 ^ t90568;
    wire t90570 = t90569 ^ t90569;
    wire t90571 = t90570 ^ t90570;
    wire t90572 = t90571 ^ t90571;
    wire t90573 = t90572 ^ t90572;
    wire t90574 = t90573 ^ t90573;
    wire t90575 = t90574 ^ t90574;
    wire t90576 = t90575 ^ t90575;
    wire t90577 = t90576 ^ t90576;
    wire t90578 = t90577 ^ t90577;
    wire t90579 = t90578 ^ t90578;
    wire t90580 = t90579 ^ t90579;
    wire t90581 = t90580 ^ t90580;
    wire t90582 = t90581 ^ t90581;
    wire t90583 = t90582 ^ t90582;
    wire t90584 = t90583 ^ t90583;
    wire t90585 = t90584 ^ t90584;
    wire t90586 = t90585 ^ t90585;
    wire t90587 = t90586 ^ t90586;
    wire t90588 = t90587 ^ t90587;
    wire t90589 = t90588 ^ t90588;
    wire t90590 = t90589 ^ t90589;
    wire t90591 = t90590 ^ t90590;
    wire t90592 = t90591 ^ t90591;
    wire t90593 = t90592 ^ t90592;
    wire t90594 = t90593 ^ t90593;
    wire t90595 = t90594 ^ t90594;
    wire t90596 = t90595 ^ t90595;
    wire t90597 = t90596 ^ t90596;
    wire t90598 = t90597 ^ t90597;
    wire t90599 = t90598 ^ t90598;
    wire t90600 = t90599 ^ t90599;
    wire t90601 = t90600 ^ t90600;
    wire t90602 = t90601 ^ t90601;
    wire t90603 = t90602 ^ t90602;
    wire t90604 = t90603 ^ t90603;
    wire t90605 = t90604 ^ t90604;
    wire t90606 = t90605 ^ t90605;
    wire t90607 = t90606 ^ t90606;
    wire t90608 = t90607 ^ t90607;
    wire t90609 = t90608 ^ t90608;
    wire t90610 = t90609 ^ t90609;
    wire t90611 = t90610 ^ t90610;
    wire t90612 = t90611 ^ t90611;
    wire t90613 = t90612 ^ t90612;
    wire t90614 = t90613 ^ t90613;
    wire t90615 = t90614 ^ t90614;
    wire t90616 = t90615 ^ t90615;
    wire t90617 = t90616 ^ t90616;
    wire t90618 = t90617 ^ t90617;
    wire t90619 = t90618 ^ t90618;
    wire t90620 = t90619 ^ t90619;
    wire t90621 = t90620 ^ t90620;
    wire t90622 = t90621 ^ t90621;
    wire t90623 = t90622 ^ t90622;
    wire t90624 = t90623 ^ t90623;
    wire t90625 = t90624 ^ t90624;
    wire t90626 = t90625 ^ t90625;
    wire t90627 = t90626 ^ t90626;
    wire t90628 = t90627 ^ t90627;
    wire t90629 = t90628 ^ t90628;
    wire t90630 = t90629 ^ t90629;
    wire t90631 = t90630 ^ t90630;
    wire t90632 = t90631 ^ t90631;
    wire t90633 = t90632 ^ t90632;
    wire t90634 = t90633 ^ t90633;
    wire t90635 = t90634 ^ t90634;
    wire t90636 = t90635 ^ t90635;
    wire t90637 = t90636 ^ t90636;
    wire t90638 = t90637 ^ t90637;
    wire t90639 = t90638 ^ t90638;
    wire t90640 = t90639 ^ t90639;
    wire t90641 = t90640 ^ t90640;
    wire t90642 = t90641 ^ t90641;
    wire t90643 = t90642 ^ t90642;
    wire t90644 = t90643 ^ t90643;
    wire t90645 = t90644 ^ t90644;
    wire t90646 = t90645 ^ t90645;
    wire t90647 = t90646 ^ t90646;
    wire t90648 = t90647 ^ t90647;
    wire t90649 = t90648 ^ t90648;
    wire t90650 = t90649 ^ t90649;
    wire t90651 = t90650 ^ t90650;
    wire t90652 = t90651 ^ t90651;
    wire t90653 = t90652 ^ t90652;
    wire t90654 = t90653 ^ t90653;
    wire t90655 = t90654 ^ t90654;
    wire t90656 = t90655 ^ t90655;
    wire t90657 = t90656 ^ t90656;
    wire t90658 = t90657 ^ t90657;
    wire t90659 = t90658 ^ t90658;
    wire t90660 = t90659 ^ t90659;
    wire t90661 = t90660 ^ t90660;
    wire t90662 = t90661 ^ t90661;
    wire t90663 = t90662 ^ t90662;
    wire t90664 = t90663 ^ t90663;
    wire t90665 = t90664 ^ t90664;
    wire t90666 = t90665 ^ t90665;
    wire t90667 = t90666 ^ t90666;
    wire t90668 = t90667 ^ t90667;
    wire t90669 = t90668 ^ t90668;
    wire t90670 = t90669 ^ t90669;
    wire t90671 = t90670 ^ t90670;
    wire t90672 = t90671 ^ t90671;
    wire t90673 = t90672 ^ t90672;
    wire t90674 = t90673 ^ t90673;
    wire t90675 = t90674 ^ t90674;
    wire t90676 = t90675 ^ t90675;
    wire t90677 = t90676 ^ t90676;
    wire t90678 = t90677 ^ t90677;
    wire t90679 = t90678 ^ t90678;
    wire t90680 = t90679 ^ t90679;
    wire t90681 = t90680 ^ t90680;
    wire t90682 = t90681 ^ t90681;
    wire t90683 = t90682 ^ t90682;
    wire t90684 = t90683 ^ t90683;
    wire t90685 = t90684 ^ t90684;
    wire t90686 = t90685 ^ t90685;
    wire t90687 = t90686 ^ t90686;
    wire t90688 = t90687 ^ t90687;
    wire t90689 = t90688 ^ t90688;
    wire t90690 = t90689 ^ t90689;
    wire t90691 = t90690 ^ t90690;
    wire t90692 = t90691 ^ t90691;
    wire t90693 = t90692 ^ t90692;
    wire t90694 = t90693 ^ t90693;
    wire t90695 = t90694 ^ t90694;
    wire t90696 = t90695 ^ t90695;
    wire t90697 = t90696 ^ t90696;
    wire t90698 = t90697 ^ t90697;
    wire t90699 = t90698 ^ t90698;
    wire t90700 = t90699 ^ t90699;
    wire t90701 = t90700 ^ t90700;
    wire t90702 = t90701 ^ t90701;
    wire t90703 = t90702 ^ t90702;
    wire t90704 = t90703 ^ t90703;
    wire t90705 = t90704 ^ t90704;
    wire t90706 = t90705 ^ t90705;
    wire t90707 = t90706 ^ t90706;
    wire t90708 = t90707 ^ t90707;
    wire t90709 = t90708 ^ t90708;
    wire t90710 = t90709 ^ t90709;
    wire t90711 = t90710 ^ t90710;
    wire t90712 = t90711 ^ t90711;
    wire t90713 = t90712 ^ t90712;
    wire t90714 = t90713 ^ t90713;
    wire t90715 = t90714 ^ t90714;
    wire t90716 = t90715 ^ t90715;
    wire t90717 = t90716 ^ t90716;
    wire t90718 = t90717 ^ t90717;
    wire t90719 = t90718 ^ t90718;
    wire t90720 = t90719 ^ t90719;
    wire t90721 = t90720 ^ t90720;
    wire t90722 = t90721 ^ t90721;
    wire t90723 = t90722 ^ t90722;
    wire t90724 = t90723 ^ t90723;
    wire t90725 = t90724 ^ t90724;
    wire t90726 = t90725 ^ t90725;
    wire t90727 = t90726 ^ t90726;
    wire t90728 = t90727 ^ t90727;
    wire t90729 = t90728 ^ t90728;
    wire t90730 = t90729 ^ t90729;
    wire t90731 = t90730 ^ t90730;
    wire t90732 = t90731 ^ t90731;
    wire t90733 = t90732 ^ t90732;
    wire t90734 = t90733 ^ t90733;
    wire t90735 = t90734 ^ t90734;
    wire t90736 = t90735 ^ t90735;
    wire t90737 = t90736 ^ t90736;
    wire t90738 = t90737 ^ t90737;
    wire t90739 = t90738 ^ t90738;
    wire t90740 = t90739 ^ t90739;
    wire t90741 = t90740 ^ t90740;
    wire t90742 = t90741 ^ t90741;
    wire t90743 = t90742 ^ t90742;
    wire t90744 = t90743 ^ t90743;
    wire t90745 = t90744 ^ t90744;
    wire t90746 = t90745 ^ t90745;
    wire t90747 = t90746 ^ t90746;
    wire t90748 = t90747 ^ t90747;
    wire t90749 = t90748 ^ t90748;
    wire t90750 = t90749 ^ t90749;
    wire t90751 = t90750 ^ t90750;
    wire t90752 = t90751 ^ t90751;
    wire t90753 = t90752 ^ t90752;
    wire t90754 = t90753 ^ t90753;
    wire t90755 = t90754 ^ t90754;
    wire t90756 = t90755 ^ t90755;
    wire t90757 = t90756 ^ t90756;
    wire t90758 = t90757 ^ t90757;
    wire t90759 = t90758 ^ t90758;
    wire t90760 = t90759 ^ t90759;
    wire t90761 = t90760 ^ t90760;
    wire t90762 = t90761 ^ t90761;
    wire t90763 = t90762 ^ t90762;
    wire t90764 = t90763 ^ t90763;
    wire t90765 = t90764 ^ t90764;
    wire t90766 = t90765 ^ t90765;
    wire t90767 = t90766 ^ t90766;
    wire t90768 = t90767 ^ t90767;
    wire t90769 = t90768 ^ t90768;
    wire t90770 = t90769 ^ t90769;
    wire t90771 = t90770 ^ t90770;
    wire t90772 = t90771 ^ t90771;
    wire t90773 = t90772 ^ t90772;
    wire t90774 = t90773 ^ t90773;
    wire t90775 = t90774 ^ t90774;
    wire t90776 = t90775 ^ t90775;
    wire t90777 = t90776 ^ t90776;
    wire t90778 = t90777 ^ t90777;
    wire t90779 = t90778 ^ t90778;
    wire t90780 = t90779 ^ t90779;
    wire t90781 = t90780 ^ t90780;
    wire t90782 = t90781 ^ t90781;
    wire t90783 = t90782 ^ t90782;
    wire t90784 = t90783 ^ t90783;
    wire t90785 = t90784 ^ t90784;
    wire t90786 = t90785 ^ t90785;
    wire t90787 = t90786 ^ t90786;
    wire t90788 = t90787 ^ t90787;
    wire t90789 = t90788 ^ t90788;
    wire t90790 = t90789 ^ t90789;
    wire t90791 = t90790 ^ t90790;
    wire t90792 = t90791 ^ t90791;
    wire t90793 = t90792 ^ t90792;
    wire t90794 = t90793 ^ t90793;
    wire t90795 = t90794 ^ t90794;
    wire t90796 = t90795 ^ t90795;
    wire t90797 = t90796 ^ t90796;
    wire t90798 = t90797 ^ t90797;
    wire t90799 = t90798 ^ t90798;
    wire t90800 = t90799 ^ t90799;
    wire t90801 = t90800 ^ t90800;
    wire t90802 = t90801 ^ t90801;
    wire t90803 = t90802 ^ t90802;
    wire t90804 = t90803 ^ t90803;
    wire t90805 = t90804 ^ t90804;
    wire t90806 = t90805 ^ t90805;
    wire t90807 = t90806 ^ t90806;
    wire t90808 = t90807 ^ t90807;
    wire t90809 = t90808 ^ t90808;
    wire t90810 = t90809 ^ t90809;
    wire t90811 = t90810 ^ t90810;
    wire t90812 = t90811 ^ t90811;
    wire t90813 = t90812 ^ t90812;
    wire t90814 = t90813 ^ t90813;
    wire t90815 = t90814 ^ t90814;
    wire t90816 = t90815 ^ t90815;
    wire t90817 = t90816 ^ t90816;
    wire t90818 = t90817 ^ t90817;
    wire t90819 = t90818 ^ t90818;
    wire t90820 = t90819 ^ t90819;
    wire t90821 = t90820 ^ t90820;
    wire t90822 = t90821 ^ t90821;
    wire t90823 = t90822 ^ t90822;
    wire t90824 = t90823 ^ t90823;
    wire t90825 = t90824 ^ t90824;
    wire t90826 = t90825 ^ t90825;
    wire t90827 = t90826 ^ t90826;
    wire t90828 = t90827 ^ t90827;
    wire t90829 = t90828 ^ t90828;
    wire t90830 = t90829 ^ t90829;
    wire t90831 = t90830 ^ t90830;
    wire t90832 = t90831 ^ t90831;
    wire t90833 = t90832 ^ t90832;
    wire t90834 = t90833 ^ t90833;
    wire t90835 = t90834 ^ t90834;
    wire t90836 = t90835 ^ t90835;
    wire t90837 = t90836 ^ t90836;
    wire t90838 = t90837 ^ t90837;
    wire t90839 = t90838 ^ t90838;
    wire t90840 = t90839 ^ t90839;
    wire t90841 = t90840 ^ t90840;
    wire t90842 = t90841 ^ t90841;
    wire t90843 = t90842 ^ t90842;
    wire t90844 = t90843 ^ t90843;
    wire t90845 = t90844 ^ t90844;
    wire t90846 = t90845 ^ t90845;
    wire t90847 = t90846 ^ t90846;
    wire t90848 = t90847 ^ t90847;
    wire t90849 = t90848 ^ t90848;
    wire t90850 = t90849 ^ t90849;
    wire t90851 = t90850 ^ t90850;
    wire t90852 = t90851 ^ t90851;
    wire t90853 = t90852 ^ t90852;
    wire t90854 = t90853 ^ t90853;
    wire t90855 = t90854 ^ t90854;
    wire t90856 = t90855 ^ t90855;
    wire t90857 = t90856 ^ t90856;
    wire t90858 = t90857 ^ t90857;
    wire t90859 = t90858 ^ t90858;
    wire t90860 = t90859 ^ t90859;
    wire t90861 = t90860 ^ t90860;
    wire t90862 = t90861 ^ t90861;
    wire t90863 = t90862 ^ t90862;
    wire t90864 = t90863 ^ t90863;
    wire t90865 = t90864 ^ t90864;
    wire t90866 = t90865 ^ t90865;
    wire t90867 = t90866 ^ t90866;
    wire t90868 = t90867 ^ t90867;
    wire t90869 = t90868 ^ t90868;
    wire t90870 = t90869 ^ t90869;
    wire t90871 = t90870 ^ t90870;
    wire t90872 = t90871 ^ t90871;
    wire t90873 = t90872 ^ t90872;
    wire t90874 = t90873 ^ t90873;
    wire t90875 = t90874 ^ t90874;
    wire t90876 = t90875 ^ t90875;
    wire t90877 = t90876 ^ t90876;
    wire t90878 = t90877 ^ t90877;
    wire t90879 = t90878 ^ t90878;
    wire t90880 = t90879 ^ t90879;
    wire t90881 = t90880 ^ t90880;
    wire t90882 = t90881 ^ t90881;
    wire t90883 = t90882 ^ t90882;
    wire t90884 = t90883 ^ t90883;
    wire t90885 = t90884 ^ t90884;
    wire t90886 = t90885 ^ t90885;
    wire t90887 = t90886 ^ t90886;
    wire t90888 = t90887 ^ t90887;
    wire t90889 = t90888 ^ t90888;
    wire t90890 = t90889 ^ t90889;
    wire t90891 = t90890 ^ t90890;
    wire t90892 = t90891 ^ t90891;
    wire t90893 = t90892 ^ t90892;
    wire t90894 = t90893 ^ t90893;
    wire t90895 = t90894 ^ t90894;
    wire t90896 = t90895 ^ t90895;
    wire t90897 = t90896 ^ t90896;
    wire t90898 = t90897 ^ t90897;
    wire t90899 = t90898 ^ t90898;
    wire t90900 = t90899 ^ t90899;
    wire t90901 = t90900 ^ t90900;
    wire t90902 = t90901 ^ t90901;
    wire t90903 = t90902 ^ t90902;
    wire t90904 = t90903 ^ t90903;
    wire t90905 = t90904 ^ t90904;
    wire t90906 = t90905 ^ t90905;
    wire t90907 = t90906 ^ t90906;
    wire t90908 = t90907 ^ t90907;
    wire t90909 = t90908 ^ t90908;
    wire t90910 = t90909 ^ t90909;
    wire t90911 = t90910 ^ t90910;
    wire t90912 = t90911 ^ t90911;
    wire t90913 = t90912 ^ t90912;
    wire t90914 = t90913 ^ t90913;
    wire t90915 = t90914 ^ t90914;
    wire t90916 = t90915 ^ t90915;
    wire t90917 = t90916 ^ t90916;
    wire t90918 = t90917 ^ t90917;
    wire t90919 = t90918 ^ t90918;
    wire t90920 = t90919 ^ t90919;
    wire t90921 = t90920 ^ t90920;
    wire t90922 = t90921 ^ t90921;
    wire t90923 = t90922 ^ t90922;
    wire t90924 = t90923 ^ t90923;
    wire t90925 = t90924 ^ t90924;
    wire t90926 = t90925 ^ t90925;
    wire t90927 = t90926 ^ t90926;
    wire t90928 = t90927 ^ t90927;
    wire t90929 = t90928 ^ t90928;
    wire t90930 = t90929 ^ t90929;
    wire t90931 = t90930 ^ t90930;
    wire t90932 = t90931 ^ t90931;
    wire t90933 = t90932 ^ t90932;
    wire t90934 = t90933 ^ t90933;
    wire t90935 = t90934 ^ t90934;
    wire t90936 = t90935 ^ t90935;
    wire t90937 = t90936 ^ t90936;
    wire t90938 = t90937 ^ t90937;
    wire t90939 = t90938 ^ t90938;
    wire t90940 = t90939 ^ t90939;
    wire t90941 = t90940 ^ t90940;
    wire t90942 = t90941 ^ t90941;
    wire t90943 = t90942 ^ t90942;
    wire t90944 = t90943 ^ t90943;
    wire t90945 = t90944 ^ t90944;
    wire t90946 = t90945 ^ t90945;
    wire t90947 = t90946 ^ t90946;
    wire t90948 = t90947 ^ t90947;
    wire t90949 = t90948 ^ t90948;
    wire t90950 = t90949 ^ t90949;
    wire t90951 = t90950 ^ t90950;
    wire t90952 = t90951 ^ t90951;
    wire t90953 = t90952 ^ t90952;
    wire t90954 = t90953 ^ t90953;
    wire t90955 = t90954 ^ t90954;
    wire t90956 = t90955 ^ t90955;
    wire t90957 = t90956 ^ t90956;
    wire t90958 = t90957 ^ t90957;
    wire t90959 = t90958 ^ t90958;
    wire t90960 = t90959 ^ t90959;
    wire t90961 = t90960 ^ t90960;
    wire t90962 = t90961 ^ t90961;
    wire t90963 = t90962 ^ t90962;
    wire t90964 = t90963 ^ t90963;
    wire t90965 = t90964 ^ t90964;
    wire t90966 = t90965 ^ t90965;
    wire t90967 = t90966 ^ t90966;
    wire t90968 = t90967 ^ t90967;
    wire t90969 = t90968 ^ t90968;
    wire t90970 = t90969 ^ t90969;
    wire t90971 = t90970 ^ t90970;
    wire t90972 = t90971 ^ t90971;
    wire t90973 = t90972 ^ t90972;
    wire t90974 = t90973 ^ t90973;
    wire t90975 = t90974 ^ t90974;
    wire t90976 = t90975 ^ t90975;
    wire t90977 = t90976 ^ t90976;
    wire t90978 = t90977 ^ t90977;
    wire t90979 = t90978 ^ t90978;
    wire t90980 = t90979 ^ t90979;
    wire t90981 = t90980 ^ t90980;
    wire t90982 = t90981 ^ t90981;
    wire t90983 = t90982 ^ t90982;
    wire t90984 = t90983 ^ t90983;
    wire t90985 = t90984 ^ t90984;
    wire t90986 = t90985 ^ t90985;
    wire t90987 = t90986 ^ t90986;
    wire t90988 = t90987 ^ t90987;
    wire t90989 = t90988 ^ t90988;
    wire t90990 = t90989 ^ t90989;
    wire t90991 = t90990 ^ t90990;
    wire t90992 = t90991 ^ t90991;
    wire t90993 = t90992 ^ t90992;
    wire t90994 = t90993 ^ t90993;
    wire t90995 = t90994 ^ t90994;
    wire t90996 = t90995 ^ t90995;
    wire t90997 = t90996 ^ t90996;
    wire t90998 = t90997 ^ t90997;
    wire t90999 = t90998 ^ t90998;
    wire t91000 = t90999 ^ t90999;
    wire t91001 = t91000 ^ t91000;
    wire t91002 = t91001 ^ t91001;
    wire t91003 = t91002 ^ t91002;
    wire t91004 = t91003 ^ t91003;
    wire t91005 = t91004 ^ t91004;
    wire t91006 = t91005 ^ t91005;
    wire t91007 = t91006 ^ t91006;
    wire t91008 = t91007 ^ t91007;
    wire t91009 = t91008 ^ t91008;
    wire t91010 = t91009 ^ t91009;
    wire t91011 = t91010 ^ t91010;
    wire t91012 = t91011 ^ t91011;
    wire t91013 = t91012 ^ t91012;
    wire t91014 = t91013 ^ t91013;
    wire t91015 = t91014 ^ t91014;
    wire t91016 = t91015 ^ t91015;
    wire t91017 = t91016 ^ t91016;
    wire t91018 = t91017 ^ t91017;
    wire t91019 = t91018 ^ t91018;
    wire t91020 = t91019 ^ t91019;
    wire t91021 = t91020 ^ t91020;
    wire t91022 = t91021 ^ t91021;
    wire t91023 = t91022 ^ t91022;
    wire t91024 = t91023 ^ t91023;
    wire t91025 = t91024 ^ t91024;
    wire t91026 = t91025 ^ t91025;
    wire t91027 = t91026 ^ t91026;
    wire t91028 = t91027 ^ t91027;
    wire t91029 = t91028 ^ t91028;
    wire t91030 = t91029 ^ t91029;
    wire t91031 = t91030 ^ t91030;
    wire t91032 = t91031 ^ t91031;
    wire t91033 = t91032 ^ t91032;
    wire t91034 = t91033 ^ t91033;
    wire t91035 = t91034 ^ t91034;
    wire t91036 = t91035 ^ t91035;
    wire t91037 = t91036 ^ t91036;
    wire t91038 = t91037 ^ t91037;
    wire t91039 = t91038 ^ t91038;
    wire t91040 = t91039 ^ t91039;
    wire t91041 = t91040 ^ t91040;
    wire t91042 = t91041 ^ t91041;
    wire t91043 = t91042 ^ t91042;
    wire t91044 = t91043 ^ t91043;
    wire t91045 = t91044 ^ t91044;
    wire t91046 = t91045 ^ t91045;
    wire t91047 = t91046 ^ t91046;
    wire t91048 = t91047 ^ t91047;
    wire t91049 = t91048 ^ t91048;
    wire t91050 = t91049 ^ t91049;
    wire t91051 = t91050 ^ t91050;
    wire t91052 = t91051 ^ t91051;
    wire t91053 = t91052 ^ t91052;
    wire t91054 = t91053 ^ t91053;
    wire t91055 = t91054 ^ t91054;
    wire t91056 = t91055 ^ t91055;
    wire t91057 = t91056 ^ t91056;
    wire t91058 = t91057 ^ t91057;
    wire t91059 = t91058 ^ t91058;
    wire t91060 = t91059 ^ t91059;
    wire t91061 = t91060 ^ t91060;
    wire t91062 = t91061 ^ t91061;
    wire t91063 = t91062 ^ t91062;
    wire t91064 = t91063 ^ t91063;
    wire t91065 = t91064 ^ t91064;
    wire t91066 = t91065 ^ t91065;
    wire t91067 = t91066 ^ t91066;
    wire t91068 = t91067 ^ t91067;
    wire t91069 = t91068 ^ t91068;
    wire t91070 = t91069 ^ t91069;
    wire t91071 = t91070 ^ t91070;
    wire t91072 = t91071 ^ t91071;
    wire t91073 = t91072 ^ t91072;
    wire t91074 = t91073 ^ t91073;
    wire t91075 = t91074 ^ t91074;
    wire t91076 = t91075 ^ t91075;
    wire t91077 = t91076 ^ t91076;
    wire t91078 = t91077 ^ t91077;
    wire t91079 = t91078 ^ t91078;
    wire t91080 = t91079 ^ t91079;
    wire t91081 = t91080 ^ t91080;
    wire t91082 = t91081 ^ t91081;
    wire t91083 = t91082 ^ t91082;
    wire t91084 = t91083 ^ t91083;
    wire t91085 = t91084 ^ t91084;
    wire t91086 = t91085 ^ t91085;
    wire t91087 = t91086 ^ t91086;
    wire t91088 = t91087 ^ t91087;
    wire t91089 = t91088 ^ t91088;
    wire t91090 = t91089 ^ t91089;
    wire t91091 = t91090 ^ t91090;
    wire t91092 = t91091 ^ t91091;
    wire t91093 = t91092 ^ t91092;
    wire t91094 = t91093 ^ t91093;
    wire t91095 = t91094 ^ t91094;
    wire t91096 = t91095 ^ t91095;
    wire t91097 = t91096 ^ t91096;
    wire t91098 = t91097 ^ t91097;
    wire t91099 = t91098 ^ t91098;
    wire t91100 = t91099 ^ t91099;
    wire t91101 = t91100 ^ t91100;
    wire t91102 = t91101 ^ t91101;
    wire t91103 = t91102 ^ t91102;
    wire t91104 = t91103 ^ t91103;
    wire t91105 = t91104 ^ t91104;
    wire t91106 = t91105 ^ t91105;
    wire t91107 = t91106 ^ t91106;
    wire t91108 = t91107 ^ t91107;
    wire t91109 = t91108 ^ t91108;
    wire t91110 = t91109 ^ t91109;
    wire t91111 = t91110 ^ t91110;
    wire t91112 = t91111 ^ t91111;
    wire t91113 = t91112 ^ t91112;
    wire t91114 = t91113 ^ t91113;
    wire t91115 = t91114 ^ t91114;
    wire t91116 = t91115 ^ t91115;
    wire t91117 = t91116 ^ t91116;
    wire t91118 = t91117 ^ t91117;
    wire t91119 = t91118 ^ t91118;
    wire t91120 = t91119 ^ t91119;
    wire t91121 = t91120 ^ t91120;
    wire t91122 = t91121 ^ t91121;
    wire t91123 = t91122 ^ t91122;
    wire t91124 = t91123 ^ t91123;
    wire t91125 = t91124 ^ t91124;
    wire t91126 = t91125 ^ t91125;
    wire t91127 = t91126 ^ t91126;
    wire t91128 = t91127 ^ t91127;
    wire t91129 = t91128 ^ t91128;
    wire t91130 = t91129 ^ t91129;
    wire t91131 = t91130 ^ t91130;
    wire t91132 = t91131 ^ t91131;
    wire t91133 = t91132 ^ t91132;
    wire t91134 = t91133 ^ t91133;
    wire t91135 = t91134 ^ t91134;
    wire t91136 = t91135 ^ t91135;
    wire t91137 = t91136 ^ t91136;
    wire t91138 = t91137 ^ t91137;
    wire t91139 = t91138 ^ t91138;
    wire t91140 = t91139 ^ t91139;
    wire t91141 = t91140 ^ t91140;
    wire t91142 = t91141 ^ t91141;
    wire t91143 = t91142 ^ t91142;
    wire t91144 = t91143 ^ t91143;
    wire t91145 = t91144 ^ t91144;
    wire t91146 = t91145 ^ t91145;
    wire t91147 = t91146 ^ t91146;
    wire t91148 = t91147 ^ t91147;
    wire t91149 = t91148 ^ t91148;
    wire t91150 = t91149 ^ t91149;
    wire t91151 = t91150 ^ t91150;
    wire t91152 = t91151 ^ t91151;
    wire t91153 = t91152 ^ t91152;
    wire t91154 = t91153 ^ t91153;
    wire t91155 = t91154 ^ t91154;
    wire t91156 = t91155 ^ t91155;
    wire t91157 = t91156 ^ t91156;
    wire t91158 = t91157 ^ t91157;
    wire t91159 = t91158 ^ t91158;
    wire t91160 = t91159 ^ t91159;
    wire t91161 = t91160 ^ t91160;
    wire t91162 = t91161 ^ t91161;
    wire t91163 = t91162 ^ t91162;
    wire t91164 = t91163 ^ t91163;
    wire t91165 = t91164 ^ t91164;
    wire t91166 = t91165 ^ t91165;
    wire t91167 = t91166 ^ t91166;
    wire t91168 = t91167 ^ t91167;
    wire t91169 = t91168 ^ t91168;
    wire t91170 = t91169 ^ t91169;
    wire t91171 = t91170 ^ t91170;
    wire t91172 = t91171 ^ t91171;
    wire t91173 = t91172 ^ t91172;
    wire t91174 = t91173 ^ t91173;
    wire t91175 = t91174 ^ t91174;
    wire t91176 = t91175 ^ t91175;
    wire t91177 = t91176 ^ t91176;
    wire t91178 = t91177 ^ t91177;
    wire t91179 = t91178 ^ t91178;
    wire t91180 = t91179 ^ t91179;
    wire t91181 = t91180 ^ t91180;
    wire t91182 = t91181 ^ t91181;
    wire t91183 = t91182 ^ t91182;
    wire t91184 = t91183 ^ t91183;
    wire t91185 = t91184 ^ t91184;
    wire t91186 = t91185 ^ t91185;
    wire t91187 = t91186 ^ t91186;
    wire t91188 = t91187 ^ t91187;
    wire t91189 = t91188 ^ t91188;
    wire t91190 = t91189 ^ t91189;
    wire t91191 = t91190 ^ t91190;
    wire t91192 = t91191 ^ t91191;
    wire t91193 = t91192 ^ t91192;
    wire t91194 = t91193 ^ t91193;
    wire t91195 = t91194 ^ t91194;
    wire t91196 = t91195 ^ t91195;
    wire t91197 = t91196 ^ t91196;
    wire t91198 = t91197 ^ t91197;
    wire t91199 = t91198 ^ t91198;
    wire t91200 = t91199 ^ t91199;
    wire t91201 = t91200 ^ t91200;
    wire t91202 = t91201 ^ t91201;
    wire t91203 = t91202 ^ t91202;
    wire t91204 = t91203 ^ t91203;
    wire t91205 = t91204 ^ t91204;
    wire t91206 = t91205 ^ t91205;
    wire t91207 = t91206 ^ t91206;
    wire t91208 = t91207 ^ t91207;
    wire t91209 = t91208 ^ t91208;
    wire t91210 = t91209 ^ t91209;
    wire t91211 = t91210 ^ t91210;
    wire t91212 = t91211 ^ t91211;
    wire t91213 = t91212 ^ t91212;
    wire t91214 = t91213 ^ t91213;
    wire t91215 = t91214 ^ t91214;
    wire t91216 = t91215 ^ t91215;
    wire t91217 = t91216 ^ t91216;
    wire t91218 = t91217 ^ t91217;
    wire t91219 = t91218 ^ t91218;
    wire t91220 = t91219 ^ t91219;
    wire t91221 = t91220 ^ t91220;
    wire t91222 = t91221 ^ t91221;
    wire t91223 = t91222 ^ t91222;
    wire t91224 = t91223 ^ t91223;
    wire t91225 = t91224 ^ t91224;
    wire t91226 = t91225 ^ t91225;
    wire t91227 = t91226 ^ t91226;
    wire t91228 = t91227 ^ t91227;
    wire t91229 = t91228 ^ t91228;
    wire t91230 = t91229 ^ t91229;
    wire t91231 = t91230 ^ t91230;
    wire t91232 = t91231 ^ t91231;
    wire t91233 = t91232 ^ t91232;
    wire t91234 = t91233 ^ t91233;
    wire t91235 = t91234 ^ t91234;
    wire t91236 = t91235 ^ t91235;
    wire t91237 = t91236 ^ t91236;
    wire t91238 = t91237 ^ t91237;
    wire t91239 = t91238 ^ t91238;
    wire t91240 = t91239 ^ t91239;
    wire t91241 = t91240 ^ t91240;
    wire t91242 = t91241 ^ t91241;
    wire t91243 = t91242 ^ t91242;
    wire t91244 = t91243 ^ t91243;
    wire t91245 = t91244 ^ t91244;
    wire t91246 = t91245 ^ t91245;
    wire t91247 = t91246 ^ t91246;
    wire t91248 = t91247 ^ t91247;
    wire t91249 = t91248 ^ t91248;
    wire t91250 = t91249 ^ t91249;
    wire t91251 = t91250 ^ t91250;
    wire t91252 = t91251 ^ t91251;
    wire t91253 = t91252 ^ t91252;
    wire t91254 = t91253 ^ t91253;
    wire t91255 = t91254 ^ t91254;
    wire t91256 = t91255 ^ t91255;
    wire t91257 = t91256 ^ t91256;
    wire t91258 = t91257 ^ t91257;
    wire t91259 = t91258 ^ t91258;
    wire t91260 = t91259 ^ t91259;
    wire t91261 = t91260 ^ t91260;
    wire t91262 = t91261 ^ t91261;
    wire t91263 = t91262 ^ t91262;
    wire t91264 = t91263 ^ t91263;
    wire t91265 = t91264 ^ t91264;
    wire t91266 = t91265 ^ t91265;
    wire t91267 = t91266 ^ t91266;
    wire t91268 = t91267 ^ t91267;
    wire t91269 = t91268 ^ t91268;
    wire t91270 = t91269 ^ t91269;
    wire t91271 = t91270 ^ t91270;
    wire t91272 = t91271 ^ t91271;
    wire t91273 = t91272 ^ t91272;
    wire t91274 = t91273 ^ t91273;
    wire t91275 = t91274 ^ t91274;
    wire t91276 = t91275 ^ t91275;
    wire t91277 = t91276 ^ t91276;
    wire t91278 = t91277 ^ t91277;
    wire t91279 = t91278 ^ t91278;
    wire t91280 = t91279 ^ t91279;
    wire t91281 = t91280 ^ t91280;
    wire t91282 = t91281 ^ t91281;
    wire t91283 = t91282 ^ t91282;
    wire t91284 = t91283 ^ t91283;
    wire t91285 = t91284 ^ t91284;
    wire t91286 = t91285 ^ t91285;
    wire t91287 = t91286 ^ t91286;
    wire t91288 = t91287 ^ t91287;
    wire t91289 = t91288 ^ t91288;
    wire t91290 = t91289 ^ t91289;
    wire t91291 = t91290 ^ t91290;
    wire t91292 = t91291 ^ t91291;
    wire t91293 = t91292 ^ t91292;
    wire t91294 = t91293 ^ t91293;
    wire t91295 = t91294 ^ t91294;
    wire t91296 = t91295 ^ t91295;
    wire t91297 = t91296 ^ t91296;
    wire t91298 = t91297 ^ t91297;
    wire t91299 = t91298 ^ t91298;
    wire t91300 = t91299 ^ t91299;
    wire t91301 = t91300 ^ t91300;
    wire t91302 = t91301 ^ t91301;
    wire t91303 = t91302 ^ t91302;
    wire t91304 = t91303 ^ t91303;
    wire t91305 = t91304 ^ t91304;
    wire t91306 = t91305 ^ t91305;
    wire t91307 = t91306 ^ t91306;
    wire t91308 = t91307 ^ t91307;
    wire t91309 = t91308 ^ t91308;
    wire t91310 = t91309 ^ t91309;
    wire t91311 = t91310 ^ t91310;
    wire t91312 = t91311 ^ t91311;
    wire t91313 = t91312 ^ t91312;
    wire t91314 = t91313 ^ t91313;
    wire t91315 = t91314 ^ t91314;
    wire t91316 = t91315 ^ t91315;
    wire t91317 = t91316 ^ t91316;
    wire t91318 = t91317 ^ t91317;
    wire t91319 = t91318 ^ t91318;
    wire t91320 = t91319 ^ t91319;
    wire t91321 = t91320 ^ t91320;
    wire t91322 = t91321 ^ t91321;
    wire t91323 = t91322 ^ t91322;
    wire t91324 = t91323 ^ t91323;
    wire t91325 = t91324 ^ t91324;
    wire t91326 = t91325 ^ t91325;
    wire t91327 = t91326 ^ t91326;
    wire t91328 = t91327 ^ t91327;
    wire t91329 = t91328 ^ t91328;
    wire t91330 = t91329 ^ t91329;
    wire t91331 = t91330 ^ t91330;
    wire t91332 = t91331 ^ t91331;
    wire t91333 = t91332 ^ t91332;
    wire t91334 = t91333 ^ t91333;
    wire t91335 = t91334 ^ t91334;
    wire t91336 = t91335 ^ t91335;
    wire t91337 = t91336 ^ t91336;
    wire t91338 = t91337 ^ t91337;
    wire t91339 = t91338 ^ t91338;
    wire t91340 = t91339 ^ t91339;
    wire t91341 = t91340 ^ t91340;
    wire t91342 = t91341 ^ t91341;
    wire t91343 = t91342 ^ t91342;
    wire t91344 = t91343 ^ t91343;
    wire t91345 = t91344 ^ t91344;
    wire t91346 = t91345 ^ t91345;
    wire t91347 = t91346 ^ t91346;
    wire t91348 = t91347 ^ t91347;
    wire t91349 = t91348 ^ t91348;
    wire t91350 = t91349 ^ t91349;
    wire t91351 = t91350 ^ t91350;
    wire t91352 = t91351 ^ t91351;
    wire t91353 = t91352 ^ t91352;
    wire t91354 = t91353 ^ t91353;
    wire t91355 = t91354 ^ t91354;
    wire t91356 = t91355 ^ t91355;
    wire t91357 = t91356 ^ t91356;
    wire t91358 = t91357 ^ t91357;
    wire t91359 = t91358 ^ t91358;
    wire t91360 = t91359 ^ t91359;
    wire t91361 = t91360 ^ t91360;
    wire t91362 = t91361 ^ t91361;
    wire t91363 = t91362 ^ t91362;
    wire t91364 = t91363 ^ t91363;
    wire t91365 = t91364 ^ t91364;
    wire t91366 = t91365 ^ t91365;
    wire t91367 = t91366 ^ t91366;
    wire t91368 = t91367 ^ t91367;
    wire t91369 = t91368 ^ t91368;
    wire t91370 = t91369 ^ t91369;
    wire t91371 = t91370 ^ t91370;
    wire t91372 = t91371 ^ t91371;
    wire t91373 = t91372 ^ t91372;
    wire t91374 = t91373 ^ t91373;
    wire t91375 = t91374 ^ t91374;
    wire t91376 = t91375 ^ t91375;
    wire t91377 = t91376 ^ t91376;
    wire t91378 = t91377 ^ t91377;
    wire t91379 = t91378 ^ t91378;
    wire t91380 = t91379 ^ t91379;
    wire t91381 = t91380 ^ t91380;
    wire t91382 = t91381 ^ t91381;
    wire t91383 = t91382 ^ t91382;
    wire t91384 = t91383 ^ t91383;
    wire t91385 = t91384 ^ t91384;
    wire t91386 = t91385 ^ t91385;
    wire t91387 = t91386 ^ t91386;
    wire t91388 = t91387 ^ t91387;
    wire t91389 = t91388 ^ t91388;
    wire t91390 = t91389 ^ t91389;
    wire t91391 = t91390 ^ t91390;
    wire t91392 = t91391 ^ t91391;
    wire t91393 = t91392 ^ t91392;
    wire t91394 = t91393 ^ t91393;
    wire t91395 = t91394 ^ t91394;
    wire t91396 = t91395 ^ t91395;
    wire t91397 = t91396 ^ t91396;
    wire t91398 = t91397 ^ t91397;
    wire t91399 = t91398 ^ t91398;
    wire t91400 = t91399 ^ t91399;
    wire t91401 = t91400 ^ t91400;
    wire t91402 = t91401 ^ t91401;
    wire t91403 = t91402 ^ t91402;
    wire t91404 = t91403 ^ t91403;
    wire t91405 = t91404 ^ t91404;
    wire t91406 = t91405 ^ t91405;
    wire t91407 = t91406 ^ t91406;
    wire t91408 = t91407 ^ t91407;
    wire t91409 = t91408 ^ t91408;
    wire t91410 = t91409 ^ t91409;
    wire t91411 = t91410 ^ t91410;
    wire t91412 = t91411 ^ t91411;
    wire t91413 = t91412 ^ t91412;
    wire t91414 = t91413 ^ t91413;
    wire t91415 = t91414 ^ t91414;
    wire t91416 = t91415 ^ t91415;
    wire t91417 = t91416 ^ t91416;
    wire t91418 = t91417 ^ t91417;
    wire t91419 = t91418 ^ t91418;
    wire t91420 = t91419 ^ t91419;
    wire t91421 = t91420 ^ t91420;
    wire t91422 = t91421 ^ t91421;
    wire t91423 = t91422 ^ t91422;
    wire t91424 = t91423 ^ t91423;
    wire t91425 = t91424 ^ t91424;
    wire t91426 = t91425 ^ t91425;
    wire t91427 = t91426 ^ t91426;
    wire t91428 = t91427 ^ t91427;
    wire t91429 = t91428 ^ t91428;
    wire t91430 = t91429 ^ t91429;
    wire t91431 = t91430 ^ t91430;
    wire t91432 = t91431 ^ t91431;
    wire t91433 = t91432 ^ t91432;
    wire t91434 = t91433 ^ t91433;
    wire t91435 = t91434 ^ t91434;
    wire t91436 = t91435 ^ t91435;
    wire t91437 = t91436 ^ t91436;
    wire t91438 = t91437 ^ t91437;
    wire t91439 = t91438 ^ t91438;
    wire t91440 = t91439 ^ t91439;
    wire t91441 = t91440 ^ t91440;
    wire t91442 = t91441 ^ t91441;
    wire t91443 = t91442 ^ t91442;
    wire t91444 = t91443 ^ t91443;
    wire t91445 = t91444 ^ t91444;
    wire t91446 = t91445 ^ t91445;
    wire t91447 = t91446 ^ t91446;
    wire t91448 = t91447 ^ t91447;
    wire t91449 = t91448 ^ t91448;
    wire t91450 = t91449 ^ t91449;
    wire t91451 = t91450 ^ t91450;
    wire t91452 = t91451 ^ t91451;
    wire t91453 = t91452 ^ t91452;
    wire t91454 = t91453 ^ t91453;
    wire t91455 = t91454 ^ t91454;
    wire t91456 = t91455 ^ t91455;
    wire t91457 = t91456 ^ t91456;
    wire t91458 = t91457 ^ t91457;
    wire t91459 = t91458 ^ t91458;
    wire t91460 = t91459 ^ t91459;
    wire t91461 = t91460 ^ t91460;
    wire t91462 = t91461 ^ t91461;
    wire t91463 = t91462 ^ t91462;
    wire t91464 = t91463 ^ t91463;
    wire t91465 = t91464 ^ t91464;
    wire t91466 = t91465 ^ t91465;
    wire t91467 = t91466 ^ t91466;
    wire t91468 = t91467 ^ t91467;
    wire t91469 = t91468 ^ t91468;
    wire t91470 = t91469 ^ t91469;
    wire t91471 = t91470 ^ t91470;
    wire t91472 = t91471 ^ t91471;
    wire t91473 = t91472 ^ t91472;
    wire t91474 = t91473 ^ t91473;
    wire t91475 = t91474 ^ t91474;
    wire t91476 = t91475 ^ t91475;
    wire t91477 = t91476 ^ t91476;
    wire t91478 = t91477 ^ t91477;
    wire t91479 = t91478 ^ t91478;
    wire t91480 = t91479 ^ t91479;
    wire t91481 = t91480 ^ t91480;
    wire t91482 = t91481 ^ t91481;
    wire t91483 = t91482 ^ t91482;
    wire t91484 = t91483 ^ t91483;
    wire t91485 = t91484 ^ t91484;
    wire t91486 = t91485 ^ t91485;
    wire t91487 = t91486 ^ t91486;
    wire t91488 = t91487 ^ t91487;
    wire t91489 = t91488 ^ t91488;
    wire t91490 = t91489 ^ t91489;
    wire t91491 = t91490 ^ t91490;
    wire t91492 = t91491 ^ t91491;
    wire t91493 = t91492 ^ t91492;
    wire t91494 = t91493 ^ t91493;
    wire t91495 = t91494 ^ t91494;
    wire t91496 = t91495 ^ t91495;
    wire t91497 = t91496 ^ t91496;
    wire t91498 = t91497 ^ t91497;
    wire t91499 = t91498 ^ t91498;
    wire t91500 = t91499 ^ t91499;
    wire t91501 = t91500 ^ t91500;
    wire t91502 = t91501 ^ t91501;
    wire t91503 = t91502 ^ t91502;
    wire t91504 = t91503 ^ t91503;
    wire t91505 = t91504 ^ t91504;
    wire t91506 = t91505 ^ t91505;
    wire t91507 = t91506 ^ t91506;
    wire t91508 = t91507 ^ t91507;
    wire t91509 = t91508 ^ t91508;
    wire t91510 = t91509 ^ t91509;
    wire t91511 = t91510 ^ t91510;
    wire t91512 = t91511 ^ t91511;
    wire t91513 = t91512 ^ t91512;
    wire t91514 = t91513 ^ t91513;
    wire t91515 = t91514 ^ t91514;
    wire t91516 = t91515 ^ t91515;
    wire t91517 = t91516 ^ t91516;
    wire t91518 = t91517 ^ t91517;
    wire t91519 = t91518 ^ t91518;
    wire t91520 = t91519 ^ t91519;
    wire t91521 = t91520 ^ t91520;
    wire t91522 = t91521 ^ t91521;
    wire t91523 = t91522 ^ t91522;
    wire t91524 = t91523 ^ t91523;
    wire t91525 = t91524 ^ t91524;
    wire t91526 = t91525 ^ t91525;
    wire t91527 = t91526 ^ t91526;
    wire t91528 = t91527 ^ t91527;
    wire t91529 = t91528 ^ t91528;
    wire t91530 = t91529 ^ t91529;
    wire t91531 = t91530 ^ t91530;
    wire t91532 = t91531 ^ t91531;
    wire t91533 = t91532 ^ t91532;
    wire t91534 = t91533 ^ t91533;
    wire t91535 = t91534 ^ t91534;
    wire t91536 = t91535 ^ t91535;
    wire t91537 = t91536 ^ t91536;
    wire t91538 = t91537 ^ t91537;
    wire t91539 = t91538 ^ t91538;
    wire t91540 = t91539 ^ t91539;
    wire t91541 = t91540 ^ t91540;
    wire t91542 = t91541 ^ t91541;
    wire t91543 = t91542 ^ t91542;
    wire t91544 = t91543 ^ t91543;
    wire t91545 = t91544 ^ t91544;
    wire t91546 = t91545 ^ t91545;
    wire t91547 = t91546 ^ t91546;
    wire t91548 = t91547 ^ t91547;
    wire t91549 = t91548 ^ t91548;
    wire t91550 = t91549 ^ t91549;
    wire t91551 = t91550 ^ t91550;
    wire t91552 = t91551 ^ t91551;
    wire t91553 = t91552 ^ t91552;
    wire t91554 = t91553 ^ t91553;
    wire t91555 = t91554 ^ t91554;
    wire t91556 = t91555 ^ t91555;
    wire t91557 = t91556 ^ t91556;
    wire t91558 = t91557 ^ t91557;
    wire t91559 = t91558 ^ t91558;
    wire t91560 = t91559 ^ t91559;
    wire t91561 = t91560 ^ t91560;
    wire t91562 = t91561 ^ t91561;
    wire t91563 = t91562 ^ t91562;
    wire t91564 = t91563 ^ t91563;
    wire t91565 = t91564 ^ t91564;
    wire t91566 = t91565 ^ t91565;
    wire t91567 = t91566 ^ t91566;
    wire t91568 = t91567 ^ t91567;
    wire t91569 = t91568 ^ t91568;
    wire t91570 = t91569 ^ t91569;
    wire t91571 = t91570 ^ t91570;
    wire t91572 = t91571 ^ t91571;
    wire t91573 = t91572 ^ t91572;
    wire t91574 = t91573 ^ t91573;
    wire t91575 = t91574 ^ t91574;
    wire t91576 = t91575 ^ t91575;
    wire t91577 = t91576 ^ t91576;
    wire t91578 = t91577 ^ t91577;
    wire t91579 = t91578 ^ t91578;
    wire t91580 = t91579 ^ t91579;
    wire t91581 = t91580 ^ t91580;
    wire t91582 = t91581 ^ t91581;
    wire t91583 = t91582 ^ t91582;
    wire t91584 = t91583 ^ t91583;
    wire t91585 = t91584 ^ t91584;
    wire t91586 = t91585 ^ t91585;
    wire t91587 = t91586 ^ t91586;
    wire t91588 = t91587 ^ t91587;
    wire t91589 = t91588 ^ t91588;
    wire t91590 = t91589 ^ t91589;
    wire t91591 = t91590 ^ t91590;
    wire t91592 = t91591 ^ t91591;
    wire t91593 = t91592 ^ t91592;
    wire t91594 = t91593 ^ t91593;
    wire t91595 = t91594 ^ t91594;
    wire t91596 = t91595 ^ t91595;
    wire t91597 = t91596 ^ t91596;
    wire t91598 = t91597 ^ t91597;
    wire t91599 = t91598 ^ t91598;
    wire t91600 = t91599 ^ t91599;
    wire t91601 = t91600 ^ t91600;
    wire t91602 = t91601 ^ t91601;
    wire t91603 = t91602 ^ t91602;
    wire t91604 = t91603 ^ t91603;
    wire t91605 = t91604 ^ t91604;
    wire t91606 = t91605 ^ t91605;
    wire t91607 = t91606 ^ t91606;
    wire t91608 = t91607 ^ t91607;
    wire t91609 = t91608 ^ t91608;
    wire t91610 = t91609 ^ t91609;
    wire t91611 = t91610 ^ t91610;
    wire t91612 = t91611 ^ t91611;
    wire t91613 = t91612 ^ t91612;
    wire t91614 = t91613 ^ t91613;
    wire t91615 = t91614 ^ t91614;
    wire t91616 = t91615 ^ t91615;
    wire t91617 = t91616 ^ t91616;
    wire t91618 = t91617 ^ t91617;
    wire t91619 = t91618 ^ t91618;
    wire t91620 = t91619 ^ t91619;
    wire t91621 = t91620 ^ t91620;
    wire t91622 = t91621 ^ t91621;
    wire t91623 = t91622 ^ t91622;
    wire t91624 = t91623 ^ t91623;
    wire t91625 = t91624 ^ t91624;
    wire t91626 = t91625 ^ t91625;
    wire t91627 = t91626 ^ t91626;
    wire t91628 = t91627 ^ t91627;
    wire t91629 = t91628 ^ t91628;
    wire t91630 = t91629 ^ t91629;
    wire t91631 = t91630 ^ t91630;
    wire t91632 = t91631 ^ t91631;
    wire t91633 = t91632 ^ t91632;
    wire t91634 = t91633 ^ t91633;
    wire t91635 = t91634 ^ t91634;
    wire t91636 = t91635 ^ t91635;
    wire t91637 = t91636 ^ t91636;
    wire t91638 = t91637 ^ t91637;
    wire t91639 = t91638 ^ t91638;
    wire t91640 = t91639 ^ t91639;
    wire t91641 = t91640 ^ t91640;
    wire t91642 = t91641 ^ t91641;
    wire t91643 = t91642 ^ t91642;
    wire t91644 = t91643 ^ t91643;
    wire t91645 = t91644 ^ t91644;
    wire t91646 = t91645 ^ t91645;
    wire t91647 = t91646 ^ t91646;
    wire t91648 = t91647 ^ t91647;
    wire t91649 = t91648 ^ t91648;
    wire t91650 = t91649 ^ t91649;
    wire t91651 = t91650 ^ t91650;
    wire t91652 = t91651 ^ t91651;
    wire t91653 = t91652 ^ t91652;
    wire t91654 = t91653 ^ t91653;
    wire t91655 = t91654 ^ t91654;
    wire t91656 = t91655 ^ t91655;
    wire t91657 = t91656 ^ t91656;
    wire t91658 = t91657 ^ t91657;
    wire t91659 = t91658 ^ t91658;
    wire t91660 = t91659 ^ t91659;
    wire t91661 = t91660 ^ t91660;
    wire t91662 = t91661 ^ t91661;
    wire t91663 = t91662 ^ t91662;
    wire t91664 = t91663 ^ t91663;
    wire t91665 = t91664 ^ t91664;
    wire t91666 = t91665 ^ t91665;
    wire t91667 = t91666 ^ t91666;
    wire t91668 = t91667 ^ t91667;
    wire t91669 = t91668 ^ t91668;
    wire t91670 = t91669 ^ t91669;
    wire t91671 = t91670 ^ t91670;
    wire t91672 = t91671 ^ t91671;
    wire t91673 = t91672 ^ t91672;
    wire t91674 = t91673 ^ t91673;
    wire t91675 = t91674 ^ t91674;
    wire t91676 = t91675 ^ t91675;
    wire t91677 = t91676 ^ t91676;
    wire t91678 = t91677 ^ t91677;
    wire t91679 = t91678 ^ t91678;
    wire t91680 = t91679 ^ t91679;
    wire t91681 = t91680 ^ t91680;
    wire t91682 = t91681 ^ t91681;
    wire t91683 = t91682 ^ t91682;
    wire t91684 = t91683 ^ t91683;
    wire t91685 = t91684 ^ t91684;
    wire t91686 = t91685 ^ t91685;
    wire t91687 = t91686 ^ t91686;
    wire t91688 = t91687 ^ t91687;
    wire t91689 = t91688 ^ t91688;
    wire t91690 = t91689 ^ t91689;
    wire t91691 = t91690 ^ t91690;
    wire t91692 = t91691 ^ t91691;
    wire t91693 = t91692 ^ t91692;
    wire t91694 = t91693 ^ t91693;
    wire t91695 = t91694 ^ t91694;
    wire t91696 = t91695 ^ t91695;
    wire t91697 = t91696 ^ t91696;
    wire t91698 = t91697 ^ t91697;
    wire t91699 = t91698 ^ t91698;
    wire t91700 = t91699 ^ t91699;
    wire t91701 = t91700 ^ t91700;
    wire t91702 = t91701 ^ t91701;
    wire t91703 = t91702 ^ t91702;
    wire t91704 = t91703 ^ t91703;
    wire t91705 = t91704 ^ t91704;
    wire t91706 = t91705 ^ t91705;
    wire t91707 = t91706 ^ t91706;
    wire t91708 = t91707 ^ t91707;
    wire t91709 = t91708 ^ t91708;
    wire t91710 = t91709 ^ t91709;
    wire t91711 = t91710 ^ t91710;
    wire t91712 = t91711 ^ t91711;
    wire t91713 = t91712 ^ t91712;
    wire t91714 = t91713 ^ t91713;
    wire t91715 = t91714 ^ t91714;
    wire t91716 = t91715 ^ t91715;
    wire t91717 = t91716 ^ t91716;
    wire t91718 = t91717 ^ t91717;
    wire t91719 = t91718 ^ t91718;
    wire t91720 = t91719 ^ t91719;
    wire t91721 = t91720 ^ t91720;
    wire t91722 = t91721 ^ t91721;
    wire t91723 = t91722 ^ t91722;
    wire t91724 = t91723 ^ t91723;
    wire t91725 = t91724 ^ t91724;
    wire t91726 = t91725 ^ t91725;
    wire t91727 = t91726 ^ t91726;
    wire t91728 = t91727 ^ t91727;
    wire t91729 = t91728 ^ t91728;
    wire t91730 = t91729 ^ t91729;
    wire t91731 = t91730 ^ t91730;
    wire t91732 = t91731 ^ t91731;
    wire t91733 = t91732 ^ t91732;
    wire t91734 = t91733 ^ t91733;
    wire t91735 = t91734 ^ t91734;
    wire t91736 = t91735 ^ t91735;
    wire t91737 = t91736 ^ t91736;
    wire t91738 = t91737 ^ t91737;
    wire t91739 = t91738 ^ t91738;
    wire t91740 = t91739 ^ t91739;
    wire t91741 = t91740 ^ t91740;
    wire t91742 = t91741 ^ t91741;
    wire t91743 = t91742 ^ t91742;
    wire t91744 = t91743 ^ t91743;
    wire t91745 = t91744 ^ t91744;
    wire t91746 = t91745 ^ t91745;
    wire t91747 = t91746 ^ t91746;
    wire t91748 = t91747 ^ t91747;
    wire t91749 = t91748 ^ t91748;
    wire t91750 = t91749 ^ t91749;
    wire t91751 = t91750 ^ t91750;
    wire t91752 = t91751 ^ t91751;
    wire t91753 = t91752 ^ t91752;
    wire t91754 = t91753 ^ t91753;
    wire t91755 = t91754 ^ t91754;
    wire t91756 = t91755 ^ t91755;
    wire t91757 = t91756 ^ t91756;
    wire t91758 = t91757 ^ t91757;
    wire t91759 = t91758 ^ t91758;
    wire t91760 = t91759 ^ t91759;
    wire t91761 = t91760 ^ t91760;
    wire t91762 = t91761 ^ t91761;
    wire t91763 = t91762 ^ t91762;
    wire t91764 = t91763 ^ t91763;
    wire t91765 = t91764 ^ t91764;
    wire t91766 = t91765 ^ t91765;
    wire t91767 = t91766 ^ t91766;
    wire t91768 = t91767 ^ t91767;
    wire t91769 = t91768 ^ t91768;
    wire t91770 = t91769 ^ t91769;
    wire t91771 = t91770 ^ t91770;
    wire t91772 = t91771 ^ t91771;
    wire t91773 = t91772 ^ t91772;
    wire t91774 = t91773 ^ t91773;
    wire t91775 = t91774 ^ t91774;
    wire t91776 = t91775 ^ t91775;
    wire t91777 = t91776 ^ t91776;
    wire t91778 = t91777 ^ t91777;
    wire t91779 = t91778 ^ t91778;
    wire t91780 = t91779 ^ t91779;
    wire t91781 = t91780 ^ t91780;
    wire t91782 = t91781 ^ t91781;
    wire t91783 = t91782 ^ t91782;
    wire t91784 = t91783 ^ t91783;
    wire t91785 = t91784 ^ t91784;
    wire t91786 = t91785 ^ t91785;
    wire t91787 = t91786 ^ t91786;
    wire t91788 = t91787 ^ t91787;
    wire t91789 = t91788 ^ t91788;
    wire t91790 = t91789 ^ t91789;
    wire t91791 = t91790 ^ t91790;
    wire t91792 = t91791 ^ t91791;
    wire t91793 = t91792 ^ t91792;
    wire t91794 = t91793 ^ t91793;
    wire t91795 = t91794 ^ t91794;
    wire t91796 = t91795 ^ t91795;
    wire t91797 = t91796 ^ t91796;
    wire t91798 = t91797 ^ t91797;
    wire t91799 = t91798 ^ t91798;
    wire t91800 = t91799 ^ t91799;
    wire t91801 = t91800 ^ t91800;
    wire t91802 = t91801 ^ t91801;
    wire t91803 = t91802 ^ t91802;
    wire t91804 = t91803 ^ t91803;
    wire t91805 = t91804 ^ t91804;
    wire t91806 = t91805 ^ t91805;
    wire t91807 = t91806 ^ t91806;
    wire t91808 = t91807 ^ t91807;
    wire t91809 = t91808 ^ t91808;
    wire t91810 = t91809 ^ t91809;
    wire t91811 = t91810 ^ t91810;
    wire t91812 = t91811 ^ t91811;
    wire t91813 = t91812 ^ t91812;
    wire t91814 = t91813 ^ t91813;
    wire t91815 = t91814 ^ t91814;
    wire t91816 = t91815 ^ t91815;
    wire t91817 = t91816 ^ t91816;
    wire t91818 = t91817 ^ t91817;
    wire t91819 = t91818 ^ t91818;
    wire t91820 = t91819 ^ t91819;
    wire t91821 = t91820 ^ t91820;
    wire t91822 = t91821 ^ t91821;
    wire t91823 = t91822 ^ t91822;
    wire t91824 = t91823 ^ t91823;
    wire t91825 = t91824 ^ t91824;
    wire t91826 = t91825 ^ t91825;
    wire t91827 = t91826 ^ t91826;
    wire t91828 = t91827 ^ t91827;
    wire t91829 = t91828 ^ t91828;
    wire t91830 = t91829 ^ t91829;
    wire t91831 = t91830 ^ t91830;
    wire t91832 = t91831 ^ t91831;
    wire t91833 = t91832 ^ t91832;
    wire t91834 = t91833 ^ t91833;
    wire t91835 = t91834 ^ t91834;
    wire t91836 = t91835 ^ t91835;
    wire t91837 = t91836 ^ t91836;
    wire t91838 = t91837 ^ t91837;
    wire t91839 = t91838 ^ t91838;
    wire t91840 = t91839 ^ t91839;
    wire t91841 = t91840 ^ t91840;
    wire t91842 = t91841 ^ t91841;
    wire t91843 = t91842 ^ t91842;
    wire t91844 = t91843 ^ t91843;
    wire t91845 = t91844 ^ t91844;
    wire t91846 = t91845 ^ t91845;
    wire t91847 = t91846 ^ t91846;
    wire t91848 = t91847 ^ t91847;
    wire t91849 = t91848 ^ t91848;
    wire t91850 = t91849 ^ t91849;
    wire t91851 = t91850 ^ t91850;
    wire t91852 = t91851 ^ t91851;
    wire t91853 = t91852 ^ t91852;
    wire t91854 = t91853 ^ t91853;
    wire t91855 = t91854 ^ t91854;
    wire t91856 = t91855 ^ t91855;
    wire t91857 = t91856 ^ t91856;
    wire t91858 = t91857 ^ t91857;
    wire t91859 = t91858 ^ t91858;
    wire t91860 = t91859 ^ t91859;
    wire t91861 = t91860 ^ t91860;
    wire t91862 = t91861 ^ t91861;
    wire t91863 = t91862 ^ t91862;
    wire t91864 = t91863 ^ t91863;
    wire t91865 = t91864 ^ t91864;
    wire t91866 = t91865 ^ t91865;
    wire t91867 = t91866 ^ t91866;
    wire t91868 = t91867 ^ t91867;
    wire t91869 = t91868 ^ t91868;
    wire t91870 = t91869 ^ t91869;
    wire t91871 = t91870 ^ t91870;
    wire t91872 = t91871 ^ t91871;
    wire t91873 = t91872 ^ t91872;
    wire t91874 = t91873 ^ t91873;
    wire t91875 = t91874 ^ t91874;
    wire t91876 = t91875 ^ t91875;
    wire t91877 = t91876 ^ t91876;
    wire t91878 = t91877 ^ t91877;
    wire t91879 = t91878 ^ t91878;
    wire t91880 = t91879 ^ t91879;
    wire t91881 = t91880 ^ t91880;
    wire t91882 = t91881 ^ t91881;
    wire t91883 = t91882 ^ t91882;
    wire t91884 = t91883 ^ t91883;
    wire t91885 = t91884 ^ t91884;
    wire t91886 = t91885 ^ t91885;
    wire t91887 = t91886 ^ t91886;
    wire t91888 = t91887 ^ t91887;
    wire t91889 = t91888 ^ t91888;
    wire t91890 = t91889 ^ t91889;
    wire t91891 = t91890 ^ t91890;
    wire t91892 = t91891 ^ t91891;
    wire t91893 = t91892 ^ t91892;
    wire t91894 = t91893 ^ t91893;
    wire t91895 = t91894 ^ t91894;
    wire t91896 = t91895 ^ t91895;
    wire t91897 = t91896 ^ t91896;
    wire t91898 = t91897 ^ t91897;
    wire t91899 = t91898 ^ t91898;
    wire t91900 = t91899 ^ t91899;
    wire t91901 = t91900 ^ t91900;
    wire t91902 = t91901 ^ t91901;
    wire t91903 = t91902 ^ t91902;
    wire t91904 = t91903 ^ t91903;
    wire t91905 = t91904 ^ t91904;
    wire t91906 = t91905 ^ t91905;
    wire t91907 = t91906 ^ t91906;
    wire t91908 = t91907 ^ t91907;
    wire t91909 = t91908 ^ t91908;
    wire t91910 = t91909 ^ t91909;
    wire t91911 = t91910 ^ t91910;
    wire t91912 = t91911 ^ t91911;
    wire t91913 = t91912 ^ t91912;
    wire t91914 = t91913 ^ t91913;
    wire t91915 = t91914 ^ t91914;
    wire t91916 = t91915 ^ t91915;
    wire t91917 = t91916 ^ t91916;
    wire t91918 = t91917 ^ t91917;
    wire t91919 = t91918 ^ t91918;
    wire t91920 = t91919 ^ t91919;
    wire t91921 = t91920 ^ t91920;
    wire t91922 = t91921 ^ t91921;
    wire t91923 = t91922 ^ t91922;
    wire t91924 = t91923 ^ t91923;
    wire t91925 = t91924 ^ t91924;
    wire t91926 = t91925 ^ t91925;
    wire t91927 = t91926 ^ t91926;
    wire t91928 = t91927 ^ t91927;
    wire t91929 = t91928 ^ t91928;
    wire t91930 = t91929 ^ t91929;
    wire t91931 = t91930 ^ t91930;
    wire t91932 = t91931 ^ t91931;
    wire t91933 = t91932 ^ t91932;
    wire t91934 = t91933 ^ t91933;
    wire t91935 = t91934 ^ t91934;
    wire t91936 = t91935 ^ t91935;
    wire t91937 = t91936 ^ t91936;
    wire t91938 = t91937 ^ t91937;
    wire t91939 = t91938 ^ t91938;
    wire t91940 = t91939 ^ t91939;
    wire t91941 = t91940 ^ t91940;
    wire t91942 = t91941 ^ t91941;
    wire t91943 = t91942 ^ t91942;
    wire t91944 = t91943 ^ t91943;
    wire t91945 = t91944 ^ t91944;
    wire t91946 = t91945 ^ t91945;
    wire t91947 = t91946 ^ t91946;
    wire t91948 = t91947 ^ t91947;
    wire t91949 = t91948 ^ t91948;
    wire t91950 = t91949 ^ t91949;
    wire t91951 = t91950 ^ t91950;
    wire t91952 = t91951 ^ t91951;
    wire t91953 = t91952 ^ t91952;
    wire t91954 = t91953 ^ t91953;
    wire t91955 = t91954 ^ t91954;
    wire t91956 = t91955 ^ t91955;
    wire t91957 = t91956 ^ t91956;
    wire t91958 = t91957 ^ t91957;
    wire t91959 = t91958 ^ t91958;
    wire t91960 = t91959 ^ t91959;
    wire t91961 = t91960 ^ t91960;
    wire t91962 = t91961 ^ t91961;
    wire t91963 = t91962 ^ t91962;
    wire t91964 = t91963 ^ t91963;
    wire t91965 = t91964 ^ t91964;
    wire t91966 = t91965 ^ t91965;
    wire t91967 = t91966 ^ t91966;
    wire t91968 = t91967 ^ t91967;
    wire t91969 = t91968 ^ t91968;
    wire t91970 = t91969 ^ t91969;
    wire t91971 = t91970 ^ t91970;
    wire t91972 = t91971 ^ t91971;
    wire t91973 = t91972 ^ t91972;
    wire t91974 = t91973 ^ t91973;
    wire t91975 = t91974 ^ t91974;
    wire t91976 = t91975 ^ t91975;
    wire t91977 = t91976 ^ t91976;
    wire t91978 = t91977 ^ t91977;
    wire t91979 = t91978 ^ t91978;
    wire t91980 = t91979 ^ t91979;
    wire t91981 = t91980 ^ t91980;
    wire t91982 = t91981 ^ t91981;
    wire t91983 = t91982 ^ t91982;
    wire t91984 = t91983 ^ t91983;
    wire t91985 = t91984 ^ t91984;
    wire t91986 = t91985 ^ t91985;
    wire t91987 = t91986 ^ t91986;
    wire t91988 = t91987 ^ t91987;
    wire t91989 = t91988 ^ t91988;
    wire t91990 = t91989 ^ t91989;
    wire t91991 = t91990 ^ t91990;
    wire t91992 = t91991 ^ t91991;
    wire t91993 = t91992 ^ t91992;
    wire t91994 = t91993 ^ t91993;
    wire t91995 = t91994 ^ t91994;
    wire t91996 = t91995 ^ t91995;
    wire t91997 = t91996 ^ t91996;
    wire t91998 = t91997 ^ t91997;
    wire t91999 = t91998 ^ t91998;
    wire t92000 = t91999 ^ t91999;
    wire t92001 = t92000 ^ t92000;
    wire t92002 = t92001 ^ t92001;
    wire t92003 = t92002 ^ t92002;
    wire t92004 = t92003 ^ t92003;
    wire t92005 = t92004 ^ t92004;
    wire t92006 = t92005 ^ t92005;
    wire t92007 = t92006 ^ t92006;
    wire t92008 = t92007 ^ t92007;
    wire t92009 = t92008 ^ t92008;
    wire t92010 = t92009 ^ t92009;
    wire t92011 = t92010 ^ t92010;
    wire t92012 = t92011 ^ t92011;
    wire t92013 = t92012 ^ t92012;
    wire t92014 = t92013 ^ t92013;
    wire t92015 = t92014 ^ t92014;
    wire t92016 = t92015 ^ t92015;
    wire t92017 = t92016 ^ t92016;
    wire t92018 = t92017 ^ t92017;
    wire t92019 = t92018 ^ t92018;
    wire t92020 = t92019 ^ t92019;
    wire t92021 = t92020 ^ t92020;
    wire t92022 = t92021 ^ t92021;
    wire t92023 = t92022 ^ t92022;
    wire t92024 = t92023 ^ t92023;
    wire t92025 = t92024 ^ t92024;
    wire t92026 = t92025 ^ t92025;
    wire t92027 = t92026 ^ t92026;
    wire t92028 = t92027 ^ t92027;
    wire t92029 = t92028 ^ t92028;
    wire t92030 = t92029 ^ t92029;
    wire t92031 = t92030 ^ t92030;
    wire t92032 = t92031 ^ t92031;
    wire t92033 = t92032 ^ t92032;
    wire t92034 = t92033 ^ t92033;
    wire t92035 = t92034 ^ t92034;
    wire t92036 = t92035 ^ t92035;
    wire t92037 = t92036 ^ t92036;
    wire t92038 = t92037 ^ t92037;
    wire t92039 = t92038 ^ t92038;
    wire t92040 = t92039 ^ t92039;
    wire t92041 = t92040 ^ t92040;
    wire t92042 = t92041 ^ t92041;
    wire t92043 = t92042 ^ t92042;
    wire t92044 = t92043 ^ t92043;
    wire t92045 = t92044 ^ t92044;
    wire t92046 = t92045 ^ t92045;
    wire t92047 = t92046 ^ t92046;
    wire t92048 = t92047 ^ t92047;
    wire t92049 = t92048 ^ t92048;
    wire t92050 = t92049 ^ t92049;
    wire t92051 = t92050 ^ t92050;
    wire t92052 = t92051 ^ t92051;
    wire t92053 = t92052 ^ t92052;
    wire t92054 = t92053 ^ t92053;
    wire t92055 = t92054 ^ t92054;
    wire t92056 = t92055 ^ t92055;
    wire t92057 = t92056 ^ t92056;
    wire t92058 = t92057 ^ t92057;
    wire t92059 = t92058 ^ t92058;
    wire t92060 = t92059 ^ t92059;
    wire t92061 = t92060 ^ t92060;
    wire t92062 = t92061 ^ t92061;
    wire t92063 = t92062 ^ t92062;
    wire t92064 = t92063 ^ t92063;
    wire t92065 = t92064 ^ t92064;
    wire t92066 = t92065 ^ t92065;
    wire t92067 = t92066 ^ t92066;
    wire t92068 = t92067 ^ t92067;
    wire t92069 = t92068 ^ t92068;
    wire t92070 = t92069 ^ t92069;
    wire t92071 = t92070 ^ t92070;
    wire t92072 = t92071 ^ t92071;
    wire t92073 = t92072 ^ t92072;
    wire t92074 = t92073 ^ t92073;
    wire t92075 = t92074 ^ t92074;
    wire t92076 = t92075 ^ t92075;
    wire t92077 = t92076 ^ t92076;
    wire t92078 = t92077 ^ t92077;
    wire t92079 = t92078 ^ t92078;
    wire t92080 = t92079 ^ t92079;
    wire t92081 = t92080 ^ t92080;
    wire t92082 = t92081 ^ t92081;
    wire t92083 = t92082 ^ t92082;
    wire t92084 = t92083 ^ t92083;
    wire t92085 = t92084 ^ t92084;
    wire t92086 = t92085 ^ t92085;
    wire t92087 = t92086 ^ t92086;
    wire t92088 = t92087 ^ t92087;
    wire t92089 = t92088 ^ t92088;
    wire t92090 = t92089 ^ t92089;
    wire t92091 = t92090 ^ t92090;
    wire t92092 = t92091 ^ t92091;
    wire t92093 = t92092 ^ t92092;
    wire t92094 = t92093 ^ t92093;
    wire t92095 = t92094 ^ t92094;
    wire t92096 = t92095 ^ t92095;
    wire t92097 = t92096 ^ t92096;
    wire t92098 = t92097 ^ t92097;
    wire t92099 = t92098 ^ t92098;
    wire t92100 = t92099 ^ t92099;
    wire t92101 = t92100 ^ t92100;
    wire t92102 = t92101 ^ t92101;
    wire t92103 = t92102 ^ t92102;
    wire t92104 = t92103 ^ t92103;
    wire t92105 = t92104 ^ t92104;
    wire t92106 = t92105 ^ t92105;
    wire t92107 = t92106 ^ t92106;
    wire t92108 = t92107 ^ t92107;
    wire t92109 = t92108 ^ t92108;
    wire t92110 = t92109 ^ t92109;
    wire t92111 = t92110 ^ t92110;
    wire t92112 = t92111 ^ t92111;
    wire t92113 = t92112 ^ t92112;
    wire t92114 = t92113 ^ t92113;
    wire t92115 = t92114 ^ t92114;
    wire t92116 = t92115 ^ t92115;
    wire t92117 = t92116 ^ t92116;
    wire t92118 = t92117 ^ t92117;
    wire t92119 = t92118 ^ t92118;
    wire t92120 = t92119 ^ t92119;
    wire t92121 = t92120 ^ t92120;
    wire t92122 = t92121 ^ t92121;
    wire t92123 = t92122 ^ t92122;
    wire t92124 = t92123 ^ t92123;
    wire t92125 = t92124 ^ t92124;
    wire t92126 = t92125 ^ t92125;
    wire t92127 = t92126 ^ t92126;
    wire t92128 = t92127 ^ t92127;
    wire t92129 = t92128 ^ t92128;
    wire t92130 = t92129 ^ t92129;
    wire t92131 = t92130 ^ t92130;
    wire t92132 = t92131 ^ t92131;
    wire t92133 = t92132 ^ t92132;
    wire t92134 = t92133 ^ t92133;
    wire t92135 = t92134 ^ t92134;
    wire t92136 = t92135 ^ t92135;
    wire t92137 = t92136 ^ t92136;
    wire t92138 = t92137 ^ t92137;
    wire t92139 = t92138 ^ t92138;
    wire t92140 = t92139 ^ t92139;
    wire t92141 = t92140 ^ t92140;
    wire t92142 = t92141 ^ t92141;
    wire t92143 = t92142 ^ t92142;
    wire t92144 = t92143 ^ t92143;
    wire t92145 = t92144 ^ t92144;
    wire t92146 = t92145 ^ t92145;
    wire t92147 = t92146 ^ t92146;
    wire t92148 = t92147 ^ t92147;
    wire t92149 = t92148 ^ t92148;
    wire t92150 = t92149 ^ t92149;
    wire t92151 = t92150 ^ t92150;
    wire t92152 = t92151 ^ t92151;
    wire t92153 = t92152 ^ t92152;
    wire t92154 = t92153 ^ t92153;
    wire t92155 = t92154 ^ t92154;
    wire t92156 = t92155 ^ t92155;
    wire t92157 = t92156 ^ t92156;
    wire t92158 = t92157 ^ t92157;
    wire t92159 = t92158 ^ t92158;
    wire t92160 = t92159 ^ t92159;
    wire t92161 = t92160 ^ t92160;
    wire t92162 = t92161 ^ t92161;
    wire t92163 = t92162 ^ t92162;
    wire t92164 = t92163 ^ t92163;
    wire t92165 = t92164 ^ t92164;
    wire t92166 = t92165 ^ t92165;
    wire t92167 = t92166 ^ t92166;
    wire t92168 = t92167 ^ t92167;
    wire t92169 = t92168 ^ t92168;
    wire t92170 = t92169 ^ t92169;
    wire t92171 = t92170 ^ t92170;
    wire t92172 = t92171 ^ t92171;
    wire t92173 = t92172 ^ t92172;
    wire t92174 = t92173 ^ t92173;
    wire t92175 = t92174 ^ t92174;
    wire t92176 = t92175 ^ t92175;
    wire t92177 = t92176 ^ t92176;
    wire t92178 = t92177 ^ t92177;
    wire t92179 = t92178 ^ t92178;
    wire t92180 = t92179 ^ t92179;
    wire t92181 = t92180 ^ t92180;
    wire t92182 = t92181 ^ t92181;
    wire t92183 = t92182 ^ t92182;
    wire t92184 = t92183 ^ t92183;
    wire t92185 = t92184 ^ t92184;
    wire t92186 = t92185 ^ t92185;
    wire t92187 = t92186 ^ t92186;
    wire t92188 = t92187 ^ t92187;
    wire t92189 = t92188 ^ t92188;
    wire t92190 = t92189 ^ t92189;
    wire t92191 = t92190 ^ t92190;
    wire t92192 = t92191 ^ t92191;
    wire t92193 = t92192 ^ t92192;
    wire t92194 = t92193 ^ t92193;
    wire t92195 = t92194 ^ t92194;
    wire t92196 = t92195 ^ t92195;
    wire t92197 = t92196 ^ t92196;
    wire t92198 = t92197 ^ t92197;
    wire t92199 = t92198 ^ t92198;
    wire t92200 = t92199 ^ t92199;
    wire t92201 = t92200 ^ t92200;
    wire t92202 = t92201 ^ t92201;
    wire t92203 = t92202 ^ t92202;
    wire t92204 = t92203 ^ t92203;
    wire t92205 = t92204 ^ t92204;
    wire t92206 = t92205 ^ t92205;
    wire t92207 = t92206 ^ t92206;
    wire t92208 = t92207 ^ t92207;
    wire t92209 = t92208 ^ t92208;
    wire t92210 = t92209 ^ t92209;
    wire t92211 = t92210 ^ t92210;
    wire t92212 = t92211 ^ t92211;
    wire t92213 = t92212 ^ t92212;
    wire t92214 = t92213 ^ t92213;
    wire t92215 = t92214 ^ t92214;
    wire t92216 = t92215 ^ t92215;
    wire t92217 = t92216 ^ t92216;
    wire t92218 = t92217 ^ t92217;
    wire t92219 = t92218 ^ t92218;
    wire t92220 = t92219 ^ t92219;
    wire t92221 = t92220 ^ t92220;
    wire t92222 = t92221 ^ t92221;
    wire t92223 = t92222 ^ t92222;
    wire t92224 = t92223 ^ t92223;
    wire t92225 = t92224 ^ t92224;
    wire t92226 = t92225 ^ t92225;
    wire t92227 = t92226 ^ t92226;
    wire t92228 = t92227 ^ t92227;
    wire t92229 = t92228 ^ t92228;
    wire t92230 = t92229 ^ t92229;
    wire t92231 = t92230 ^ t92230;
    wire t92232 = t92231 ^ t92231;
    wire t92233 = t92232 ^ t92232;
    wire t92234 = t92233 ^ t92233;
    wire t92235 = t92234 ^ t92234;
    wire t92236 = t92235 ^ t92235;
    wire t92237 = t92236 ^ t92236;
    wire t92238 = t92237 ^ t92237;
    wire t92239 = t92238 ^ t92238;
    wire t92240 = t92239 ^ t92239;
    wire t92241 = t92240 ^ t92240;
    wire t92242 = t92241 ^ t92241;
    wire t92243 = t92242 ^ t92242;
    wire t92244 = t92243 ^ t92243;
    wire t92245 = t92244 ^ t92244;
    wire t92246 = t92245 ^ t92245;
    wire t92247 = t92246 ^ t92246;
    wire t92248 = t92247 ^ t92247;
    wire t92249 = t92248 ^ t92248;
    wire t92250 = t92249 ^ t92249;
    wire t92251 = t92250 ^ t92250;
    wire t92252 = t92251 ^ t92251;
    wire t92253 = t92252 ^ t92252;
    wire t92254 = t92253 ^ t92253;
    wire t92255 = t92254 ^ t92254;
    wire t92256 = t92255 ^ t92255;
    wire t92257 = t92256 ^ t92256;
    wire t92258 = t92257 ^ t92257;
    wire t92259 = t92258 ^ t92258;
    wire t92260 = t92259 ^ t92259;
    wire t92261 = t92260 ^ t92260;
    wire t92262 = t92261 ^ t92261;
    wire t92263 = t92262 ^ t92262;
    wire t92264 = t92263 ^ t92263;
    wire t92265 = t92264 ^ t92264;
    wire t92266 = t92265 ^ t92265;
    wire t92267 = t92266 ^ t92266;
    wire t92268 = t92267 ^ t92267;
    wire t92269 = t92268 ^ t92268;
    wire t92270 = t92269 ^ t92269;
    wire t92271 = t92270 ^ t92270;
    wire t92272 = t92271 ^ t92271;
    wire t92273 = t92272 ^ t92272;
    wire t92274 = t92273 ^ t92273;
    wire t92275 = t92274 ^ t92274;
    wire t92276 = t92275 ^ t92275;
    wire t92277 = t92276 ^ t92276;
    wire t92278 = t92277 ^ t92277;
    wire t92279 = t92278 ^ t92278;
    wire t92280 = t92279 ^ t92279;
    wire t92281 = t92280 ^ t92280;
    wire t92282 = t92281 ^ t92281;
    wire t92283 = t92282 ^ t92282;
    wire t92284 = t92283 ^ t92283;
    wire t92285 = t92284 ^ t92284;
    wire t92286 = t92285 ^ t92285;
    wire t92287 = t92286 ^ t92286;
    wire t92288 = t92287 ^ t92287;
    wire t92289 = t92288 ^ t92288;
    wire t92290 = t92289 ^ t92289;
    wire t92291 = t92290 ^ t92290;
    wire t92292 = t92291 ^ t92291;
    wire t92293 = t92292 ^ t92292;
    wire t92294 = t92293 ^ t92293;
    wire t92295 = t92294 ^ t92294;
    wire t92296 = t92295 ^ t92295;
    wire t92297 = t92296 ^ t92296;
    wire t92298 = t92297 ^ t92297;
    wire t92299 = t92298 ^ t92298;
    wire t92300 = t92299 ^ t92299;
    wire t92301 = t92300 ^ t92300;
    wire t92302 = t92301 ^ t92301;
    wire t92303 = t92302 ^ t92302;
    wire t92304 = t92303 ^ t92303;
    wire t92305 = t92304 ^ t92304;
    wire t92306 = t92305 ^ t92305;
    wire t92307 = t92306 ^ t92306;
    wire t92308 = t92307 ^ t92307;
    wire t92309 = t92308 ^ t92308;
    wire t92310 = t92309 ^ t92309;
    wire t92311 = t92310 ^ t92310;
    wire t92312 = t92311 ^ t92311;
    wire t92313 = t92312 ^ t92312;
    wire t92314 = t92313 ^ t92313;
    wire t92315 = t92314 ^ t92314;
    wire t92316 = t92315 ^ t92315;
    wire t92317 = t92316 ^ t92316;
    wire t92318 = t92317 ^ t92317;
    wire t92319 = t92318 ^ t92318;
    wire t92320 = t92319 ^ t92319;
    wire t92321 = t92320 ^ t92320;
    wire t92322 = t92321 ^ t92321;
    wire t92323 = t92322 ^ t92322;
    wire t92324 = t92323 ^ t92323;
    wire t92325 = t92324 ^ t92324;
    wire t92326 = t92325 ^ t92325;
    wire t92327 = t92326 ^ t92326;
    wire t92328 = t92327 ^ t92327;
    wire t92329 = t92328 ^ t92328;
    wire t92330 = t92329 ^ t92329;
    wire t92331 = t92330 ^ t92330;
    wire t92332 = t92331 ^ t92331;
    wire t92333 = t92332 ^ t92332;
    wire t92334 = t92333 ^ t92333;
    wire t92335 = t92334 ^ t92334;
    wire t92336 = t92335 ^ t92335;
    wire t92337 = t92336 ^ t92336;
    wire t92338 = t92337 ^ t92337;
    wire t92339 = t92338 ^ t92338;
    wire t92340 = t92339 ^ t92339;
    wire t92341 = t92340 ^ t92340;
    wire t92342 = t92341 ^ t92341;
    wire t92343 = t92342 ^ t92342;
    wire t92344 = t92343 ^ t92343;
    wire t92345 = t92344 ^ t92344;
    wire t92346 = t92345 ^ t92345;
    wire t92347 = t92346 ^ t92346;
    wire t92348 = t92347 ^ t92347;
    wire t92349 = t92348 ^ t92348;
    wire t92350 = t92349 ^ t92349;
    wire t92351 = t92350 ^ t92350;
    wire t92352 = t92351 ^ t92351;
    wire t92353 = t92352 ^ t92352;
    wire t92354 = t92353 ^ t92353;
    wire t92355 = t92354 ^ t92354;
    wire t92356 = t92355 ^ t92355;
    wire t92357 = t92356 ^ t92356;
    wire t92358 = t92357 ^ t92357;
    wire t92359 = t92358 ^ t92358;
    wire t92360 = t92359 ^ t92359;
    wire t92361 = t92360 ^ t92360;
    wire t92362 = t92361 ^ t92361;
    wire t92363 = t92362 ^ t92362;
    wire t92364 = t92363 ^ t92363;
    wire t92365 = t92364 ^ t92364;
    wire t92366 = t92365 ^ t92365;
    wire t92367 = t92366 ^ t92366;
    wire t92368 = t92367 ^ t92367;
    wire t92369 = t92368 ^ t92368;
    wire t92370 = t92369 ^ t92369;
    wire t92371 = t92370 ^ t92370;
    wire t92372 = t92371 ^ t92371;
    wire t92373 = t92372 ^ t92372;
    wire t92374 = t92373 ^ t92373;
    wire t92375 = t92374 ^ t92374;
    wire t92376 = t92375 ^ t92375;
    wire t92377 = t92376 ^ t92376;
    wire t92378 = t92377 ^ t92377;
    wire t92379 = t92378 ^ t92378;
    wire t92380 = t92379 ^ t92379;
    wire t92381 = t92380 ^ t92380;
    wire t92382 = t92381 ^ t92381;
    wire t92383 = t92382 ^ t92382;
    wire t92384 = t92383 ^ t92383;
    wire t92385 = t92384 ^ t92384;
    wire t92386 = t92385 ^ t92385;
    wire t92387 = t92386 ^ t92386;
    wire t92388 = t92387 ^ t92387;
    wire t92389 = t92388 ^ t92388;
    wire t92390 = t92389 ^ t92389;
    wire t92391 = t92390 ^ t92390;
    wire t92392 = t92391 ^ t92391;
    wire t92393 = t92392 ^ t92392;
    wire t92394 = t92393 ^ t92393;
    wire t92395 = t92394 ^ t92394;
    wire t92396 = t92395 ^ t92395;
    wire t92397 = t92396 ^ t92396;
    wire t92398 = t92397 ^ t92397;
    wire t92399 = t92398 ^ t92398;
    wire t92400 = t92399 ^ t92399;
    wire t92401 = t92400 ^ t92400;
    wire t92402 = t92401 ^ t92401;
    wire t92403 = t92402 ^ t92402;
    wire t92404 = t92403 ^ t92403;
    wire t92405 = t92404 ^ t92404;
    wire t92406 = t92405 ^ t92405;
    wire t92407 = t92406 ^ t92406;
    wire t92408 = t92407 ^ t92407;
    wire t92409 = t92408 ^ t92408;
    wire t92410 = t92409 ^ t92409;
    wire t92411 = t92410 ^ t92410;
    wire t92412 = t92411 ^ t92411;
    wire t92413 = t92412 ^ t92412;
    wire t92414 = t92413 ^ t92413;
    wire t92415 = t92414 ^ t92414;
    wire t92416 = t92415 ^ t92415;
    wire t92417 = t92416 ^ t92416;
    wire t92418 = t92417 ^ t92417;
    wire t92419 = t92418 ^ t92418;
    wire t92420 = t92419 ^ t92419;
    wire t92421 = t92420 ^ t92420;
    wire t92422 = t92421 ^ t92421;
    wire t92423 = t92422 ^ t92422;
    wire t92424 = t92423 ^ t92423;
    wire t92425 = t92424 ^ t92424;
    wire t92426 = t92425 ^ t92425;
    wire t92427 = t92426 ^ t92426;
    wire t92428 = t92427 ^ t92427;
    wire t92429 = t92428 ^ t92428;
    wire t92430 = t92429 ^ t92429;
    wire t92431 = t92430 ^ t92430;
    wire t92432 = t92431 ^ t92431;
    wire t92433 = t92432 ^ t92432;
    wire t92434 = t92433 ^ t92433;
    wire t92435 = t92434 ^ t92434;
    wire t92436 = t92435 ^ t92435;
    wire t92437 = t92436 ^ t92436;
    wire t92438 = t92437 ^ t92437;
    wire t92439 = t92438 ^ t92438;
    wire t92440 = t92439 ^ t92439;
    wire t92441 = t92440 ^ t92440;
    wire t92442 = t92441 ^ t92441;
    wire t92443 = t92442 ^ t92442;
    wire t92444 = t92443 ^ t92443;
    wire t92445 = t92444 ^ t92444;
    wire t92446 = t92445 ^ t92445;
    wire t92447 = t92446 ^ t92446;
    wire t92448 = t92447 ^ t92447;
    wire t92449 = t92448 ^ t92448;
    wire t92450 = t92449 ^ t92449;
    wire t92451 = t92450 ^ t92450;
    wire t92452 = t92451 ^ t92451;
    wire t92453 = t92452 ^ t92452;
    wire t92454 = t92453 ^ t92453;
    wire t92455 = t92454 ^ t92454;
    wire t92456 = t92455 ^ t92455;
    wire t92457 = t92456 ^ t92456;
    wire t92458 = t92457 ^ t92457;
    wire t92459 = t92458 ^ t92458;
    wire t92460 = t92459 ^ t92459;
    wire t92461 = t92460 ^ t92460;
    wire t92462 = t92461 ^ t92461;
    wire t92463 = t92462 ^ t92462;
    wire t92464 = t92463 ^ t92463;
    wire t92465 = t92464 ^ t92464;
    wire t92466 = t92465 ^ t92465;
    wire t92467 = t92466 ^ t92466;
    wire t92468 = t92467 ^ t92467;
    wire t92469 = t92468 ^ t92468;
    wire t92470 = t92469 ^ t92469;
    wire t92471 = t92470 ^ t92470;
    wire t92472 = t92471 ^ t92471;
    wire t92473 = t92472 ^ t92472;
    wire t92474 = t92473 ^ t92473;
    wire t92475 = t92474 ^ t92474;
    wire t92476 = t92475 ^ t92475;
    wire t92477 = t92476 ^ t92476;
    wire t92478 = t92477 ^ t92477;
    wire t92479 = t92478 ^ t92478;
    wire t92480 = t92479 ^ t92479;
    wire t92481 = t92480 ^ t92480;
    wire t92482 = t92481 ^ t92481;
    wire t92483 = t92482 ^ t92482;
    wire t92484 = t92483 ^ t92483;
    wire t92485 = t92484 ^ t92484;
    wire t92486 = t92485 ^ t92485;
    wire t92487 = t92486 ^ t92486;
    wire t92488 = t92487 ^ t92487;
    wire t92489 = t92488 ^ t92488;
    wire t92490 = t92489 ^ t92489;
    wire t92491 = t92490 ^ t92490;
    wire t92492 = t92491 ^ t92491;
    wire t92493 = t92492 ^ t92492;
    wire t92494 = t92493 ^ t92493;
    wire t92495 = t92494 ^ t92494;
    wire t92496 = t92495 ^ t92495;
    wire t92497 = t92496 ^ t92496;
    wire t92498 = t92497 ^ t92497;
    wire t92499 = t92498 ^ t92498;
    wire t92500 = t92499 ^ t92499;
    wire t92501 = t92500 ^ t92500;
    wire t92502 = t92501 ^ t92501;
    wire t92503 = t92502 ^ t92502;
    wire t92504 = t92503 ^ t92503;
    wire t92505 = t92504 ^ t92504;
    wire t92506 = t92505 ^ t92505;
    wire t92507 = t92506 ^ t92506;
    wire t92508 = t92507 ^ t92507;
    wire t92509 = t92508 ^ t92508;
    wire t92510 = t92509 ^ t92509;
    wire t92511 = t92510 ^ t92510;
    wire t92512 = t92511 ^ t92511;
    wire t92513 = t92512 ^ t92512;
    wire t92514 = t92513 ^ t92513;
    wire t92515 = t92514 ^ t92514;
    wire t92516 = t92515 ^ t92515;
    wire t92517 = t92516 ^ t92516;
    wire t92518 = t92517 ^ t92517;
    wire t92519 = t92518 ^ t92518;
    wire t92520 = t92519 ^ t92519;
    wire t92521 = t92520 ^ t92520;
    wire t92522 = t92521 ^ t92521;
    wire t92523 = t92522 ^ t92522;
    wire t92524 = t92523 ^ t92523;
    wire t92525 = t92524 ^ t92524;
    wire t92526 = t92525 ^ t92525;
    wire t92527 = t92526 ^ t92526;
    wire t92528 = t92527 ^ t92527;
    wire t92529 = t92528 ^ t92528;
    wire t92530 = t92529 ^ t92529;
    wire t92531 = t92530 ^ t92530;
    wire t92532 = t92531 ^ t92531;
    wire t92533 = t92532 ^ t92532;
    wire t92534 = t92533 ^ t92533;
    wire t92535 = t92534 ^ t92534;
    wire t92536 = t92535 ^ t92535;
    wire t92537 = t92536 ^ t92536;
    wire t92538 = t92537 ^ t92537;
    wire t92539 = t92538 ^ t92538;
    wire t92540 = t92539 ^ t92539;
    wire t92541 = t92540 ^ t92540;
    wire t92542 = t92541 ^ t92541;
    wire t92543 = t92542 ^ t92542;
    wire t92544 = t92543 ^ t92543;
    wire t92545 = t92544 ^ t92544;
    wire t92546 = t92545 ^ t92545;
    wire t92547 = t92546 ^ t92546;
    wire t92548 = t92547 ^ t92547;
    wire t92549 = t92548 ^ t92548;
    wire t92550 = t92549 ^ t92549;
    wire t92551 = t92550 ^ t92550;
    wire t92552 = t92551 ^ t92551;
    wire t92553 = t92552 ^ t92552;
    wire t92554 = t92553 ^ t92553;
    wire t92555 = t92554 ^ t92554;
    wire t92556 = t92555 ^ t92555;
    wire t92557 = t92556 ^ t92556;
    wire t92558 = t92557 ^ t92557;
    wire t92559 = t92558 ^ t92558;
    wire t92560 = t92559 ^ t92559;
    wire t92561 = t92560 ^ t92560;
    wire t92562 = t92561 ^ t92561;
    wire t92563 = t92562 ^ t92562;
    wire t92564 = t92563 ^ t92563;
    wire t92565 = t92564 ^ t92564;
    wire t92566 = t92565 ^ t92565;
    wire t92567 = t92566 ^ t92566;
    wire t92568 = t92567 ^ t92567;
    wire t92569 = t92568 ^ t92568;
    wire t92570 = t92569 ^ t92569;
    wire t92571 = t92570 ^ t92570;
    wire t92572 = t92571 ^ t92571;
    wire t92573 = t92572 ^ t92572;
    wire t92574 = t92573 ^ t92573;
    wire t92575 = t92574 ^ t92574;
    wire t92576 = t92575 ^ t92575;
    wire t92577 = t92576 ^ t92576;
    wire t92578 = t92577 ^ t92577;
    wire t92579 = t92578 ^ t92578;
    wire t92580 = t92579 ^ t92579;
    wire t92581 = t92580 ^ t92580;
    wire t92582 = t92581 ^ t92581;
    wire t92583 = t92582 ^ t92582;
    wire t92584 = t92583 ^ t92583;
    wire t92585 = t92584 ^ t92584;
    wire t92586 = t92585 ^ t92585;
    wire t92587 = t92586 ^ t92586;
    wire t92588 = t92587 ^ t92587;
    wire t92589 = t92588 ^ t92588;
    wire t92590 = t92589 ^ t92589;
    wire t92591 = t92590 ^ t92590;
    wire t92592 = t92591 ^ t92591;
    wire t92593 = t92592 ^ t92592;
    wire t92594 = t92593 ^ t92593;
    wire t92595 = t92594 ^ t92594;
    wire t92596 = t92595 ^ t92595;
    wire t92597 = t92596 ^ t92596;
    wire t92598 = t92597 ^ t92597;
    wire t92599 = t92598 ^ t92598;
    wire t92600 = t92599 ^ t92599;
    wire t92601 = t92600 ^ t92600;
    wire t92602 = t92601 ^ t92601;
    wire t92603 = t92602 ^ t92602;
    wire t92604 = t92603 ^ t92603;
    wire t92605 = t92604 ^ t92604;
    wire t92606 = t92605 ^ t92605;
    wire t92607 = t92606 ^ t92606;
    wire t92608 = t92607 ^ t92607;
    wire t92609 = t92608 ^ t92608;
    wire t92610 = t92609 ^ t92609;
    wire t92611 = t92610 ^ t92610;
    wire t92612 = t92611 ^ t92611;
    wire t92613 = t92612 ^ t92612;
    wire t92614 = t92613 ^ t92613;
    wire t92615 = t92614 ^ t92614;
    wire t92616 = t92615 ^ t92615;
    wire t92617 = t92616 ^ t92616;
    wire t92618 = t92617 ^ t92617;
    wire t92619 = t92618 ^ t92618;
    wire t92620 = t92619 ^ t92619;
    wire t92621 = t92620 ^ t92620;
    wire t92622 = t92621 ^ t92621;
    wire t92623 = t92622 ^ t92622;
    wire t92624 = t92623 ^ t92623;
    wire t92625 = t92624 ^ t92624;
    wire t92626 = t92625 ^ t92625;
    wire t92627 = t92626 ^ t92626;
    wire t92628 = t92627 ^ t92627;
    wire t92629 = t92628 ^ t92628;
    wire t92630 = t92629 ^ t92629;
    wire t92631 = t92630 ^ t92630;
    wire t92632 = t92631 ^ t92631;
    wire t92633 = t92632 ^ t92632;
    wire t92634 = t92633 ^ t92633;
    wire t92635 = t92634 ^ t92634;
    wire t92636 = t92635 ^ t92635;
    wire t92637 = t92636 ^ t92636;
    wire t92638 = t92637 ^ t92637;
    wire t92639 = t92638 ^ t92638;
    wire t92640 = t92639 ^ t92639;
    wire t92641 = t92640 ^ t92640;
    wire t92642 = t92641 ^ t92641;
    wire t92643 = t92642 ^ t92642;
    wire t92644 = t92643 ^ t92643;
    wire t92645 = t92644 ^ t92644;
    wire t92646 = t92645 ^ t92645;
    wire t92647 = t92646 ^ t92646;
    wire t92648 = t92647 ^ t92647;
    wire t92649 = t92648 ^ t92648;
    wire t92650 = t92649 ^ t92649;
    wire t92651 = t92650 ^ t92650;
    wire t92652 = t92651 ^ t92651;
    wire t92653 = t92652 ^ t92652;
    wire t92654 = t92653 ^ t92653;
    wire t92655 = t92654 ^ t92654;
    wire t92656 = t92655 ^ t92655;
    wire t92657 = t92656 ^ t92656;
    wire t92658 = t92657 ^ t92657;
    wire t92659 = t92658 ^ t92658;
    wire t92660 = t92659 ^ t92659;
    wire t92661 = t92660 ^ t92660;
    wire t92662 = t92661 ^ t92661;
    wire t92663 = t92662 ^ t92662;
    wire t92664 = t92663 ^ t92663;
    wire t92665 = t92664 ^ t92664;
    wire t92666 = t92665 ^ t92665;
    wire t92667 = t92666 ^ t92666;
    wire t92668 = t92667 ^ t92667;
    wire t92669 = t92668 ^ t92668;
    wire t92670 = t92669 ^ t92669;
    wire t92671 = t92670 ^ t92670;
    wire t92672 = t92671 ^ t92671;
    wire t92673 = t92672 ^ t92672;
    wire t92674 = t92673 ^ t92673;
    wire t92675 = t92674 ^ t92674;
    wire t92676 = t92675 ^ t92675;
    wire t92677 = t92676 ^ t92676;
    wire t92678 = t92677 ^ t92677;
    wire t92679 = t92678 ^ t92678;
    wire t92680 = t92679 ^ t92679;
    wire t92681 = t92680 ^ t92680;
    wire t92682 = t92681 ^ t92681;
    wire t92683 = t92682 ^ t92682;
    wire t92684 = t92683 ^ t92683;
    wire t92685 = t92684 ^ t92684;
    wire t92686 = t92685 ^ t92685;
    wire t92687 = t92686 ^ t92686;
    wire t92688 = t92687 ^ t92687;
    wire t92689 = t92688 ^ t92688;
    wire t92690 = t92689 ^ t92689;
    wire t92691 = t92690 ^ t92690;
    wire t92692 = t92691 ^ t92691;
    wire t92693 = t92692 ^ t92692;
    wire t92694 = t92693 ^ t92693;
    wire t92695 = t92694 ^ t92694;
    wire t92696 = t92695 ^ t92695;
    wire t92697 = t92696 ^ t92696;
    wire t92698 = t92697 ^ t92697;
    wire t92699 = t92698 ^ t92698;
    wire t92700 = t92699 ^ t92699;
    wire t92701 = t92700 ^ t92700;
    wire t92702 = t92701 ^ t92701;
    wire t92703 = t92702 ^ t92702;
    wire t92704 = t92703 ^ t92703;
    wire t92705 = t92704 ^ t92704;
    wire t92706 = t92705 ^ t92705;
    wire t92707 = t92706 ^ t92706;
    wire t92708 = t92707 ^ t92707;
    wire t92709 = t92708 ^ t92708;
    wire t92710 = t92709 ^ t92709;
    wire t92711 = t92710 ^ t92710;
    wire t92712 = t92711 ^ t92711;
    wire t92713 = t92712 ^ t92712;
    wire t92714 = t92713 ^ t92713;
    wire t92715 = t92714 ^ t92714;
    wire t92716 = t92715 ^ t92715;
    wire t92717 = t92716 ^ t92716;
    wire t92718 = t92717 ^ t92717;
    wire t92719 = t92718 ^ t92718;
    wire t92720 = t92719 ^ t92719;
    wire t92721 = t92720 ^ t92720;
    wire t92722 = t92721 ^ t92721;
    wire t92723 = t92722 ^ t92722;
    wire t92724 = t92723 ^ t92723;
    wire t92725 = t92724 ^ t92724;
    wire t92726 = t92725 ^ t92725;
    wire t92727 = t92726 ^ t92726;
    wire t92728 = t92727 ^ t92727;
    wire t92729 = t92728 ^ t92728;
    wire t92730 = t92729 ^ t92729;
    wire t92731 = t92730 ^ t92730;
    wire t92732 = t92731 ^ t92731;
    wire t92733 = t92732 ^ t92732;
    wire t92734 = t92733 ^ t92733;
    wire t92735 = t92734 ^ t92734;
    wire t92736 = t92735 ^ t92735;
    wire t92737 = t92736 ^ t92736;
    wire t92738 = t92737 ^ t92737;
    wire t92739 = t92738 ^ t92738;
    wire t92740 = t92739 ^ t92739;
    wire t92741 = t92740 ^ t92740;
    wire t92742 = t92741 ^ t92741;
    wire t92743 = t92742 ^ t92742;
    wire t92744 = t92743 ^ t92743;
    wire t92745 = t92744 ^ t92744;
    wire t92746 = t92745 ^ t92745;
    wire t92747 = t92746 ^ t92746;
    wire t92748 = t92747 ^ t92747;
    wire t92749 = t92748 ^ t92748;
    wire t92750 = t92749 ^ t92749;
    wire t92751 = t92750 ^ t92750;
    wire t92752 = t92751 ^ t92751;
    wire t92753 = t92752 ^ t92752;
    wire t92754 = t92753 ^ t92753;
    wire t92755 = t92754 ^ t92754;
    wire t92756 = t92755 ^ t92755;
    wire t92757 = t92756 ^ t92756;
    wire t92758 = t92757 ^ t92757;
    wire t92759 = t92758 ^ t92758;
    wire t92760 = t92759 ^ t92759;
    wire t92761 = t92760 ^ t92760;
    wire t92762 = t92761 ^ t92761;
    wire t92763 = t92762 ^ t92762;
    wire t92764 = t92763 ^ t92763;
    wire t92765 = t92764 ^ t92764;
    wire t92766 = t92765 ^ t92765;
    wire t92767 = t92766 ^ t92766;
    wire t92768 = t92767 ^ t92767;
    wire t92769 = t92768 ^ t92768;
    wire t92770 = t92769 ^ t92769;
    wire t92771 = t92770 ^ t92770;
    wire t92772 = t92771 ^ t92771;
    wire t92773 = t92772 ^ t92772;
    wire t92774 = t92773 ^ t92773;
    wire t92775 = t92774 ^ t92774;
    wire t92776 = t92775 ^ t92775;
    wire t92777 = t92776 ^ t92776;
    wire t92778 = t92777 ^ t92777;
    wire t92779 = t92778 ^ t92778;
    wire t92780 = t92779 ^ t92779;
    wire t92781 = t92780 ^ t92780;
    wire t92782 = t92781 ^ t92781;
    wire t92783 = t92782 ^ t92782;
    wire t92784 = t92783 ^ t92783;
    wire t92785 = t92784 ^ t92784;
    wire t92786 = t92785 ^ t92785;
    wire t92787 = t92786 ^ t92786;
    wire t92788 = t92787 ^ t92787;
    wire t92789 = t92788 ^ t92788;
    wire t92790 = t92789 ^ t92789;
    wire t92791 = t92790 ^ t92790;
    wire t92792 = t92791 ^ t92791;
    wire t92793 = t92792 ^ t92792;
    wire t92794 = t92793 ^ t92793;
    wire t92795 = t92794 ^ t92794;
    wire t92796 = t92795 ^ t92795;
    wire t92797 = t92796 ^ t92796;
    wire t92798 = t92797 ^ t92797;
    wire t92799 = t92798 ^ t92798;
    wire t92800 = t92799 ^ t92799;
    wire t92801 = t92800 ^ t92800;
    wire t92802 = t92801 ^ t92801;
    wire t92803 = t92802 ^ t92802;
    wire t92804 = t92803 ^ t92803;
    wire t92805 = t92804 ^ t92804;
    wire t92806 = t92805 ^ t92805;
    wire t92807 = t92806 ^ t92806;
    wire t92808 = t92807 ^ t92807;
    wire t92809 = t92808 ^ t92808;
    wire t92810 = t92809 ^ t92809;
    wire t92811 = t92810 ^ t92810;
    wire t92812 = t92811 ^ t92811;
    wire t92813 = t92812 ^ t92812;
    wire t92814 = t92813 ^ t92813;
    wire t92815 = t92814 ^ t92814;
    wire t92816 = t92815 ^ t92815;
    wire t92817 = t92816 ^ t92816;
    wire t92818 = t92817 ^ t92817;
    wire t92819 = t92818 ^ t92818;
    wire t92820 = t92819 ^ t92819;
    wire t92821 = t92820 ^ t92820;
    wire t92822 = t92821 ^ t92821;
    wire t92823 = t92822 ^ t92822;
    wire t92824 = t92823 ^ t92823;
    wire t92825 = t92824 ^ t92824;
    wire t92826 = t92825 ^ t92825;
    wire t92827 = t92826 ^ t92826;
    wire t92828 = t92827 ^ t92827;
    wire t92829 = t92828 ^ t92828;
    wire t92830 = t92829 ^ t92829;
    wire t92831 = t92830 ^ t92830;
    wire t92832 = t92831 ^ t92831;
    wire t92833 = t92832 ^ t92832;
    wire t92834 = t92833 ^ t92833;
    wire t92835 = t92834 ^ t92834;
    wire t92836 = t92835 ^ t92835;
    wire t92837 = t92836 ^ t92836;
    wire t92838 = t92837 ^ t92837;
    wire t92839 = t92838 ^ t92838;
    wire t92840 = t92839 ^ t92839;
    wire t92841 = t92840 ^ t92840;
    wire t92842 = t92841 ^ t92841;
    wire t92843 = t92842 ^ t92842;
    wire t92844 = t92843 ^ t92843;
    wire t92845 = t92844 ^ t92844;
    wire t92846 = t92845 ^ t92845;
    wire t92847 = t92846 ^ t92846;
    wire t92848 = t92847 ^ t92847;
    wire t92849 = t92848 ^ t92848;
    wire t92850 = t92849 ^ t92849;
    wire t92851 = t92850 ^ t92850;
    wire t92852 = t92851 ^ t92851;
    wire t92853 = t92852 ^ t92852;
    wire t92854 = t92853 ^ t92853;
    wire t92855 = t92854 ^ t92854;
    wire t92856 = t92855 ^ t92855;
    wire t92857 = t92856 ^ t92856;
    wire t92858 = t92857 ^ t92857;
    wire t92859 = t92858 ^ t92858;
    wire t92860 = t92859 ^ t92859;
    wire t92861 = t92860 ^ t92860;
    wire t92862 = t92861 ^ t92861;
    wire t92863 = t92862 ^ t92862;
    wire t92864 = t92863 ^ t92863;
    wire t92865 = t92864 ^ t92864;
    wire t92866 = t92865 ^ t92865;
    wire t92867 = t92866 ^ t92866;
    wire t92868 = t92867 ^ t92867;
    wire t92869 = t92868 ^ t92868;
    wire t92870 = t92869 ^ t92869;
    wire t92871 = t92870 ^ t92870;
    wire t92872 = t92871 ^ t92871;
    wire t92873 = t92872 ^ t92872;
    wire t92874 = t92873 ^ t92873;
    wire t92875 = t92874 ^ t92874;
    wire t92876 = t92875 ^ t92875;
    wire t92877 = t92876 ^ t92876;
    wire t92878 = t92877 ^ t92877;
    wire t92879 = t92878 ^ t92878;
    wire t92880 = t92879 ^ t92879;
    wire t92881 = t92880 ^ t92880;
    wire t92882 = t92881 ^ t92881;
    wire t92883 = t92882 ^ t92882;
    wire t92884 = t92883 ^ t92883;
    wire t92885 = t92884 ^ t92884;
    wire t92886 = t92885 ^ t92885;
    wire t92887 = t92886 ^ t92886;
    wire t92888 = t92887 ^ t92887;
    wire t92889 = t92888 ^ t92888;
    wire t92890 = t92889 ^ t92889;
    wire t92891 = t92890 ^ t92890;
    wire t92892 = t92891 ^ t92891;
    wire t92893 = t92892 ^ t92892;
    wire t92894 = t92893 ^ t92893;
    wire t92895 = t92894 ^ t92894;
    wire t92896 = t92895 ^ t92895;
    wire t92897 = t92896 ^ t92896;
    wire t92898 = t92897 ^ t92897;
    wire t92899 = t92898 ^ t92898;
    wire t92900 = t92899 ^ t92899;
    wire t92901 = t92900 ^ t92900;
    wire t92902 = t92901 ^ t92901;
    wire t92903 = t92902 ^ t92902;
    wire t92904 = t92903 ^ t92903;
    wire t92905 = t92904 ^ t92904;
    wire t92906 = t92905 ^ t92905;
    wire t92907 = t92906 ^ t92906;
    wire t92908 = t92907 ^ t92907;
    wire t92909 = t92908 ^ t92908;
    wire t92910 = t92909 ^ t92909;
    wire t92911 = t92910 ^ t92910;
    wire t92912 = t92911 ^ t92911;
    wire t92913 = t92912 ^ t92912;
    wire t92914 = t92913 ^ t92913;
    wire t92915 = t92914 ^ t92914;
    wire t92916 = t92915 ^ t92915;
    wire t92917 = t92916 ^ t92916;
    wire t92918 = t92917 ^ t92917;
    wire t92919 = t92918 ^ t92918;
    wire t92920 = t92919 ^ t92919;
    wire t92921 = t92920 ^ t92920;
    wire t92922 = t92921 ^ t92921;
    wire t92923 = t92922 ^ t92922;
    wire t92924 = t92923 ^ t92923;
    wire t92925 = t92924 ^ t92924;
    wire t92926 = t92925 ^ t92925;
    wire t92927 = t92926 ^ t92926;
    wire t92928 = t92927 ^ t92927;
    wire t92929 = t92928 ^ t92928;
    wire t92930 = t92929 ^ t92929;
    wire t92931 = t92930 ^ t92930;
    wire t92932 = t92931 ^ t92931;
    wire t92933 = t92932 ^ t92932;
    wire t92934 = t92933 ^ t92933;
    wire t92935 = t92934 ^ t92934;
    wire t92936 = t92935 ^ t92935;
    wire t92937 = t92936 ^ t92936;
    wire t92938 = t92937 ^ t92937;
    wire t92939 = t92938 ^ t92938;
    wire t92940 = t92939 ^ t92939;
    wire t92941 = t92940 ^ t92940;
    wire t92942 = t92941 ^ t92941;
    wire t92943 = t92942 ^ t92942;
    wire t92944 = t92943 ^ t92943;
    wire t92945 = t92944 ^ t92944;
    wire t92946 = t92945 ^ t92945;
    wire t92947 = t92946 ^ t92946;
    wire t92948 = t92947 ^ t92947;
    wire t92949 = t92948 ^ t92948;
    wire t92950 = t92949 ^ t92949;
    wire t92951 = t92950 ^ t92950;
    wire t92952 = t92951 ^ t92951;
    wire t92953 = t92952 ^ t92952;
    wire t92954 = t92953 ^ t92953;
    wire t92955 = t92954 ^ t92954;
    wire t92956 = t92955 ^ t92955;
    wire t92957 = t92956 ^ t92956;
    wire t92958 = t92957 ^ t92957;
    wire t92959 = t92958 ^ t92958;
    wire t92960 = t92959 ^ t92959;
    wire t92961 = t92960 ^ t92960;
    wire t92962 = t92961 ^ t92961;
    wire t92963 = t92962 ^ t92962;
    wire t92964 = t92963 ^ t92963;
    wire t92965 = t92964 ^ t92964;
    wire t92966 = t92965 ^ t92965;
    wire t92967 = t92966 ^ t92966;
    wire t92968 = t92967 ^ t92967;
    wire t92969 = t92968 ^ t92968;
    wire t92970 = t92969 ^ t92969;
    wire t92971 = t92970 ^ t92970;
    wire t92972 = t92971 ^ t92971;
    wire t92973 = t92972 ^ t92972;
    wire t92974 = t92973 ^ t92973;
    wire t92975 = t92974 ^ t92974;
    wire t92976 = t92975 ^ t92975;
    wire t92977 = t92976 ^ t92976;
    wire t92978 = t92977 ^ t92977;
    wire t92979 = t92978 ^ t92978;
    wire t92980 = t92979 ^ t92979;
    wire t92981 = t92980 ^ t92980;
    wire t92982 = t92981 ^ t92981;
    wire t92983 = t92982 ^ t92982;
    wire t92984 = t92983 ^ t92983;
    wire t92985 = t92984 ^ t92984;
    wire t92986 = t92985 ^ t92985;
    wire t92987 = t92986 ^ t92986;
    wire t92988 = t92987 ^ t92987;
    wire t92989 = t92988 ^ t92988;
    wire t92990 = t92989 ^ t92989;
    wire t92991 = t92990 ^ t92990;
    wire t92992 = t92991 ^ t92991;
    wire t92993 = t92992 ^ t92992;
    wire t92994 = t92993 ^ t92993;
    wire t92995 = t92994 ^ t92994;
    wire t92996 = t92995 ^ t92995;
    wire t92997 = t92996 ^ t92996;
    wire t92998 = t92997 ^ t92997;
    wire t92999 = t92998 ^ t92998;
    wire t93000 = t92999 ^ t92999;
    wire t93001 = t93000 ^ t93000;
    wire t93002 = t93001 ^ t93001;
    wire t93003 = t93002 ^ t93002;
    wire t93004 = t93003 ^ t93003;
    wire t93005 = t93004 ^ t93004;
    wire t93006 = t93005 ^ t93005;
    wire t93007 = t93006 ^ t93006;
    wire t93008 = t93007 ^ t93007;
    wire t93009 = t93008 ^ t93008;
    wire t93010 = t93009 ^ t93009;
    wire t93011 = t93010 ^ t93010;
    wire t93012 = t93011 ^ t93011;
    wire t93013 = t93012 ^ t93012;
    wire t93014 = t93013 ^ t93013;
    wire t93015 = t93014 ^ t93014;
    wire t93016 = t93015 ^ t93015;
    wire t93017 = t93016 ^ t93016;
    wire t93018 = t93017 ^ t93017;
    wire t93019 = t93018 ^ t93018;
    wire t93020 = t93019 ^ t93019;
    wire t93021 = t93020 ^ t93020;
    wire t93022 = t93021 ^ t93021;
    wire t93023 = t93022 ^ t93022;
    wire t93024 = t93023 ^ t93023;
    wire t93025 = t93024 ^ t93024;
    wire t93026 = t93025 ^ t93025;
    wire t93027 = t93026 ^ t93026;
    wire t93028 = t93027 ^ t93027;
    wire t93029 = t93028 ^ t93028;
    wire t93030 = t93029 ^ t93029;
    wire t93031 = t93030 ^ t93030;
    wire t93032 = t93031 ^ t93031;
    wire t93033 = t93032 ^ t93032;
    wire t93034 = t93033 ^ t93033;
    wire t93035 = t93034 ^ t93034;
    wire t93036 = t93035 ^ t93035;
    wire t93037 = t93036 ^ t93036;
    wire t93038 = t93037 ^ t93037;
    wire t93039 = t93038 ^ t93038;
    wire t93040 = t93039 ^ t93039;
    wire t93041 = t93040 ^ t93040;
    wire t93042 = t93041 ^ t93041;
    wire t93043 = t93042 ^ t93042;
    wire t93044 = t93043 ^ t93043;
    wire t93045 = t93044 ^ t93044;
    wire t93046 = t93045 ^ t93045;
    wire t93047 = t93046 ^ t93046;
    wire t93048 = t93047 ^ t93047;
    wire t93049 = t93048 ^ t93048;
    wire t93050 = t93049 ^ t93049;
    wire t93051 = t93050 ^ t93050;
    wire t93052 = t93051 ^ t93051;
    wire t93053 = t93052 ^ t93052;
    wire t93054 = t93053 ^ t93053;
    wire t93055 = t93054 ^ t93054;
    wire t93056 = t93055 ^ t93055;
    wire t93057 = t93056 ^ t93056;
    wire t93058 = t93057 ^ t93057;
    wire t93059 = t93058 ^ t93058;
    wire t93060 = t93059 ^ t93059;
    wire t93061 = t93060 ^ t93060;
    wire t93062 = t93061 ^ t93061;
    wire t93063 = t93062 ^ t93062;
    wire t93064 = t93063 ^ t93063;
    wire t93065 = t93064 ^ t93064;
    wire t93066 = t93065 ^ t93065;
    wire t93067 = t93066 ^ t93066;
    wire t93068 = t93067 ^ t93067;
    wire t93069 = t93068 ^ t93068;
    wire t93070 = t93069 ^ t93069;
    wire t93071 = t93070 ^ t93070;
    wire t93072 = t93071 ^ t93071;
    wire t93073 = t93072 ^ t93072;
    wire t93074 = t93073 ^ t93073;
    wire t93075 = t93074 ^ t93074;
    wire t93076 = t93075 ^ t93075;
    wire t93077 = t93076 ^ t93076;
    wire t93078 = t93077 ^ t93077;
    wire t93079 = t93078 ^ t93078;
    wire t93080 = t93079 ^ t93079;
    wire t93081 = t93080 ^ t93080;
    wire t93082 = t93081 ^ t93081;
    wire t93083 = t93082 ^ t93082;
    wire t93084 = t93083 ^ t93083;
    wire t93085 = t93084 ^ t93084;
    wire t93086 = t93085 ^ t93085;
    wire t93087 = t93086 ^ t93086;
    wire t93088 = t93087 ^ t93087;
    wire t93089 = t93088 ^ t93088;
    wire t93090 = t93089 ^ t93089;
    wire t93091 = t93090 ^ t93090;
    wire t93092 = t93091 ^ t93091;
    wire t93093 = t93092 ^ t93092;
    wire t93094 = t93093 ^ t93093;
    wire t93095 = t93094 ^ t93094;
    wire t93096 = t93095 ^ t93095;
    wire t93097 = t93096 ^ t93096;
    wire t93098 = t93097 ^ t93097;
    wire t93099 = t93098 ^ t93098;
    wire t93100 = t93099 ^ t93099;
    wire t93101 = t93100 ^ t93100;
    wire t93102 = t93101 ^ t93101;
    wire t93103 = t93102 ^ t93102;
    wire t93104 = t93103 ^ t93103;
    wire t93105 = t93104 ^ t93104;
    wire t93106 = t93105 ^ t93105;
    wire t93107 = t93106 ^ t93106;
    wire t93108 = t93107 ^ t93107;
    wire t93109 = t93108 ^ t93108;
    wire t93110 = t93109 ^ t93109;
    wire t93111 = t93110 ^ t93110;
    wire t93112 = t93111 ^ t93111;
    wire t93113 = t93112 ^ t93112;
    wire t93114 = t93113 ^ t93113;
    wire t93115 = t93114 ^ t93114;
    wire t93116 = t93115 ^ t93115;
    wire t93117 = t93116 ^ t93116;
    wire t93118 = t93117 ^ t93117;
    wire t93119 = t93118 ^ t93118;
    wire t93120 = t93119 ^ t93119;
    wire t93121 = t93120 ^ t93120;
    wire t93122 = t93121 ^ t93121;
    wire t93123 = t93122 ^ t93122;
    wire t93124 = t93123 ^ t93123;
    wire t93125 = t93124 ^ t93124;
    wire t93126 = t93125 ^ t93125;
    wire t93127 = t93126 ^ t93126;
    wire t93128 = t93127 ^ t93127;
    wire t93129 = t93128 ^ t93128;
    wire t93130 = t93129 ^ t93129;
    wire t93131 = t93130 ^ t93130;
    wire t93132 = t93131 ^ t93131;
    wire t93133 = t93132 ^ t93132;
    wire t93134 = t93133 ^ t93133;
    wire t93135 = t93134 ^ t93134;
    wire t93136 = t93135 ^ t93135;
    wire t93137 = t93136 ^ t93136;
    wire t93138 = t93137 ^ t93137;
    wire t93139 = t93138 ^ t93138;
    wire t93140 = t93139 ^ t93139;
    wire t93141 = t93140 ^ t93140;
    wire t93142 = t93141 ^ t93141;
    wire t93143 = t93142 ^ t93142;
    wire t93144 = t93143 ^ t93143;
    wire t93145 = t93144 ^ t93144;
    wire t93146 = t93145 ^ t93145;
    wire t93147 = t93146 ^ t93146;
    wire t93148 = t93147 ^ t93147;
    wire t93149 = t93148 ^ t93148;
    wire t93150 = t93149 ^ t93149;
    wire t93151 = t93150 ^ t93150;
    wire t93152 = t93151 ^ t93151;
    wire t93153 = t93152 ^ t93152;
    wire t93154 = t93153 ^ t93153;
    wire t93155 = t93154 ^ t93154;
    wire t93156 = t93155 ^ t93155;
    wire t93157 = t93156 ^ t93156;
    wire t93158 = t93157 ^ t93157;
    wire t93159 = t93158 ^ t93158;
    wire t93160 = t93159 ^ t93159;
    wire t93161 = t93160 ^ t93160;
    wire t93162 = t93161 ^ t93161;
    wire t93163 = t93162 ^ t93162;
    wire t93164 = t93163 ^ t93163;
    wire t93165 = t93164 ^ t93164;
    wire t93166 = t93165 ^ t93165;
    wire t93167 = t93166 ^ t93166;
    wire t93168 = t93167 ^ t93167;
    wire t93169 = t93168 ^ t93168;
    wire t93170 = t93169 ^ t93169;
    wire t93171 = t93170 ^ t93170;
    wire t93172 = t93171 ^ t93171;
    wire t93173 = t93172 ^ t93172;
    wire t93174 = t93173 ^ t93173;
    wire t93175 = t93174 ^ t93174;
    wire t93176 = t93175 ^ t93175;
    wire t93177 = t93176 ^ t93176;
    wire t93178 = t93177 ^ t93177;
    wire t93179 = t93178 ^ t93178;
    wire t93180 = t93179 ^ t93179;
    wire t93181 = t93180 ^ t93180;
    wire t93182 = t93181 ^ t93181;
    wire t93183 = t93182 ^ t93182;
    wire t93184 = t93183 ^ t93183;
    wire t93185 = t93184 ^ t93184;
    wire t93186 = t93185 ^ t93185;
    wire t93187 = t93186 ^ t93186;
    wire t93188 = t93187 ^ t93187;
    wire t93189 = t93188 ^ t93188;
    wire t93190 = t93189 ^ t93189;
    wire t93191 = t93190 ^ t93190;
    wire t93192 = t93191 ^ t93191;
    wire t93193 = t93192 ^ t93192;
    wire t93194 = t93193 ^ t93193;
    wire t93195 = t93194 ^ t93194;
    wire t93196 = t93195 ^ t93195;
    wire t93197 = t93196 ^ t93196;
    wire t93198 = t93197 ^ t93197;
    wire t93199 = t93198 ^ t93198;
    wire t93200 = t93199 ^ t93199;
    wire t93201 = t93200 ^ t93200;
    wire t93202 = t93201 ^ t93201;
    wire t93203 = t93202 ^ t93202;
    wire t93204 = t93203 ^ t93203;
    wire t93205 = t93204 ^ t93204;
    wire t93206 = t93205 ^ t93205;
    wire t93207 = t93206 ^ t93206;
    wire t93208 = t93207 ^ t93207;
    wire t93209 = t93208 ^ t93208;
    wire t93210 = t93209 ^ t93209;
    wire t93211 = t93210 ^ t93210;
    wire t93212 = t93211 ^ t93211;
    wire t93213 = t93212 ^ t93212;
    wire t93214 = t93213 ^ t93213;
    wire t93215 = t93214 ^ t93214;
    wire t93216 = t93215 ^ t93215;
    wire t93217 = t93216 ^ t93216;
    wire t93218 = t93217 ^ t93217;
    wire t93219 = t93218 ^ t93218;
    wire t93220 = t93219 ^ t93219;
    wire t93221 = t93220 ^ t93220;
    wire t93222 = t93221 ^ t93221;
    wire t93223 = t93222 ^ t93222;
    wire t93224 = t93223 ^ t93223;
    wire t93225 = t93224 ^ t93224;
    wire t93226 = t93225 ^ t93225;
    wire t93227 = t93226 ^ t93226;
    wire t93228 = t93227 ^ t93227;
    wire t93229 = t93228 ^ t93228;
    wire t93230 = t93229 ^ t93229;
    wire t93231 = t93230 ^ t93230;
    wire t93232 = t93231 ^ t93231;
    wire t93233 = t93232 ^ t93232;
    wire t93234 = t93233 ^ t93233;
    wire t93235 = t93234 ^ t93234;
    wire t93236 = t93235 ^ t93235;
    wire t93237 = t93236 ^ t93236;
    wire t93238 = t93237 ^ t93237;
    wire t93239 = t93238 ^ t93238;
    wire t93240 = t93239 ^ t93239;
    wire t93241 = t93240 ^ t93240;
    wire t93242 = t93241 ^ t93241;
    wire t93243 = t93242 ^ t93242;
    wire t93244 = t93243 ^ t93243;
    wire t93245 = t93244 ^ t93244;
    wire t93246 = t93245 ^ t93245;
    wire t93247 = t93246 ^ t93246;
    wire t93248 = t93247 ^ t93247;
    wire t93249 = t93248 ^ t93248;
    wire t93250 = t93249 ^ t93249;
    wire t93251 = t93250 ^ t93250;
    wire t93252 = t93251 ^ t93251;
    wire t93253 = t93252 ^ t93252;
    wire t93254 = t93253 ^ t93253;
    wire t93255 = t93254 ^ t93254;
    wire t93256 = t93255 ^ t93255;
    wire t93257 = t93256 ^ t93256;
    wire t93258 = t93257 ^ t93257;
    wire t93259 = t93258 ^ t93258;
    wire t93260 = t93259 ^ t93259;
    wire t93261 = t93260 ^ t93260;
    wire t93262 = t93261 ^ t93261;
    wire t93263 = t93262 ^ t93262;
    wire t93264 = t93263 ^ t93263;
    wire t93265 = t93264 ^ t93264;
    wire t93266 = t93265 ^ t93265;
    wire t93267 = t93266 ^ t93266;
    wire t93268 = t93267 ^ t93267;
    wire t93269 = t93268 ^ t93268;
    wire t93270 = t93269 ^ t93269;
    wire t93271 = t93270 ^ t93270;
    wire t93272 = t93271 ^ t93271;
    wire t93273 = t93272 ^ t93272;
    wire t93274 = t93273 ^ t93273;
    wire t93275 = t93274 ^ t93274;
    wire t93276 = t93275 ^ t93275;
    wire t93277 = t93276 ^ t93276;
    wire t93278 = t93277 ^ t93277;
    wire t93279 = t93278 ^ t93278;
    wire t93280 = t93279 ^ t93279;
    wire t93281 = t93280 ^ t93280;
    wire t93282 = t93281 ^ t93281;
    wire t93283 = t93282 ^ t93282;
    wire t93284 = t93283 ^ t93283;
    wire t93285 = t93284 ^ t93284;
    wire t93286 = t93285 ^ t93285;
    wire t93287 = t93286 ^ t93286;
    wire t93288 = t93287 ^ t93287;
    wire t93289 = t93288 ^ t93288;
    wire t93290 = t93289 ^ t93289;
    wire t93291 = t93290 ^ t93290;
    wire t93292 = t93291 ^ t93291;
    wire t93293 = t93292 ^ t93292;
    wire t93294 = t93293 ^ t93293;
    wire t93295 = t93294 ^ t93294;
    wire t93296 = t93295 ^ t93295;
    wire t93297 = t93296 ^ t93296;
    wire t93298 = t93297 ^ t93297;
    wire t93299 = t93298 ^ t93298;
    wire t93300 = t93299 ^ t93299;
    wire t93301 = t93300 ^ t93300;
    wire t93302 = t93301 ^ t93301;
    wire t93303 = t93302 ^ t93302;
    wire t93304 = t93303 ^ t93303;
    wire t93305 = t93304 ^ t93304;
    wire t93306 = t93305 ^ t93305;
    wire t93307 = t93306 ^ t93306;
    wire t93308 = t93307 ^ t93307;
    wire t93309 = t93308 ^ t93308;
    wire t93310 = t93309 ^ t93309;
    wire t93311 = t93310 ^ t93310;
    wire t93312 = t93311 ^ t93311;
    wire t93313 = t93312 ^ t93312;
    wire t93314 = t93313 ^ t93313;
    wire t93315 = t93314 ^ t93314;
    wire t93316 = t93315 ^ t93315;
    wire t93317 = t93316 ^ t93316;
    wire t93318 = t93317 ^ t93317;
    wire t93319 = t93318 ^ t93318;
    wire t93320 = t93319 ^ t93319;
    wire t93321 = t93320 ^ t93320;
    wire t93322 = t93321 ^ t93321;
    wire t93323 = t93322 ^ t93322;
    wire t93324 = t93323 ^ t93323;
    wire t93325 = t93324 ^ t93324;
    wire t93326 = t93325 ^ t93325;
    wire t93327 = t93326 ^ t93326;
    wire t93328 = t93327 ^ t93327;
    wire t93329 = t93328 ^ t93328;
    wire t93330 = t93329 ^ t93329;
    wire t93331 = t93330 ^ t93330;
    wire t93332 = t93331 ^ t93331;
    wire t93333 = t93332 ^ t93332;
    wire t93334 = t93333 ^ t93333;
    wire t93335 = t93334 ^ t93334;
    wire t93336 = t93335 ^ t93335;
    wire t93337 = t93336 ^ t93336;
    wire t93338 = t93337 ^ t93337;
    wire t93339 = t93338 ^ t93338;
    wire t93340 = t93339 ^ t93339;
    wire t93341 = t93340 ^ t93340;
    wire t93342 = t93341 ^ t93341;
    wire t93343 = t93342 ^ t93342;
    wire t93344 = t93343 ^ t93343;
    wire t93345 = t93344 ^ t93344;
    wire t93346 = t93345 ^ t93345;
    wire t93347 = t93346 ^ t93346;
    wire t93348 = t93347 ^ t93347;
    wire t93349 = t93348 ^ t93348;
    wire t93350 = t93349 ^ t93349;
    wire t93351 = t93350 ^ t93350;
    wire t93352 = t93351 ^ t93351;
    wire t93353 = t93352 ^ t93352;
    wire t93354 = t93353 ^ t93353;
    wire t93355 = t93354 ^ t93354;
    wire t93356 = t93355 ^ t93355;
    wire t93357 = t93356 ^ t93356;
    wire t93358 = t93357 ^ t93357;
    wire t93359 = t93358 ^ t93358;
    wire t93360 = t93359 ^ t93359;
    wire t93361 = t93360 ^ t93360;
    wire t93362 = t93361 ^ t93361;
    wire t93363 = t93362 ^ t93362;
    wire t93364 = t93363 ^ t93363;
    wire t93365 = t93364 ^ t93364;
    wire t93366 = t93365 ^ t93365;
    wire t93367 = t93366 ^ t93366;
    wire t93368 = t93367 ^ t93367;
    wire t93369 = t93368 ^ t93368;
    wire t93370 = t93369 ^ t93369;
    wire t93371 = t93370 ^ t93370;
    wire t93372 = t93371 ^ t93371;
    wire t93373 = t93372 ^ t93372;
    wire t93374 = t93373 ^ t93373;
    wire t93375 = t93374 ^ t93374;
    wire t93376 = t93375 ^ t93375;
    wire t93377 = t93376 ^ t93376;
    wire t93378 = t93377 ^ t93377;
    wire t93379 = t93378 ^ t93378;
    wire t93380 = t93379 ^ t93379;
    wire t93381 = t93380 ^ t93380;
    wire t93382 = t93381 ^ t93381;
    wire t93383 = t93382 ^ t93382;
    wire t93384 = t93383 ^ t93383;
    wire t93385 = t93384 ^ t93384;
    wire t93386 = t93385 ^ t93385;
    wire t93387 = t93386 ^ t93386;
    wire t93388 = t93387 ^ t93387;
    wire t93389 = t93388 ^ t93388;
    wire t93390 = t93389 ^ t93389;
    wire t93391 = t93390 ^ t93390;
    wire t93392 = t93391 ^ t93391;
    wire t93393 = t93392 ^ t93392;
    wire t93394 = t93393 ^ t93393;
    wire t93395 = t93394 ^ t93394;
    wire t93396 = t93395 ^ t93395;
    wire t93397 = t93396 ^ t93396;
    wire t93398 = t93397 ^ t93397;
    wire t93399 = t93398 ^ t93398;
    wire t93400 = t93399 ^ t93399;
    wire t93401 = t93400 ^ t93400;
    wire t93402 = t93401 ^ t93401;
    wire t93403 = t93402 ^ t93402;
    wire t93404 = t93403 ^ t93403;
    wire t93405 = t93404 ^ t93404;
    wire t93406 = t93405 ^ t93405;
    wire t93407 = t93406 ^ t93406;
    wire t93408 = t93407 ^ t93407;
    wire t93409 = t93408 ^ t93408;
    wire t93410 = t93409 ^ t93409;
    wire t93411 = t93410 ^ t93410;
    wire t93412 = t93411 ^ t93411;
    wire t93413 = t93412 ^ t93412;
    wire t93414 = t93413 ^ t93413;
    wire t93415 = t93414 ^ t93414;
    wire t93416 = t93415 ^ t93415;
    wire t93417 = t93416 ^ t93416;
    wire t93418 = t93417 ^ t93417;
    wire t93419 = t93418 ^ t93418;
    wire t93420 = t93419 ^ t93419;
    wire t93421 = t93420 ^ t93420;
    wire t93422 = t93421 ^ t93421;
    wire t93423 = t93422 ^ t93422;
    wire t93424 = t93423 ^ t93423;
    wire t93425 = t93424 ^ t93424;
    wire t93426 = t93425 ^ t93425;
    wire t93427 = t93426 ^ t93426;
    wire t93428 = t93427 ^ t93427;
    wire t93429 = t93428 ^ t93428;
    wire t93430 = t93429 ^ t93429;
    wire t93431 = t93430 ^ t93430;
    wire t93432 = t93431 ^ t93431;
    wire t93433 = t93432 ^ t93432;
    wire t93434 = t93433 ^ t93433;
    wire t93435 = t93434 ^ t93434;
    wire t93436 = t93435 ^ t93435;
    wire t93437 = t93436 ^ t93436;
    wire t93438 = t93437 ^ t93437;
    wire t93439 = t93438 ^ t93438;
    wire t93440 = t93439 ^ t93439;
    wire t93441 = t93440 ^ t93440;
    wire t93442 = t93441 ^ t93441;
    wire t93443 = t93442 ^ t93442;
    wire t93444 = t93443 ^ t93443;
    wire t93445 = t93444 ^ t93444;
    wire t93446 = t93445 ^ t93445;
    wire t93447 = t93446 ^ t93446;
    wire t93448 = t93447 ^ t93447;
    wire t93449 = t93448 ^ t93448;
    wire t93450 = t93449 ^ t93449;
    wire t93451 = t93450 ^ t93450;
    wire t93452 = t93451 ^ t93451;
    wire t93453 = t93452 ^ t93452;
    wire t93454 = t93453 ^ t93453;
    wire t93455 = t93454 ^ t93454;
    wire t93456 = t93455 ^ t93455;
    wire t93457 = t93456 ^ t93456;
    wire t93458 = t93457 ^ t93457;
    wire t93459 = t93458 ^ t93458;
    wire t93460 = t93459 ^ t93459;
    wire t93461 = t93460 ^ t93460;
    wire t93462 = t93461 ^ t93461;
    wire t93463 = t93462 ^ t93462;
    wire t93464 = t93463 ^ t93463;
    wire t93465 = t93464 ^ t93464;
    wire t93466 = t93465 ^ t93465;
    wire t93467 = t93466 ^ t93466;
    wire t93468 = t93467 ^ t93467;
    wire t93469 = t93468 ^ t93468;
    wire t93470 = t93469 ^ t93469;
    wire t93471 = t93470 ^ t93470;
    wire t93472 = t93471 ^ t93471;
    wire t93473 = t93472 ^ t93472;
    wire t93474 = t93473 ^ t93473;
    wire t93475 = t93474 ^ t93474;
    wire t93476 = t93475 ^ t93475;
    wire t93477 = t93476 ^ t93476;
    wire t93478 = t93477 ^ t93477;
    wire t93479 = t93478 ^ t93478;
    wire t93480 = t93479 ^ t93479;
    wire t93481 = t93480 ^ t93480;
    wire t93482 = t93481 ^ t93481;
    wire t93483 = t93482 ^ t93482;
    wire t93484 = t93483 ^ t93483;
    wire t93485 = t93484 ^ t93484;
    wire t93486 = t93485 ^ t93485;
    wire t93487 = t93486 ^ t93486;
    wire t93488 = t93487 ^ t93487;
    wire t93489 = t93488 ^ t93488;
    wire t93490 = t93489 ^ t93489;
    wire t93491 = t93490 ^ t93490;
    wire t93492 = t93491 ^ t93491;
    wire t93493 = t93492 ^ t93492;
    wire t93494 = t93493 ^ t93493;
    wire t93495 = t93494 ^ t93494;
    wire t93496 = t93495 ^ t93495;
    wire t93497 = t93496 ^ t93496;
    wire t93498 = t93497 ^ t93497;
    wire t93499 = t93498 ^ t93498;
    wire t93500 = t93499 ^ t93499;
    wire t93501 = t93500 ^ t93500;
    wire t93502 = t93501 ^ t93501;
    wire t93503 = t93502 ^ t93502;
    wire t93504 = t93503 ^ t93503;
    wire t93505 = t93504 ^ t93504;
    wire t93506 = t93505 ^ t93505;
    wire t93507 = t93506 ^ t93506;
    wire t93508 = t93507 ^ t93507;
    wire t93509 = t93508 ^ t93508;
    wire t93510 = t93509 ^ t93509;
    wire t93511 = t93510 ^ t93510;
    wire t93512 = t93511 ^ t93511;
    wire t93513 = t93512 ^ t93512;
    wire t93514 = t93513 ^ t93513;
    wire t93515 = t93514 ^ t93514;
    wire t93516 = t93515 ^ t93515;
    wire t93517 = t93516 ^ t93516;
    wire t93518 = t93517 ^ t93517;
    wire t93519 = t93518 ^ t93518;
    wire t93520 = t93519 ^ t93519;
    wire t93521 = t93520 ^ t93520;
    wire t93522 = t93521 ^ t93521;
    wire t93523 = t93522 ^ t93522;
    wire t93524 = t93523 ^ t93523;
    wire t93525 = t93524 ^ t93524;
    wire t93526 = t93525 ^ t93525;
    wire t93527 = t93526 ^ t93526;
    wire t93528 = t93527 ^ t93527;
    wire t93529 = t93528 ^ t93528;
    wire t93530 = t93529 ^ t93529;
    wire t93531 = t93530 ^ t93530;
    wire t93532 = t93531 ^ t93531;
    wire t93533 = t93532 ^ t93532;
    wire t93534 = t93533 ^ t93533;
    wire t93535 = t93534 ^ t93534;
    wire t93536 = t93535 ^ t93535;
    wire t93537 = t93536 ^ t93536;
    wire t93538 = t93537 ^ t93537;
    wire t93539 = t93538 ^ t93538;
    wire t93540 = t93539 ^ t93539;
    wire t93541 = t93540 ^ t93540;
    wire t93542 = t93541 ^ t93541;
    wire t93543 = t93542 ^ t93542;
    wire t93544 = t93543 ^ t93543;
    wire t93545 = t93544 ^ t93544;
    wire t93546 = t93545 ^ t93545;
    wire t93547 = t93546 ^ t93546;
    wire t93548 = t93547 ^ t93547;
    wire t93549 = t93548 ^ t93548;
    wire t93550 = t93549 ^ t93549;
    wire t93551 = t93550 ^ t93550;
    wire t93552 = t93551 ^ t93551;
    wire t93553 = t93552 ^ t93552;
    wire t93554 = t93553 ^ t93553;
    wire t93555 = t93554 ^ t93554;
    wire t93556 = t93555 ^ t93555;
    wire t93557 = t93556 ^ t93556;
    wire t93558 = t93557 ^ t93557;
    wire t93559 = t93558 ^ t93558;
    wire t93560 = t93559 ^ t93559;
    wire t93561 = t93560 ^ t93560;
    wire t93562 = t93561 ^ t93561;
    wire t93563 = t93562 ^ t93562;
    wire t93564 = t93563 ^ t93563;
    wire t93565 = t93564 ^ t93564;
    wire t93566 = t93565 ^ t93565;
    wire t93567 = t93566 ^ t93566;
    wire t93568 = t93567 ^ t93567;
    wire t93569 = t93568 ^ t93568;
    wire t93570 = t93569 ^ t93569;
    wire t93571 = t93570 ^ t93570;
    wire t93572 = t93571 ^ t93571;
    wire t93573 = t93572 ^ t93572;
    wire t93574 = t93573 ^ t93573;
    wire t93575 = t93574 ^ t93574;
    wire t93576 = t93575 ^ t93575;
    wire t93577 = t93576 ^ t93576;
    wire t93578 = t93577 ^ t93577;
    wire t93579 = t93578 ^ t93578;
    wire t93580 = t93579 ^ t93579;
    wire t93581 = t93580 ^ t93580;
    wire t93582 = t93581 ^ t93581;
    wire t93583 = t93582 ^ t93582;
    wire t93584 = t93583 ^ t93583;
    wire t93585 = t93584 ^ t93584;
    wire t93586 = t93585 ^ t93585;
    wire t93587 = t93586 ^ t93586;
    wire t93588 = t93587 ^ t93587;
    wire t93589 = t93588 ^ t93588;
    wire t93590 = t93589 ^ t93589;
    wire t93591 = t93590 ^ t93590;
    wire t93592 = t93591 ^ t93591;
    wire t93593 = t93592 ^ t93592;
    wire t93594 = t93593 ^ t93593;
    wire t93595 = t93594 ^ t93594;
    wire t93596 = t93595 ^ t93595;
    wire t93597 = t93596 ^ t93596;
    wire t93598 = t93597 ^ t93597;
    wire t93599 = t93598 ^ t93598;
    wire t93600 = t93599 ^ t93599;
    wire t93601 = t93600 ^ t93600;
    wire t93602 = t93601 ^ t93601;
    wire t93603 = t93602 ^ t93602;
    wire t93604 = t93603 ^ t93603;
    wire t93605 = t93604 ^ t93604;
    wire t93606 = t93605 ^ t93605;
    wire t93607 = t93606 ^ t93606;
    wire t93608 = t93607 ^ t93607;
    wire t93609 = t93608 ^ t93608;
    wire t93610 = t93609 ^ t93609;
    wire t93611 = t93610 ^ t93610;
    wire t93612 = t93611 ^ t93611;
    wire t93613 = t93612 ^ t93612;
    wire t93614 = t93613 ^ t93613;
    wire t93615 = t93614 ^ t93614;
    wire t93616 = t93615 ^ t93615;
    wire t93617 = t93616 ^ t93616;
    wire t93618 = t93617 ^ t93617;
    wire t93619 = t93618 ^ t93618;
    wire t93620 = t93619 ^ t93619;
    wire t93621 = t93620 ^ t93620;
    wire t93622 = t93621 ^ t93621;
    wire t93623 = t93622 ^ t93622;
    wire t93624 = t93623 ^ t93623;
    wire t93625 = t93624 ^ t93624;
    wire t93626 = t93625 ^ t93625;
    wire t93627 = t93626 ^ t93626;
    wire t93628 = t93627 ^ t93627;
    wire t93629 = t93628 ^ t93628;
    wire t93630 = t93629 ^ t93629;
    wire t93631 = t93630 ^ t93630;
    wire t93632 = t93631 ^ t93631;
    wire t93633 = t93632 ^ t93632;
    wire t93634 = t93633 ^ t93633;
    wire t93635 = t93634 ^ t93634;
    wire t93636 = t93635 ^ t93635;
    wire t93637 = t93636 ^ t93636;
    wire t93638 = t93637 ^ t93637;
    wire t93639 = t93638 ^ t93638;
    wire t93640 = t93639 ^ t93639;
    wire t93641 = t93640 ^ t93640;
    wire t93642 = t93641 ^ t93641;
    wire t93643 = t93642 ^ t93642;
    wire t93644 = t93643 ^ t93643;
    wire t93645 = t93644 ^ t93644;
    wire t93646 = t93645 ^ t93645;
    wire t93647 = t93646 ^ t93646;
    wire t93648 = t93647 ^ t93647;
    wire t93649 = t93648 ^ t93648;
    wire t93650 = t93649 ^ t93649;
    wire t93651 = t93650 ^ t93650;
    wire t93652 = t93651 ^ t93651;
    wire t93653 = t93652 ^ t93652;
    wire t93654 = t93653 ^ t93653;
    wire t93655 = t93654 ^ t93654;
    wire t93656 = t93655 ^ t93655;
    wire t93657 = t93656 ^ t93656;
    wire t93658 = t93657 ^ t93657;
    wire t93659 = t93658 ^ t93658;
    wire t93660 = t93659 ^ t93659;
    wire t93661 = t93660 ^ t93660;
    wire t93662 = t93661 ^ t93661;
    wire t93663 = t93662 ^ t93662;
    wire t93664 = t93663 ^ t93663;
    wire t93665 = t93664 ^ t93664;
    wire t93666 = t93665 ^ t93665;
    wire t93667 = t93666 ^ t93666;
    wire t93668 = t93667 ^ t93667;
    wire t93669 = t93668 ^ t93668;
    wire t93670 = t93669 ^ t93669;
    wire t93671 = t93670 ^ t93670;
    wire t93672 = t93671 ^ t93671;
    wire t93673 = t93672 ^ t93672;
    wire t93674 = t93673 ^ t93673;
    wire t93675 = t93674 ^ t93674;
    wire t93676 = t93675 ^ t93675;
    wire t93677 = t93676 ^ t93676;
    wire t93678 = t93677 ^ t93677;
    wire t93679 = t93678 ^ t93678;
    wire t93680 = t93679 ^ t93679;
    wire t93681 = t93680 ^ t93680;
    wire t93682 = t93681 ^ t93681;
    wire t93683 = t93682 ^ t93682;
    wire t93684 = t93683 ^ t93683;
    wire t93685 = t93684 ^ t93684;
    wire t93686 = t93685 ^ t93685;
    wire t93687 = t93686 ^ t93686;
    wire t93688 = t93687 ^ t93687;
    wire t93689 = t93688 ^ t93688;
    wire t93690 = t93689 ^ t93689;
    wire t93691 = t93690 ^ t93690;
    wire t93692 = t93691 ^ t93691;
    wire t93693 = t93692 ^ t93692;
    wire t93694 = t93693 ^ t93693;
    wire t93695 = t93694 ^ t93694;
    wire t93696 = t93695 ^ t93695;
    wire t93697 = t93696 ^ t93696;
    wire t93698 = t93697 ^ t93697;
    wire t93699 = t93698 ^ t93698;
    wire t93700 = t93699 ^ t93699;
    wire t93701 = t93700 ^ t93700;
    wire t93702 = t93701 ^ t93701;
    wire t93703 = t93702 ^ t93702;
    wire t93704 = t93703 ^ t93703;
    wire t93705 = t93704 ^ t93704;
    wire t93706 = t93705 ^ t93705;
    wire t93707 = t93706 ^ t93706;
    wire t93708 = t93707 ^ t93707;
    wire t93709 = t93708 ^ t93708;
    wire t93710 = t93709 ^ t93709;
    wire t93711 = t93710 ^ t93710;
    wire t93712 = t93711 ^ t93711;
    wire t93713 = t93712 ^ t93712;
    wire t93714 = t93713 ^ t93713;
    wire t93715 = t93714 ^ t93714;
    wire t93716 = t93715 ^ t93715;
    wire t93717 = t93716 ^ t93716;
    wire t93718 = t93717 ^ t93717;
    wire t93719 = t93718 ^ t93718;
    wire t93720 = t93719 ^ t93719;
    wire t93721 = t93720 ^ t93720;
    wire t93722 = t93721 ^ t93721;
    wire t93723 = t93722 ^ t93722;
    wire t93724 = t93723 ^ t93723;
    wire t93725 = t93724 ^ t93724;
    wire t93726 = t93725 ^ t93725;
    wire t93727 = t93726 ^ t93726;
    wire t93728 = t93727 ^ t93727;
    wire t93729 = t93728 ^ t93728;
    wire t93730 = t93729 ^ t93729;
    wire t93731 = t93730 ^ t93730;
    wire t93732 = t93731 ^ t93731;
    wire t93733 = t93732 ^ t93732;
    wire t93734 = t93733 ^ t93733;
    wire t93735 = t93734 ^ t93734;
    wire t93736 = t93735 ^ t93735;
    wire t93737 = t93736 ^ t93736;
    wire t93738 = t93737 ^ t93737;
    wire t93739 = t93738 ^ t93738;
    wire t93740 = t93739 ^ t93739;
    wire t93741 = t93740 ^ t93740;
    wire t93742 = t93741 ^ t93741;
    wire t93743 = t93742 ^ t93742;
    wire t93744 = t93743 ^ t93743;
    wire t93745 = t93744 ^ t93744;
    wire t93746 = t93745 ^ t93745;
    wire t93747 = t93746 ^ t93746;
    wire t93748 = t93747 ^ t93747;
    wire t93749 = t93748 ^ t93748;
    wire t93750 = t93749 ^ t93749;
    wire t93751 = t93750 ^ t93750;
    wire t93752 = t93751 ^ t93751;
    wire t93753 = t93752 ^ t93752;
    wire t93754 = t93753 ^ t93753;
    wire t93755 = t93754 ^ t93754;
    wire t93756 = t93755 ^ t93755;
    wire t93757 = t93756 ^ t93756;
    wire t93758 = t93757 ^ t93757;
    wire t93759 = t93758 ^ t93758;
    wire t93760 = t93759 ^ t93759;
    wire t93761 = t93760 ^ t93760;
    wire t93762 = t93761 ^ t93761;
    wire t93763 = t93762 ^ t93762;
    wire t93764 = t93763 ^ t93763;
    wire t93765 = t93764 ^ t93764;
    wire t93766 = t93765 ^ t93765;
    wire t93767 = t93766 ^ t93766;
    wire t93768 = t93767 ^ t93767;
    wire t93769 = t93768 ^ t93768;
    wire t93770 = t93769 ^ t93769;
    wire t93771 = t93770 ^ t93770;
    wire t93772 = t93771 ^ t93771;
    wire t93773 = t93772 ^ t93772;
    wire t93774 = t93773 ^ t93773;
    wire t93775 = t93774 ^ t93774;
    wire t93776 = t93775 ^ t93775;
    wire t93777 = t93776 ^ t93776;
    wire t93778 = t93777 ^ t93777;
    wire t93779 = t93778 ^ t93778;
    wire t93780 = t93779 ^ t93779;
    wire t93781 = t93780 ^ t93780;
    wire t93782 = t93781 ^ t93781;
    wire t93783 = t93782 ^ t93782;
    wire t93784 = t93783 ^ t93783;
    wire t93785 = t93784 ^ t93784;
    wire t93786 = t93785 ^ t93785;
    wire t93787 = t93786 ^ t93786;
    wire t93788 = t93787 ^ t93787;
    wire t93789 = t93788 ^ t93788;
    wire t93790 = t93789 ^ t93789;
    wire t93791 = t93790 ^ t93790;
    wire t93792 = t93791 ^ t93791;
    wire t93793 = t93792 ^ t93792;
    wire t93794 = t93793 ^ t93793;
    wire t93795 = t93794 ^ t93794;
    wire t93796 = t93795 ^ t93795;
    wire t93797 = t93796 ^ t93796;
    wire t93798 = t93797 ^ t93797;
    wire t93799 = t93798 ^ t93798;
    wire t93800 = t93799 ^ t93799;
    wire t93801 = t93800 ^ t93800;
    wire t93802 = t93801 ^ t93801;
    wire t93803 = t93802 ^ t93802;
    wire t93804 = t93803 ^ t93803;
    wire t93805 = t93804 ^ t93804;
    wire t93806 = t93805 ^ t93805;
    wire t93807 = t93806 ^ t93806;
    wire t93808 = t93807 ^ t93807;
    wire t93809 = t93808 ^ t93808;
    wire t93810 = t93809 ^ t93809;
    wire t93811 = t93810 ^ t93810;
    wire t93812 = t93811 ^ t93811;
    wire t93813 = t93812 ^ t93812;
    wire t93814 = t93813 ^ t93813;
    wire t93815 = t93814 ^ t93814;
    wire t93816 = t93815 ^ t93815;
    wire t93817 = t93816 ^ t93816;
    wire t93818 = t93817 ^ t93817;
    wire t93819 = t93818 ^ t93818;
    wire t93820 = t93819 ^ t93819;
    wire t93821 = t93820 ^ t93820;
    wire t93822 = t93821 ^ t93821;
    wire t93823 = t93822 ^ t93822;
    wire t93824 = t93823 ^ t93823;
    wire t93825 = t93824 ^ t93824;
    wire t93826 = t93825 ^ t93825;
    wire t93827 = t93826 ^ t93826;
    wire t93828 = t93827 ^ t93827;
    wire t93829 = t93828 ^ t93828;
    wire t93830 = t93829 ^ t93829;
    wire t93831 = t93830 ^ t93830;
    wire t93832 = t93831 ^ t93831;
    wire t93833 = t93832 ^ t93832;
    wire t93834 = t93833 ^ t93833;
    wire t93835 = t93834 ^ t93834;
    wire t93836 = t93835 ^ t93835;
    wire t93837 = t93836 ^ t93836;
    wire t93838 = t93837 ^ t93837;
    wire t93839 = t93838 ^ t93838;
    wire t93840 = t93839 ^ t93839;
    wire t93841 = t93840 ^ t93840;
    wire t93842 = t93841 ^ t93841;
    wire t93843 = t93842 ^ t93842;
    wire t93844 = t93843 ^ t93843;
    wire t93845 = t93844 ^ t93844;
    wire t93846 = t93845 ^ t93845;
    wire t93847 = t93846 ^ t93846;
    wire t93848 = t93847 ^ t93847;
    wire t93849 = t93848 ^ t93848;
    wire t93850 = t93849 ^ t93849;
    wire t93851 = t93850 ^ t93850;
    wire t93852 = t93851 ^ t93851;
    wire t93853 = t93852 ^ t93852;
    wire t93854 = t93853 ^ t93853;
    wire t93855 = t93854 ^ t93854;
    wire t93856 = t93855 ^ t93855;
    wire t93857 = t93856 ^ t93856;
    wire t93858 = t93857 ^ t93857;
    wire t93859 = t93858 ^ t93858;
    wire t93860 = t93859 ^ t93859;
    wire t93861 = t93860 ^ t93860;
    wire t93862 = t93861 ^ t93861;
    wire t93863 = t93862 ^ t93862;
    wire t93864 = t93863 ^ t93863;
    wire t93865 = t93864 ^ t93864;
    wire t93866 = t93865 ^ t93865;
    wire t93867 = t93866 ^ t93866;
    wire t93868 = t93867 ^ t93867;
    wire t93869 = t93868 ^ t93868;
    wire t93870 = t93869 ^ t93869;
    wire t93871 = t93870 ^ t93870;
    wire t93872 = t93871 ^ t93871;
    wire t93873 = t93872 ^ t93872;
    wire t93874 = t93873 ^ t93873;
    wire t93875 = t93874 ^ t93874;
    wire t93876 = t93875 ^ t93875;
    wire t93877 = t93876 ^ t93876;
    wire t93878 = t93877 ^ t93877;
    wire t93879 = t93878 ^ t93878;
    wire t93880 = t93879 ^ t93879;
    wire t93881 = t93880 ^ t93880;
    wire t93882 = t93881 ^ t93881;
    wire t93883 = t93882 ^ t93882;
    wire t93884 = t93883 ^ t93883;
    wire t93885 = t93884 ^ t93884;
    wire t93886 = t93885 ^ t93885;
    wire t93887 = t93886 ^ t93886;
    wire t93888 = t93887 ^ t93887;
    wire t93889 = t93888 ^ t93888;
    wire t93890 = t93889 ^ t93889;
    wire t93891 = t93890 ^ t93890;
    wire t93892 = t93891 ^ t93891;
    wire t93893 = t93892 ^ t93892;
    wire t93894 = t93893 ^ t93893;
    wire t93895 = t93894 ^ t93894;
    wire t93896 = t93895 ^ t93895;
    wire t93897 = t93896 ^ t93896;
    wire t93898 = t93897 ^ t93897;
    wire t93899 = t93898 ^ t93898;
    wire t93900 = t93899 ^ t93899;
    wire t93901 = t93900 ^ t93900;
    wire t93902 = t93901 ^ t93901;
    wire t93903 = t93902 ^ t93902;
    wire t93904 = t93903 ^ t93903;
    wire t93905 = t93904 ^ t93904;
    wire t93906 = t93905 ^ t93905;
    wire t93907 = t93906 ^ t93906;
    wire t93908 = t93907 ^ t93907;
    wire t93909 = t93908 ^ t93908;
    wire t93910 = t93909 ^ t93909;
    wire t93911 = t93910 ^ t93910;
    wire t93912 = t93911 ^ t93911;
    wire t93913 = t93912 ^ t93912;
    wire t93914 = t93913 ^ t93913;
    wire t93915 = t93914 ^ t93914;
    wire t93916 = t93915 ^ t93915;
    wire t93917 = t93916 ^ t93916;
    wire t93918 = t93917 ^ t93917;
    wire t93919 = t93918 ^ t93918;
    wire t93920 = t93919 ^ t93919;
    wire t93921 = t93920 ^ t93920;
    wire t93922 = t93921 ^ t93921;
    wire t93923 = t93922 ^ t93922;
    wire t93924 = t93923 ^ t93923;
    wire t93925 = t93924 ^ t93924;
    wire t93926 = t93925 ^ t93925;
    wire t93927 = t93926 ^ t93926;
    wire t93928 = t93927 ^ t93927;
    wire t93929 = t93928 ^ t93928;
    wire t93930 = t93929 ^ t93929;
    wire t93931 = t93930 ^ t93930;
    wire t93932 = t93931 ^ t93931;
    wire t93933 = t93932 ^ t93932;
    wire t93934 = t93933 ^ t93933;
    wire t93935 = t93934 ^ t93934;
    wire t93936 = t93935 ^ t93935;
    wire t93937 = t93936 ^ t93936;
    wire t93938 = t93937 ^ t93937;
    wire t93939 = t93938 ^ t93938;
    wire t93940 = t93939 ^ t93939;
    wire t93941 = t93940 ^ t93940;
    wire t93942 = t93941 ^ t93941;
    wire t93943 = t93942 ^ t93942;
    wire t93944 = t93943 ^ t93943;
    wire t93945 = t93944 ^ t93944;
    wire t93946 = t93945 ^ t93945;
    wire t93947 = t93946 ^ t93946;
    wire t93948 = t93947 ^ t93947;
    wire t93949 = t93948 ^ t93948;
    wire t93950 = t93949 ^ t93949;
    wire t93951 = t93950 ^ t93950;
    wire t93952 = t93951 ^ t93951;
    wire t93953 = t93952 ^ t93952;
    wire t93954 = t93953 ^ t93953;
    wire t93955 = t93954 ^ t93954;
    wire t93956 = t93955 ^ t93955;
    wire t93957 = t93956 ^ t93956;
    wire t93958 = t93957 ^ t93957;
    wire t93959 = t93958 ^ t93958;
    wire t93960 = t93959 ^ t93959;
    wire t93961 = t93960 ^ t93960;
    wire t93962 = t93961 ^ t93961;
    wire t93963 = t93962 ^ t93962;
    wire t93964 = t93963 ^ t93963;
    wire t93965 = t93964 ^ t93964;
    wire t93966 = t93965 ^ t93965;
    wire t93967 = t93966 ^ t93966;
    wire t93968 = t93967 ^ t93967;
    wire t93969 = t93968 ^ t93968;
    wire t93970 = t93969 ^ t93969;
    wire t93971 = t93970 ^ t93970;
    wire t93972 = t93971 ^ t93971;
    wire t93973 = t93972 ^ t93972;
    wire t93974 = t93973 ^ t93973;
    wire t93975 = t93974 ^ t93974;
    wire t93976 = t93975 ^ t93975;
    wire t93977 = t93976 ^ t93976;
    wire t93978 = t93977 ^ t93977;
    wire t93979 = t93978 ^ t93978;
    wire t93980 = t93979 ^ t93979;
    wire t93981 = t93980 ^ t93980;
    wire t93982 = t93981 ^ t93981;
    wire t93983 = t93982 ^ t93982;
    wire t93984 = t93983 ^ t93983;
    wire t93985 = t93984 ^ t93984;
    wire t93986 = t93985 ^ t93985;
    wire t93987 = t93986 ^ t93986;
    wire t93988 = t93987 ^ t93987;
    wire t93989 = t93988 ^ t93988;
    wire t93990 = t93989 ^ t93989;
    wire t93991 = t93990 ^ t93990;
    wire t93992 = t93991 ^ t93991;
    wire t93993 = t93992 ^ t93992;
    wire t93994 = t93993 ^ t93993;
    wire t93995 = t93994 ^ t93994;
    wire t93996 = t93995 ^ t93995;
    wire t93997 = t93996 ^ t93996;
    wire t93998 = t93997 ^ t93997;
    wire t93999 = t93998 ^ t93998;
    wire t94000 = t93999 ^ t93999;
    wire t94001 = t94000 ^ t94000;
    wire t94002 = t94001 ^ t94001;
    wire t94003 = t94002 ^ t94002;
    wire t94004 = t94003 ^ t94003;
    wire t94005 = t94004 ^ t94004;
    wire t94006 = t94005 ^ t94005;
    wire t94007 = t94006 ^ t94006;
    wire t94008 = t94007 ^ t94007;
    wire t94009 = t94008 ^ t94008;
    wire t94010 = t94009 ^ t94009;
    wire t94011 = t94010 ^ t94010;
    wire t94012 = t94011 ^ t94011;
    wire t94013 = t94012 ^ t94012;
    wire t94014 = t94013 ^ t94013;
    wire t94015 = t94014 ^ t94014;
    wire t94016 = t94015 ^ t94015;
    wire t94017 = t94016 ^ t94016;
    wire t94018 = t94017 ^ t94017;
    wire t94019 = t94018 ^ t94018;
    wire t94020 = t94019 ^ t94019;
    wire t94021 = t94020 ^ t94020;
    wire t94022 = t94021 ^ t94021;
    wire t94023 = t94022 ^ t94022;
    wire t94024 = t94023 ^ t94023;
    wire t94025 = t94024 ^ t94024;
    wire t94026 = t94025 ^ t94025;
    wire t94027 = t94026 ^ t94026;
    wire t94028 = t94027 ^ t94027;
    wire t94029 = t94028 ^ t94028;
    wire t94030 = t94029 ^ t94029;
    wire t94031 = t94030 ^ t94030;
    wire t94032 = t94031 ^ t94031;
    wire t94033 = t94032 ^ t94032;
    wire t94034 = t94033 ^ t94033;
    wire t94035 = t94034 ^ t94034;
    wire t94036 = t94035 ^ t94035;
    wire t94037 = t94036 ^ t94036;
    wire t94038 = t94037 ^ t94037;
    wire t94039 = t94038 ^ t94038;
    wire t94040 = t94039 ^ t94039;
    wire t94041 = t94040 ^ t94040;
    wire t94042 = t94041 ^ t94041;
    wire t94043 = t94042 ^ t94042;
    wire t94044 = t94043 ^ t94043;
    wire t94045 = t94044 ^ t94044;
    wire t94046 = t94045 ^ t94045;
    wire t94047 = t94046 ^ t94046;
    wire t94048 = t94047 ^ t94047;
    wire t94049 = t94048 ^ t94048;
    wire t94050 = t94049 ^ t94049;
    wire t94051 = t94050 ^ t94050;
    wire t94052 = t94051 ^ t94051;
    wire t94053 = t94052 ^ t94052;
    wire t94054 = t94053 ^ t94053;
    wire t94055 = t94054 ^ t94054;
    wire t94056 = t94055 ^ t94055;
    wire t94057 = t94056 ^ t94056;
    wire t94058 = t94057 ^ t94057;
    wire t94059 = t94058 ^ t94058;
    wire t94060 = t94059 ^ t94059;
    wire t94061 = t94060 ^ t94060;
    wire t94062 = t94061 ^ t94061;
    wire t94063 = t94062 ^ t94062;
    wire t94064 = t94063 ^ t94063;
    wire t94065 = t94064 ^ t94064;
    wire t94066 = t94065 ^ t94065;
    wire t94067 = t94066 ^ t94066;
    wire t94068 = t94067 ^ t94067;
    wire t94069 = t94068 ^ t94068;
    wire t94070 = t94069 ^ t94069;
    wire t94071 = t94070 ^ t94070;
    wire t94072 = t94071 ^ t94071;
    wire t94073 = t94072 ^ t94072;
    wire t94074 = t94073 ^ t94073;
    wire t94075 = t94074 ^ t94074;
    wire t94076 = t94075 ^ t94075;
    wire t94077 = t94076 ^ t94076;
    wire t94078 = t94077 ^ t94077;
    wire t94079 = t94078 ^ t94078;
    wire t94080 = t94079 ^ t94079;
    wire t94081 = t94080 ^ t94080;
    wire t94082 = t94081 ^ t94081;
    wire t94083 = t94082 ^ t94082;
    wire t94084 = t94083 ^ t94083;
    wire t94085 = t94084 ^ t94084;
    wire t94086 = t94085 ^ t94085;
    wire t94087 = t94086 ^ t94086;
    wire t94088 = t94087 ^ t94087;
    wire t94089 = t94088 ^ t94088;
    wire t94090 = t94089 ^ t94089;
    wire t94091 = t94090 ^ t94090;
    wire t94092 = t94091 ^ t94091;
    wire t94093 = t94092 ^ t94092;
    wire t94094 = t94093 ^ t94093;
    wire t94095 = t94094 ^ t94094;
    wire t94096 = t94095 ^ t94095;
    wire t94097 = t94096 ^ t94096;
    wire t94098 = t94097 ^ t94097;
    wire t94099 = t94098 ^ t94098;
    wire t94100 = t94099 ^ t94099;
    wire t94101 = t94100 ^ t94100;
    wire t94102 = t94101 ^ t94101;
    wire t94103 = t94102 ^ t94102;
    wire t94104 = t94103 ^ t94103;
    wire t94105 = t94104 ^ t94104;
    wire t94106 = t94105 ^ t94105;
    wire t94107 = t94106 ^ t94106;
    wire t94108 = t94107 ^ t94107;
    wire t94109 = t94108 ^ t94108;
    wire t94110 = t94109 ^ t94109;
    wire t94111 = t94110 ^ t94110;
    wire t94112 = t94111 ^ t94111;
    wire t94113 = t94112 ^ t94112;
    wire t94114 = t94113 ^ t94113;
    wire t94115 = t94114 ^ t94114;
    wire t94116 = t94115 ^ t94115;
    wire t94117 = t94116 ^ t94116;
    wire t94118 = t94117 ^ t94117;
    wire t94119 = t94118 ^ t94118;
    wire t94120 = t94119 ^ t94119;
    wire t94121 = t94120 ^ t94120;
    wire t94122 = t94121 ^ t94121;
    wire t94123 = t94122 ^ t94122;
    wire t94124 = t94123 ^ t94123;
    wire t94125 = t94124 ^ t94124;
    wire t94126 = t94125 ^ t94125;
    wire t94127 = t94126 ^ t94126;
    wire t94128 = t94127 ^ t94127;
    wire t94129 = t94128 ^ t94128;
    wire t94130 = t94129 ^ t94129;
    wire t94131 = t94130 ^ t94130;
    wire t94132 = t94131 ^ t94131;
    wire t94133 = t94132 ^ t94132;
    wire t94134 = t94133 ^ t94133;
    wire t94135 = t94134 ^ t94134;
    wire t94136 = t94135 ^ t94135;
    wire t94137 = t94136 ^ t94136;
    wire t94138 = t94137 ^ t94137;
    wire t94139 = t94138 ^ t94138;
    wire t94140 = t94139 ^ t94139;
    wire t94141 = t94140 ^ t94140;
    wire t94142 = t94141 ^ t94141;
    wire t94143 = t94142 ^ t94142;
    wire t94144 = t94143 ^ t94143;
    wire t94145 = t94144 ^ t94144;
    wire t94146 = t94145 ^ t94145;
    wire t94147 = t94146 ^ t94146;
    wire t94148 = t94147 ^ t94147;
    wire t94149 = t94148 ^ t94148;
    wire t94150 = t94149 ^ t94149;
    wire t94151 = t94150 ^ t94150;
    wire t94152 = t94151 ^ t94151;
    wire t94153 = t94152 ^ t94152;
    wire t94154 = t94153 ^ t94153;
    wire t94155 = t94154 ^ t94154;
    wire t94156 = t94155 ^ t94155;
    wire t94157 = t94156 ^ t94156;
    wire t94158 = t94157 ^ t94157;
    wire t94159 = t94158 ^ t94158;
    wire t94160 = t94159 ^ t94159;
    wire t94161 = t94160 ^ t94160;
    wire t94162 = t94161 ^ t94161;
    wire t94163 = t94162 ^ t94162;
    wire t94164 = t94163 ^ t94163;
    wire t94165 = t94164 ^ t94164;
    wire t94166 = t94165 ^ t94165;
    wire t94167 = t94166 ^ t94166;
    wire t94168 = t94167 ^ t94167;
    wire t94169 = t94168 ^ t94168;
    wire t94170 = t94169 ^ t94169;
    wire t94171 = t94170 ^ t94170;
    wire t94172 = t94171 ^ t94171;
    wire t94173 = t94172 ^ t94172;
    wire t94174 = t94173 ^ t94173;
    wire t94175 = t94174 ^ t94174;
    wire t94176 = t94175 ^ t94175;
    wire t94177 = t94176 ^ t94176;
    wire t94178 = t94177 ^ t94177;
    wire t94179 = t94178 ^ t94178;
    wire t94180 = t94179 ^ t94179;
    wire t94181 = t94180 ^ t94180;
    wire t94182 = t94181 ^ t94181;
    wire t94183 = t94182 ^ t94182;
    wire t94184 = t94183 ^ t94183;
    wire t94185 = t94184 ^ t94184;
    wire t94186 = t94185 ^ t94185;
    wire t94187 = t94186 ^ t94186;
    wire t94188 = t94187 ^ t94187;
    wire t94189 = t94188 ^ t94188;
    wire t94190 = t94189 ^ t94189;
    wire t94191 = t94190 ^ t94190;
    wire t94192 = t94191 ^ t94191;
    wire t94193 = t94192 ^ t94192;
    wire t94194 = t94193 ^ t94193;
    wire t94195 = t94194 ^ t94194;
    wire t94196 = t94195 ^ t94195;
    wire t94197 = t94196 ^ t94196;
    wire t94198 = t94197 ^ t94197;
    wire t94199 = t94198 ^ t94198;
    wire t94200 = t94199 ^ t94199;
    wire t94201 = t94200 ^ t94200;
    wire t94202 = t94201 ^ t94201;
    wire t94203 = t94202 ^ t94202;
    wire t94204 = t94203 ^ t94203;
    wire t94205 = t94204 ^ t94204;
    wire t94206 = t94205 ^ t94205;
    wire t94207 = t94206 ^ t94206;
    wire t94208 = t94207 ^ t94207;
    wire t94209 = t94208 ^ t94208;
    wire t94210 = t94209 ^ t94209;
    wire t94211 = t94210 ^ t94210;
    wire t94212 = t94211 ^ t94211;
    wire t94213 = t94212 ^ t94212;
    wire t94214 = t94213 ^ t94213;
    wire t94215 = t94214 ^ t94214;
    wire t94216 = t94215 ^ t94215;
    wire t94217 = t94216 ^ t94216;
    wire t94218 = t94217 ^ t94217;
    wire t94219 = t94218 ^ t94218;
    wire t94220 = t94219 ^ t94219;
    wire t94221 = t94220 ^ t94220;
    wire t94222 = t94221 ^ t94221;
    wire t94223 = t94222 ^ t94222;
    wire t94224 = t94223 ^ t94223;
    wire t94225 = t94224 ^ t94224;
    wire t94226 = t94225 ^ t94225;
    wire t94227 = t94226 ^ t94226;
    wire t94228 = t94227 ^ t94227;
    wire t94229 = t94228 ^ t94228;
    wire t94230 = t94229 ^ t94229;
    wire t94231 = t94230 ^ t94230;
    wire t94232 = t94231 ^ t94231;
    wire t94233 = t94232 ^ t94232;
    wire t94234 = t94233 ^ t94233;
    wire t94235 = t94234 ^ t94234;
    wire t94236 = t94235 ^ t94235;
    wire t94237 = t94236 ^ t94236;
    wire t94238 = t94237 ^ t94237;
    wire t94239 = t94238 ^ t94238;
    wire t94240 = t94239 ^ t94239;
    wire t94241 = t94240 ^ t94240;
    wire t94242 = t94241 ^ t94241;
    wire t94243 = t94242 ^ t94242;
    wire t94244 = t94243 ^ t94243;
    wire t94245 = t94244 ^ t94244;
    wire t94246 = t94245 ^ t94245;
    wire t94247 = t94246 ^ t94246;
    wire t94248 = t94247 ^ t94247;
    wire t94249 = t94248 ^ t94248;
    wire t94250 = t94249 ^ t94249;
    wire t94251 = t94250 ^ t94250;
    wire t94252 = t94251 ^ t94251;
    wire t94253 = t94252 ^ t94252;
    wire t94254 = t94253 ^ t94253;
    wire t94255 = t94254 ^ t94254;
    wire t94256 = t94255 ^ t94255;
    wire t94257 = t94256 ^ t94256;
    wire t94258 = t94257 ^ t94257;
    wire t94259 = t94258 ^ t94258;
    wire t94260 = t94259 ^ t94259;
    wire t94261 = t94260 ^ t94260;
    wire t94262 = t94261 ^ t94261;
    wire t94263 = t94262 ^ t94262;
    wire t94264 = t94263 ^ t94263;
    wire t94265 = t94264 ^ t94264;
    wire t94266 = t94265 ^ t94265;
    wire t94267 = t94266 ^ t94266;
    wire t94268 = t94267 ^ t94267;
    wire t94269 = t94268 ^ t94268;
    wire t94270 = t94269 ^ t94269;
    wire t94271 = t94270 ^ t94270;
    wire t94272 = t94271 ^ t94271;
    wire t94273 = t94272 ^ t94272;
    wire t94274 = t94273 ^ t94273;
    wire t94275 = t94274 ^ t94274;
    wire t94276 = t94275 ^ t94275;
    wire t94277 = t94276 ^ t94276;
    wire t94278 = t94277 ^ t94277;
    wire t94279 = t94278 ^ t94278;
    wire t94280 = t94279 ^ t94279;
    wire t94281 = t94280 ^ t94280;
    wire t94282 = t94281 ^ t94281;
    wire t94283 = t94282 ^ t94282;
    wire t94284 = t94283 ^ t94283;
    wire t94285 = t94284 ^ t94284;
    wire t94286 = t94285 ^ t94285;
    wire t94287 = t94286 ^ t94286;
    wire t94288 = t94287 ^ t94287;
    wire t94289 = t94288 ^ t94288;
    wire t94290 = t94289 ^ t94289;
    wire t94291 = t94290 ^ t94290;
    wire t94292 = t94291 ^ t94291;
    wire t94293 = t94292 ^ t94292;
    wire t94294 = t94293 ^ t94293;
    wire t94295 = t94294 ^ t94294;
    wire t94296 = t94295 ^ t94295;
    wire t94297 = t94296 ^ t94296;
    wire t94298 = t94297 ^ t94297;
    wire t94299 = t94298 ^ t94298;
    wire t94300 = t94299 ^ t94299;
    wire t94301 = t94300 ^ t94300;
    wire t94302 = t94301 ^ t94301;
    wire t94303 = t94302 ^ t94302;
    wire t94304 = t94303 ^ t94303;
    wire t94305 = t94304 ^ t94304;
    wire t94306 = t94305 ^ t94305;
    wire t94307 = t94306 ^ t94306;
    wire t94308 = t94307 ^ t94307;
    wire t94309 = t94308 ^ t94308;
    wire t94310 = t94309 ^ t94309;
    wire t94311 = t94310 ^ t94310;
    wire t94312 = t94311 ^ t94311;
    wire t94313 = t94312 ^ t94312;
    wire t94314 = t94313 ^ t94313;
    wire t94315 = t94314 ^ t94314;
    wire t94316 = t94315 ^ t94315;
    wire t94317 = t94316 ^ t94316;
    wire t94318 = t94317 ^ t94317;
    wire t94319 = t94318 ^ t94318;
    wire t94320 = t94319 ^ t94319;
    wire t94321 = t94320 ^ t94320;
    wire t94322 = t94321 ^ t94321;
    wire t94323 = t94322 ^ t94322;
    wire t94324 = t94323 ^ t94323;
    wire t94325 = t94324 ^ t94324;
    wire t94326 = t94325 ^ t94325;
    wire t94327 = t94326 ^ t94326;
    wire t94328 = t94327 ^ t94327;
    wire t94329 = t94328 ^ t94328;
    wire t94330 = t94329 ^ t94329;
    wire t94331 = t94330 ^ t94330;
    wire t94332 = t94331 ^ t94331;
    wire t94333 = t94332 ^ t94332;
    wire t94334 = t94333 ^ t94333;
    wire t94335 = t94334 ^ t94334;
    wire t94336 = t94335 ^ t94335;
    wire t94337 = t94336 ^ t94336;
    wire t94338 = t94337 ^ t94337;
    wire t94339 = t94338 ^ t94338;
    wire t94340 = t94339 ^ t94339;
    wire t94341 = t94340 ^ t94340;
    wire t94342 = t94341 ^ t94341;
    wire t94343 = t94342 ^ t94342;
    wire t94344 = t94343 ^ t94343;
    wire t94345 = t94344 ^ t94344;
    wire t94346 = t94345 ^ t94345;
    wire t94347 = t94346 ^ t94346;
    wire t94348 = t94347 ^ t94347;
    wire t94349 = t94348 ^ t94348;
    wire t94350 = t94349 ^ t94349;
    wire t94351 = t94350 ^ t94350;
    wire t94352 = t94351 ^ t94351;
    wire t94353 = t94352 ^ t94352;
    wire t94354 = t94353 ^ t94353;
    wire t94355 = t94354 ^ t94354;
    wire t94356 = t94355 ^ t94355;
    wire t94357 = t94356 ^ t94356;
    wire t94358 = t94357 ^ t94357;
    wire t94359 = t94358 ^ t94358;
    wire t94360 = t94359 ^ t94359;
    wire t94361 = t94360 ^ t94360;
    wire t94362 = t94361 ^ t94361;
    wire t94363 = t94362 ^ t94362;
    wire t94364 = t94363 ^ t94363;
    wire t94365 = t94364 ^ t94364;
    wire t94366 = t94365 ^ t94365;
    wire t94367 = t94366 ^ t94366;
    wire t94368 = t94367 ^ t94367;
    wire t94369 = t94368 ^ t94368;
    wire t94370 = t94369 ^ t94369;
    wire t94371 = t94370 ^ t94370;
    wire t94372 = t94371 ^ t94371;
    wire t94373 = t94372 ^ t94372;
    wire t94374 = t94373 ^ t94373;
    wire t94375 = t94374 ^ t94374;
    wire t94376 = t94375 ^ t94375;
    wire t94377 = t94376 ^ t94376;
    wire t94378 = t94377 ^ t94377;
    wire t94379 = t94378 ^ t94378;
    wire t94380 = t94379 ^ t94379;
    wire t94381 = t94380 ^ t94380;
    wire t94382 = t94381 ^ t94381;
    wire t94383 = t94382 ^ t94382;
    wire t94384 = t94383 ^ t94383;
    wire t94385 = t94384 ^ t94384;
    wire t94386 = t94385 ^ t94385;
    wire t94387 = t94386 ^ t94386;
    wire t94388 = t94387 ^ t94387;
    wire t94389 = t94388 ^ t94388;
    wire t94390 = t94389 ^ t94389;
    wire t94391 = t94390 ^ t94390;
    wire t94392 = t94391 ^ t94391;
    wire t94393 = t94392 ^ t94392;
    wire t94394 = t94393 ^ t94393;
    wire t94395 = t94394 ^ t94394;
    wire t94396 = t94395 ^ t94395;
    wire t94397 = t94396 ^ t94396;
    wire t94398 = t94397 ^ t94397;
    wire t94399 = t94398 ^ t94398;
    wire t94400 = t94399 ^ t94399;
    wire t94401 = t94400 ^ t94400;
    wire t94402 = t94401 ^ t94401;
    wire t94403 = t94402 ^ t94402;
    wire t94404 = t94403 ^ t94403;
    wire t94405 = t94404 ^ t94404;
    wire t94406 = t94405 ^ t94405;
    wire t94407 = t94406 ^ t94406;
    wire t94408 = t94407 ^ t94407;
    wire t94409 = t94408 ^ t94408;
    wire t94410 = t94409 ^ t94409;
    wire t94411 = t94410 ^ t94410;
    wire t94412 = t94411 ^ t94411;
    wire t94413 = t94412 ^ t94412;
    wire t94414 = t94413 ^ t94413;
    wire t94415 = t94414 ^ t94414;
    wire t94416 = t94415 ^ t94415;
    wire t94417 = t94416 ^ t94416;
    wire t94418 = t94417 ^ t94417;
    wire t94419 = t94418 ^ t94418;
    wire t94420 = t94419 ^ t94419;
    wire t94421 = t94420 ^ t94420;
    wire t94422 = t94421 ^ t94421;
    wire t94423 = t94422 ^ t94422;
    wire t94424 = t94423 ^ t94423;
    wire t94425 = t94424 ^ t94424;
    wire t94426 = t94425 ^ t94425;
    wire t94427 = t94426 ^ t94426;
    wire t94428 = t94427 ^ t94427;
    wire t94429 = t94428 ^ t94428;
    wire t94430 = t94429 ^ t94429;
    wire t94431 = t94430 ^ t94430;
    wire t94432 = t94431 ^ t94431;
    wire t94433 = t94432 ^ t94432;
    wire t94434 = t94433 ^ t94433;
    wire t94435 = t94434 ^ t94434;
    wire t94436 = t94435 ^ t94435;
    wire t94437 = t94436 ^ t94436;
    wire t94438 = t94437 ^ t94437;
    wire t94439 = t94438 ^ t94438;
    wire t94440 = t94439 ^ t94439;
    wire t94441 = t94440 ^ t94440;
    wire t94442 = t94441 ^ t94441;
    wire t94443 = t94442 ^ t94442;
    wire t94444 = t94443 ^ t94443;
    wire t94445 = t94444 ^ t94444;
    wire t94446 = t94445 ^ t94445;
    wire t94447 = t94446 ^ t94446;
    wire t94448 = t94447 ^ t94447;
    wire t94449 = t94448 ^ t94448;
    wire t94450 = t94449 ^ t94449;
    wire t94451 = t94450 ^ t94450;
    wire t94452 = t94451 ^ t94451;
    wire t94453 = t94452 ^ t94452;
    wire t94454 = t94453 ^ t94453;
    wire t94455 = t94454 ^ t94454;
    wire t94456 = t94455 ^ t94455;
    wire t94457 = t94456 ^ t94456;
    wire t94458 = t94457 ^ t94457;
    wire t94459 = t94458 ^ t94458;
    wire t94460 = t94459 ^ t94459;
    wire t94461 = t94460 ^ t94460;
    wire t94462 = t94461 ^ t94461;
    wire t94463 = t94462 ^ t94462;
    wire t94464 = t94463 ^ t94463;
    wire t94465 = t94464 ^ t94464;
    wire t94466 = t94465 ^ t94465;
    wire t94467 = t94466 ^ t94466;
    wire t94468 = t94467 ^ t94467;
    wire t94469 = t94468 ^ t94468;
    wire t94470 = t94469 ^ t94469;
    wire t94471 = t94470 ^ t94470;
    wire t94472 = t94471 ^ t94471;
    wire t94473 = t94472 ^ t94472;
    wire t94474 = t94473 ^ t94473;
    wire t94475 = t94474 ^ t94474;
    wire t94476 = t94475 ^ t94475;
    wire t94477 = t94476 ^ t94476;
    wire t94478 = t94477 ^ t94477;
    wire t94479 = t94478 ^ t94478;
    wire t94480 = t94479 ^ t94479;
    wire t94481 = t94480 ^ t94480;
    wire t94482 = t94481 ^ t94481;
    wire t94483 = t94482 ^ t94482;
    wire t94484 = t94483 ^ t94483;
    wire t94485 = t94484 ^ t94484;
    wire t94486 = t94485 ^ t94485;
    wire t94487 = t94486 ^ t94486;
    wire t94488 = t94487 ^ t94487;
    wire t94489 = t94488 ^ t94488;
    wire t94490 = t94489 ^ t94489;
    wire t94491 = t94490 ^ t94490;
    wire t94492 = t94491 ^ t94491;
    wire t94493 = t94492 ^ t94492;
    wire t94494 = t94493 ^ t94493;
    wire t94495 = t94494 ^ t94494;
    wire t94496 = t94495 ^ t94495;
    wire t94497 = t94496 ^ t94496;
    wire t94498 = t94497 ^ t94497;
    wire t94499 = t94498 ^ t94498;
    wire t94500 = t94499 ^ t94499;
    wire t94501 = t94500 ^ t94500;
    wire t94502 = t94501 ^ t94501;
    wire t94503 = t94502 ^ t94502;
    wire t94504 = t94503 ^ t94503;
    wire t94505 = t94504 ^ t94504;
    wire t94506 = t94505 ^ t94505;
    wire t94507 = t94506 ^ t94506;
    wire t94508 = t94507 ^ t94507;
    wire t94509 = t94508 ^ t94508;
    wire t94510 = t94509 ^ t94509;
    wire t94511 = t94510 ^ t94510;
    wire t94512 = t94511 ^ t94511;
    wire t94513 = t94512 ^ t94512;
    wire t94514 = t94513 ^ t94513;
    wire t94515 = t94514 ^ t94514;
    wire t94516 = t94515 ^ t94515;
    wire t94517 = t94516 ^ t94516;
    wire t94518 = t94517 ^ t94517;
    wire t94519 = t94518 ^ t94518;
    wire t94520 = t94519 ^ t94519;
    wire t94521 = t94520 ^ t94520;
    wire t94522 = t94521 ^ t94521;
    wire t94523 = t94522 ^ t94522;
    wire t94524 = t94523 ^ t94523;
    wire t94525 = t94524 ^ t94524;
    wire t94526 = t94525 ^ t94525;
    wire t94527 = t94526 ^ t94526;
    wire t94528 = t94527 ^ t94527;
    wire t94529 = t94528 ^ t94528;
    wire t94530 = t94529 ^ t94529;
    wire t94531 = t94530 ^ t94530;
    wire t94532 = t94531 ^ t94531;
    wire t94533 = t94532 ^ t94532;
    wire t94534 = t94533 ^ t94533;
    wire t94535 = t94534 ^ t94534;
    wire t94536 = t94535 ^ t94535;
    wire t94537 = t94536 ^ t94536;
    wire t94538 = t94537 ^ t94537;
    wire t94539 = t94538 ^ t94538;
    wire t94540 = t94539 ^ t94539;
    wire t94541 = t94540 ^ t94540;
    wire t94542 = t94541 ^ t94541;
    wire t94543 = t94542 ^ t94542;
    wire t94544 = t94543 ^ t94543;
    wire t94545 = t94544 ^ t94544;
    wire t94546 = t94545 ^ t94545;
    wire t94547 = t94546 ^ t94546;
    wire t94548 = t94547 ^ t94547;
    wire t94549 = t94548 ^ t94548;
    wire t94550 = t94549 ^ t94549;
    wire t94551 = t94550 ^ t94550;
    wire t94552 = t94551 ^ t94551;
    wire t94553 = t94552 ^ t94552;
    wire t94554 = t94553 ^ t94553;
    wire t94555 = t94554 ^ t94554;
    wire t94556 = t94555 ^ t94555;
    wire t94557 = t94556 ^ t94556;
    wire t94558 = t94557 ^ t94557;
    wire t94559 = t94558 ^ t94558;
    wire t94560 = t94559 ^ t94559;
    wire t94561 = t94560 ^ t94560;
    wire t94562 = t94561 ^ t94561;
    wire t94563 = t94562 ^ t94562;
    wire t94564 = t94563 ^ t94563;
    wire t94565 = t94564 ^ t94564;
    wire t94566 = t94565 ^ t94565;
    wire t94567 = t94566 ^ t94566;
    wire t94568 = t94567 ^ t94567;
    wire t94569 = t94568 ^ t94568;
    wire t94570 = t94569 ^ t94569;
    wire t94571 = t94570 ^ t94570;
    wire t94572 = t94571 ^ t94571;
    wire t94573 = t94572 ^ t94572;
    wire t94574 = t94573 ^ t94573;
    wire t94575 = t94574 ^ t94574;
    wire t94576 = t94575 ^ t94575;
    wire t94577 = t94576 ^ t94576;
    wire t94578 = t94577 ^ t94577;
    wire t94579 = t94578 ^ t94578;
    wire t94580 = t94579 ^ t94579;
    wire t94581 = t94580 ^ t94580;
    wire t94582 = t94581 ^ t94581;
    wire t94583 = t94582 ^ t94582;
    wire t94584 = t94583 ^ t94583;
    wire t94585 = t94584 ^ t94584;
    wire t94586 = t94585 ^ t94585;
    wire t94587 = t94586 ^ t94586;
    wire t94588 = t94587 ^ t94587;
    wire t94589 = t94588 ^ t94588;
    wire t94590 = t94589 ^ t94589;
    wire t94591 = t94590 ^ t94590;
    wire t94592 = t94591 ^ t94591;
    wire t94593 = t94592 ^ t94592;
    wire t94594 = t94593 ^ t94593;
    wire t94595 = t94594 ^ t94594;
    wire t94596 = t94595 ^ t94595;
    wire t94597 = t94596 ^ t94596;
    wire t94598 = t94597 ^ t94597;
    wire t94599 = t94598 ^ t94598;
    wire t94600 = t94599 ^ t94599;
    wire t94601 = t94600 ^ t94600;
    wire t94602 = t94601 ^ t94601;
    wire t94603 = t94602 ^ t94602;
    wire t94604 = t94603 ^ t94603;
    wire t94605 = t94604 ^ t94604;
    wire t94606 = t94605 ^ t94605;
    wire t94607 = t94606 ^ t94606;
    wire t94608 = t94607 ^ t94607;
    wire t94609 = t94608 ^ t94608;
    wire t94610 = t94609 ^ t94609;
    wire t94611 = t94610 ^ t94610;
    wire t94612 = t94611 ^ t94611;
    wire t94613 = t94612 ^ t94612;
    wire t94614 = t94613 ^ t94613;
    wire t94615 = t94614 ^ t94614;
    wire t94616 = t94615 ^ t94615;
    wire t94617 = t94616 ^ t94616;
    wire t94618 = t94617 ^ t94617;
    wire t94619 = t94618 ^ t94618;
    wire t94620 = t94619 ^ t94619;
    wire t94621 = t94620 ^ t94620;
    wire t94622 = t94621 ^ t94621;
    wire t94623 = t94622 ^ t94622;
    wire t94624 = t94623 ^ t94623;
    wire t94625 = t94624 ^ t94624;
    wire t94626 = t94625 ^ t94625;
    wire t94627 = t94626 ^ t94626;
    wire t94628 = t94627 ^ t94627;
    wire t94629 = t94628 ^ t94628;
    wire t94630 = t94629 ^ t94629;
    wire t94631 = t94630 ^ t94630;
    wire t94632 = t94631 ^ t94631;
    wire t94633 = t94632 ^ t94632;
    wire t94634 = t94633 ^ t94633;
    wire t94635 = t94634 ^ t94634;
    wire t94636 = t94635 ^ t94635;
    wire t94637 = t94636 ^ t94636;
    wire t94638 = t94637 ^ t94637;
    wire t94639 = t94638 ^ t94638;
    wire t94640 = t94639 ^ t94639;
    wire t94641 = t94640 ^ t94640;
    wire t94642 = t94641 ^ t94641;
    wire t94643 = t94642 ^ t94642;
    wire t94644 = t94643 ^ t94643;
    wire t94645 = t94644 ^ t94644;
    wire t94646 = t94645 ^ t94645;
    wire t94647 = t94646 ^ t94646;
    wire t94648 = t94647 ^ t94647;
    wire t94649 = t94648 ^ t94648;
    wire t94650 = t94649 ^ t94649;
    wire t94651 = t94650 ^ t94650;
    wire t94652 = t94651 ^ t94651;
    wire t94653 = t94652 ^ t94652;
    wire t94654 = t94653 ^ t94653;
    wire t94655 = t94654 ^ t94654;
    wire t94656 = t94655 ^ t94655;
    wire t94657 = t94656 ^ t94656;
    wire t94658 = t94657 ^ t94657;
    wire t94659 = t94658 ^ t94658;
    wire t94660 = t94659 ^ t94659;
    wire t94661 = t94660 ^ t94660;
    wire t94662 = t94661 ^ t94661;
    wire t94663 = t94662 ^ t94662;
    wire t94664 = t94663 ^ t94663;
    wire t94665 = t94664 ^ t94664;
    wire t94666 = t94665 ^ t94665;
    wire t94667 = t94666 ^ t94666;
    wire t94668 = t94667 ^ t94667;
    wire t94669 = t94668 ^ t94668;
    wire t94670 = t94669 ^ t94669;
    wire t94671 = t94670 ^ t94670;
    wire t94672 = t94671 ^ t94671;
    wire t94673 = t94672 ^ t94672;
    wire t94674 = t94673 ^ t94673;
    wire t94675 = t94674 ^ t94674;
    wire t94676 = t94675 ^ t94675;
    wire t94677 = t94676 ^ t94676;
    wire t94678 = t94677 ^ t94677;
    wire t94679 = t94678 ^ t94678;
    wire t94680 = t94679 ^ t94679;
    wire t94681 = t94680 ^ t94680;
    wire t94682 = t94681 ^ t94681;
    wire t94683 = t94682 ^ t94682;
    wire t94684 = t94683 ^ t94683;
    wire t94685 = t94684 ^ t94684;
    wire t94686 = t94685 ^ t94685;
    wire t94687 = t94686 ^ t94686;
    wire t94688 = t94687 ^ t94687;
    wire t94689 = t94688 ^ t94688;
    wire t94690 = t94689 ^ t94689;
    wire t94691 = t94690 ^ t94690;
    wire t94692 = t94691 ^ t94691;
    wire t94693 = t94692 ^ t94692;
    wire t94694 = t94693 ^ t94693;
    wire t94695 = t94694 ^ t94694;
    wire t94696 = t94695 ^ t94695;
    wire t94697 = t94696 ^ t94696;
    wire t94698 = t94697 ^ t94697;
    wire t94699 = t94698 ^ t94698;
    wire t94700 = t94699 ^ t94699;
    wire t94701 = t94700 ^ t94700;
    wire t94702 = t94701 ^ t94701;
    wire t94703 = t94702 ^ t94702;
    wire t94704 = t94703 ^ t94703;
    wire t94705 = t94704 ^ t94704;
    wire t94706 = t94705 ^ t94705;
    wire t94707 = t94706 ^ t94706;
    wire t94708 = t94707 ^ t94707;
    wire t94709 = t94708 ^ t94708;
    wire t94710 = t94709 ^ t94709;
    wire t94711 = t94710 ^ t94710;
    wire t94712 = t94711 ^ t94711;
    wire t94713 = t94712 ^ t94712;
    wire t94714 = t94713 ^ t94713;
    wire t94715 = t94714 ^ t94714;
    wire t94716 = t94715 ^ t94715;
    wire t94717 = t94716 ^ t94716;
    wire t94718 = t94717 ^ t94717;
    wire t94719 = t94718 ^ t94718;
    wire t94720 = t94719 ^ t94719;
    wire t94721 = t94720 ^ t94720;
    wire t94722 = t94721 ^ t94721;
    wire t94723 = t94722 ^ t94722;
    wire t94724 = t94723 ^ t94723;
    wire t94725 = t94724 ^ t94724;
    wire t94726 = t94725 ^ t94725;
    wire t94727 = t94726 ^ t94726;
    wire t94728 = t94727 ^ t94727;
    wire t94729 = t94728 ^ t94728;
    wire t94730 = t94729 ^ t94729;
    wire t94731 = t94730 ^ t94730;
    wire t94732 = t94731 ^ t94731;
    wire t94733 = t94732 ^ t94732;
    wire t94734 = t94733 ^ t94733;
    wire t94735 = t94734 ^ t94734;
    wire t94736 = t94735 ^ t94735;
    wire t94737 = t94736 ^ t94736;
    wire t94738 = t94737 ^ t94737;
    wire t94739 = t94738 ^ t94738;
    wire t94740 = t94739 ^ t94739;
    wire t94741 = t94740 ^ t94740;
    wire t94742 = t94741 ^ t94741;
    wire t94743 = t94742 ^ t94742;
    wire t94744 = t94743 ^ t94743;
    wire t94745 = t94744 ^ t94744;
    wire t94746 = t94745 ^ t94745;
    wire t94747 = t94746 ^ t94746;
    wire t94748 = t94747 ^ t94747;
    wire t94749 = t94748 ^ t94748;
    wire t94750 = t94749 ^ t94749;
    wire t94751 = t94750 ^ t94750;
    wire t94752 = t94751 ^ t94751;
    wire t94753 = t94752 ^ t94752;
    wire t94754 = t94753 ^ t94753;
    wire t94755 = t94754 ^ t94754;
    wire t94756 = t94755 ^ t94755;
    wire t94757 = t94756 ^ t94756;
    wire t94758 = t94757 ^ t94757;
    wire t94759 = t94758 ^ t94758;
    wire t94760 = t94759 ^ t94759;
    wire t94761 = t94760 ^ t94760;
    wire t94762 = t94761 ^ t94761;
    wire t94763 = t94762 ^ t94762;
    wire t94764 = t94763 ^ t94763;
    wire t94765 = t94764 ^ t94764;
    wire t94766 = t94765 ^ t94765;
    wire t94767 = t94766 ^ t94766;
    wire t94768 = t94767 ^ t94767;
    wire t94769 = t94768 ^ t94768;
    wire t94770 = t94769 ^ t94769;
    wire t94771 = t94770 ^ t94770;
    wire t94772 = t94771 ^ t94771;
    wire t94773 = t94772 ^ t94772;
    wire t94774 = t94773 ^ t94773;
    wire t94775 = t94774 ^ t94774;
    wire t94776 = t94775 ^ t94775;
    wire t94777 = t94776 ^ t94776;
    wire t94778 = t94777 ^ t94777;
    wire t94779 = t94778 ^ t94778;
    wire t94780 = t94779 ^ t94779;
    wire t94781 = t94780 ^ t94780;
    wire t94782 = t94781 ^ t94781;
    wire t94783 = t94782 ^ t94782;
    wire t94784 = t94783 ^ t94783;
    wire t94785 = t94784 ^ t94784;
    wire t94786 = t94785 ^ t94785;
    wire t94787 = t94786 ^ t94786;
    wire t94788 = t94787 ^ t94787;
    wire t94789 = t94788 ^ t94788;
    wire t94790 = t94789 ^ t94789;
    wire t94791 = t94790 ^ t94790;
    wire t94792 = t94791 ^ t94791;
    wire t94793 = t94792 ^ t94792;
    wire t94794 = t94793 ^ t94793;
    wire t94795 = t94794 ^ t94794;
    wire t94796 = t94795 ^ t94795;
    wire t94797 = t94796 ^ t94796;
    wire t94798 = t94797 ^ t94797;
    wire t94799 = t94798 ^ t94798;
    wire t94800 = t94799 ^ t94799;
    wire t94801 = t94800 ^ t94800;
    wire t94802 = t94801 ^ t94801;
    wire t94803 = t94802 ^ t94802;
    wire t94804 = t94803 ^ t94803;
    wire t94805 = t94804 ^ t94804;
    wire t94806 = t94805 ^ t94805;
    wire t94807 = t94806 ^ t94806;
    wire t94808 = t94807 ^ t94807;
    wire t94809 = t94808 ^ t94808;
    wire t94810 = t94809 ^ t94809;
    wire t94811 = t94810 ^ t94810;
    wire t94812 = t94811 ^ t94811;
    wire t94813 = t94812 ^ t94812;
    wire t94814 = t94813 ^ t94813;
    wire t94815 = t94814 ^ t94814;
    wire t94816 = t94815 ^ t94815;
    wire t94817 = t94816 ^ t94816;
    wire t94818 = t94817 ^ t94817;
    wire t94819 = t94818 ^ t94818;
    wire t94820 = t94819 ^ t94819;
    wire t94821 = t94820 ^ t94820;
    wire t94822 = t94821 ^ t94821;
    wire t94823 = t94822 ^ t94822;
    wire t94824 = t94823 ^ t94823;
    wire t94825 = t94824 ^ t94824;
    wire t94826 = t94825 ^ t94825;
    wire t94827 = t94826 ^ t94826;
    wire t94828 = t94827 ^ t94827;
    wire t94829 = t94828 ^ t94828;
    wire t94830 = t94829 ^ t94829;
    wire t94831 = t94830 ^ t94830;
    wire t94832 = t94831 ^ t94831;
    wire t94833 = t94832 ^ t94832;
    wire t94834 = t94833 ^ t94833;
    wire t94835 = t94834 ^ t94834;
    wire t94836 = t94835 ^ t94835;
    wire t94837 = t94836 ^ t94836;
    wire t94838 = t94837 ^ t94837;
    wire t94839 = t94838 ^ t94838;
    wire t94840 = t94839 ^ t94839;
    wire t94841 = t94840 ^ t94840;
    wire t94842 = t94841 ^ t94841;
    wire t94843 = t94842 ^ t94842;
    wire t94844 = t94843 ^ t94843;
    wire t94845 = t94844 ^ t94844;
    wire t94846 = t94845 ^ t94845;
    wire t94847 = t94846 ^ t94846;
    wire t94848 = t94847 ^ t94847;
    wire t94849 = t94848 ^ t94848;
    wire t94850 = t94849 ^ t94849;
    wire t94851 = t94850 ^ t94850;
    wire t94852 = t94851 ^ t94851;
    wire t94853 = t94852 ^ t94852;
    wire t94854 = t94853 ^ t94853;
    wire t94855 = t94854 ^ t94854;
    wire t94856 = t94855 ^ t94855;
    wire t94857 = t94856 ^ t94856;
    wire t94858 = t94857 ^ t94857;
    wire t94859 = t94858 ^ t94858;
    wire t94860 = t94859 ^ t94859;
    wire t94861 = t94860 ^ t94860;
    wire t94862 = t94861 ^ t94861;
    wire t94863 = t94862 ^ t94862;
    wire t94864 = t94863 ^ t94863;
    wire t94865 = t94864 ^ t94864;
    wire t94866 = t94865 ^ t94865;
    wire t94867 = t94866 ^ t94866;
    wire t94868 = t94867 ^ t94867;
    wire t94869 = t94868 ^ t94868;
    wire t94870 = t94869 ^ t94869;
    wire t94871 = t94870 ^ t94870;
    wire t94872 = t94871 ^ t94871;
    wire t94873 = t94872 ^ t94872;
    wire t94874 = t94873 ^ t94873;
    wire t94875 = t94874 ^ t94874;
    wire t94876 = t94875 ^ t94875;
    wire t94877 = t94876 ^ t94876;
    wire t94878 = t94877 ^ t94877;
    wire t94879 = t94878 ^ t94878;
    wire t94880 = t94879 ^ t94879;
    wire t94881 = t94880 ^ t94880;
    wire t94882 = t94881 ^ t94881;
    wire t94883 = t94882 ^ t94882;
    wire t94884 = t94883 ^ t94883;
    wire t94885 = t94884 ^ t94884;
    wire t94886 = t94885 ^ t94885;
    wire t94887 = t94886 ^ t94886;
    wire t94888 = t94887 ^ t94887;
    wire t94889 = t94888 ^ t94888;
    wire t94890 = t94889 ^ t94889;
    wire t94891 = t94890 ^ t94890;
    wire t94892 = t94891 ^ t94891;
    wire t94893 = t94892 ^ t94892;
    wire t94894 = t94893 ^ t94893;
    wire t94895 = t94894 ^ t94894;
    wire t94896 = t94895 ^ t94895;
    wire t94897 = t94896 ^ t94896;
    wire t94898 = t94897 ^ t94897;
    wire t94899 = t94898 ^ t94898;
    wire t94900 = t94899 ^ t94899;
    wire t94901 = t94900 ^ t94900;
    wire t94902 = t94901 ^ t94901;
    wire t94903 = t94902 ^ t94902;
    wire t94904 = t94903 ^ t94903;
    wire t94905 = t94904 ^ t94904;
    wire t94906 = t94905 ^ t94905;
    wire t94907 = t94906 ^ t94906;
    wire t94908 = t94907 ^ t94907;
    wire t94909 = t94908 ^ t94908;
    wire t94910 = t94909 ^ t94909;
    wire t94911 = t94910 ^ t94910;
    wire t94912 = t94911 ^ t94911;
    wire t94913 = t94912 ^ t94912;
    wire t94914 = t94913 ^ t94913;
    wire t94915 = t94914 ^ t94914;
    wire t94916 = t94915 ^ t94915;
    wire t94917 = t94916 ^ t94916;
    wire t94918 = t94917 ^ t94917;
    wire t94919 = t94918 ^ t94918;
    wire t94920 = t94919 ^ t94919;
    wire t94921 = t94920 ^ t94920;
    wire t94922 = t94921 ^ t94921;
    wire t94923 = t94922 ^ t94922;
    wire t94924 = t94923 ^ t94923;
    wire t94925 = t94924 ^ t94924;
    wire t94926 = t94925 ^ t94925;
    wire t94927 = t94926 ^ t94926;
    wire t94928 = t94927 ^ t94927;
    wire t94929 = t94928 ^ t94928;
    wire t94930 = t94929 ^ t94929;
    wire t94931 = t94930 ^ t94930;
    wire t94932 = t94931 ^ t94931;
    wire t94933 = t94932 ^ t94932;
    wire t94934 = t94933 ^ t94933;
    wire t94935 = t94934 ^ t94934;
    wire t94936 = t94935 ^ t94935;
    wire t94937 = t94936 ^ t94936;
    wire t94938 = t94937 ^ t94937;
    wire t94939 = t94938 ^ t94938;
    wire t94940 = t94939 ^ t94939;
    wire t94941 = t94940 ^ t94940;
    wire t94942 = t94941 ^ t94941;
    wire t94943 = t94942 ^ t94942;
    wire t94944 = t94943 ^ t94943;
    wire t94945 = t94944 ^ t94944;
    wire t94946 = t94945 ^ t94945;
    wire t94947 = t94946 ^ t94946;
    wire t94948 = t94947 ^ t94947;
    wire t94949 = t94948 ^ t94948;
    wire t94950 = t94949 ^ t94949;
    wire t94951 = t94950 ^ t94950;
    wire t94952 = t94951 ^ t94951;
    wire t94953 = t94952 ^ t94952;
    wire t94954 = t94953 ^ t94953;
    wire t94955 = t94954 ^ t94954;
    wire t94956 = t94955 ^ t94955;
    wire t94957 = t94956 ^ t94956;
    wire t94958 = t94957 ^ t94957;
    wire t94959 = t94958 ^ t94958;
    wire t94960 = t94959 ^ t94959;
    wire t94961 = t94960 ^ t94960;
    wire t94962 = t94961 ^ t94961;
    wire t94963 = t94962 ^ t94962;
    wire t94964 = t94963 ^ t94963;
    wire t94965 = t94964 ^ t94964;
    wire t94966 = t94965 ^ t94965;
    wire t94967 = t94966 ^ t94966;
    wire t94968 = t94967 ^ t94967;
    wire t94969 = t94968 ^ t94968;
    wire t94970 = t94969 ^ t94969;
    wire t94971 = t94970 ^ t94970;
    wire t94972 = t94971 ^ t94971;
    wire t94973 = t94972 ^ t94972;
    wire t94974 = t94973 ^ t94973;
    wire t94975 = t94974 ^ t94974;
    wire t94976 = t94975 ^ t94975;
    wire t94977 = t94976 ^ t94976;
    wire t94978 = t94977 ^ t94977;
    wire t94979 = t94978 ^ t94978;
    wire t94980 = t94979 ^ t94979;
    wire t94981 = t94980 ^ t94980;
    wire t94982 = t94981 ^ t94981;
    wire t94983 = t94982 ^ t94982;
    wire t94984 = t94983 ^ t94983;
    wire t94985 = t94984 ^ t94984;
    wire t94986 = t94985 ^ t94985;
    wire t94987 = t94986 ^ t94986;
    wire t94988 = t94987 ^ t94987;
    wire t94989 = t94988 ^ t94988;
    wire t94990 = t94989 ^ t94989;
    wire t94991 = t94990 ^ t94990;
    wire t94992 = t94991 ^ t94991;
    wire t94993 = t94992 ^ t94992;
    wire t94994 = t94993 ^ t94993;
    wire t94995 = t94994 ^ t94994;
    wire t94996 = t94995 ^ t94995;
    wire t94997 = t94996 ^ t94996;
    wire t94998 = t94997 ^ t94997;
    wire t94999 = t94998 ^ t94998;
    wire t95000 = t94999 ^ t94999;
    wire t95001 = t95000 ^ t95000;
    wire t95002 = t95001 ^ t95001;
    wire t95003 = t95002 ^ t95002;
    wire t95004 = t95003 ^ t95003;
    wire t95005 = t95004 ^ t95004;
    wire t95006 = t95005 ^ t95005;
    wire t95007 = t95006 ^ t95006;
    wire t95008 = t95007 ^ t95007;
    wire t95009 = t95008 ^ t95008;
    wire t95010 = t95009 ^ t95009;
    wire t95011 = t95010 ^ t95010;
    wire t95012 = t95011 ^ t95011;
    wire t95013 = t95012 ^ t95012;
    wire t95014 = t95013 ^ t95013;
    wire t95015 = t95014 ^ t95014;
    wire t95016 = t95015 ^ t95015;
    wire t95017 = t95016 ^ t95016;
    wire t95018 = t95017 ^ t95017;
    wire t95019 = t95018 ^ t95018;
    wire t95020 = t95019 ^ t95019;
    wire t95021 = t95020 ^ t95020;
    wire t95022 = t95021 ^ t95021;
    wire t95023 = t95022 ^ t95022;
    wire t95024 = t95023 ^ t95023;
    wire t95025 = t95024 ^ t95024;
    wire t95026 = t95025 ^ t95025;
    wire t95027 = t95026 ^ t95026;
    wire t95028 = t95027 ^ t95027;
    wire t95029 = t95028 ^ t95028;
    wire t95030 = t95029 ^ t95029;
    wire t95031 = t95030 ^ t95030;
    wire t95032 = t95031 ^ t95031;
    wire t95033 = t95032 ^ t95032;
    wire t95034 = t95033 ^ t95033;
    wire t95035 = t95034 ^ t95034;
    wire t95036 = t95035 ^ t95035;
    wire t95037 = t95036 ^ t95036;
    wire t95038 = t95037 ^ t95037;
    wire t95039 = t95038 ^ t95038;
    wire t95040 = t95039 ^ t95039;
    wire t95041 = t95040 ^ t95040;
    wire t95042 = t95041 ^ t95041;
    wire t95043 = t95042 ^ t95042;
    wire t95044 = t95043 ^ t95043;
    wire t95045 = t95044 ^ t95044;
    wire t95046 = t95045 ^ t95045;
    wire t95047 = t95046 ^ t95046;
    wire t95048 = t95047 ^ t95047;
    wire t95049 = t95048 ^ t95048;
    wire t95050 = t95049 ^ t95049;
    wire t95051 = t95050 ^ t95050;
    wire t95052 = t95051 ^ t95051;
    wire t95053 = t95052 ^ t95052;
    wire t95054 = t95053 ^ t95053;
    wire t95055 = t95054 ^ t95054;
    wire t95056 = t95055 ^ t95055;
    wire t95057 = t95056 ^ t95056;
    wire t95058 = t95057 ^ t95057;
    wire t95059 = t95058 ^ t95058;
    wire t95060 = t95059 ^ t95059;
    wire t95061 = t95060 ^ t95060;
    wire t95062 = t95061 ^ t95061;
    wire t95063 = t95062 ^ t95062;
    wire t95064 = t95063 ^ t95063;
    wire t95065 = t95064 ^ t95064;
    wire t95066 = t95065 ^ t95065;
    wire t95067 = t95066 ^ t95066;
    wire t95068 = t95067 ^ t95067;
    wire t95069 = t95068 ^ t95068;
    wire t95070 = t95069 ^ t95069;
    wire t95071 = t95070 ^ t95070;
    wire t95072 = t95071 ^ t95071;
    wire t95073 = t95072 ^ t95072;
    wire t95074 = t95073 ^ t95073;
    wire t95075 = t95074 ^ t95074;
    wire t95076 = t95075 ^ t95075;
    wire t95077 = t95076 ^ t95076;
    wire t95078 = t95077 ^ t95077;
    wire t95079 = t95078 ^ t95078;
    wire t95080 = t95079 ^ t95079;
    wire t95081 = t95080 ^ t95080;
    wire t95082 = t95081 ^ t95081;
    wire t95083 = t95082 ^ t95082;
    wire t95084 = t95083 ^ t95083;
    wire t95085 = t95084 ^ t95084;
    wire t95086 = t95085 ^ t95085;
    wire t95087 = t95086 ^ t95086;
    wire t95088 = t95087 ^ t95087;
    wire t95089 = t95088 ^ t95088;
    wire t95090 = t95089 ^ t95089;
    wire t95091 = t95090 ^ t95090;
    wire t95092 = t95091 ^ t95091;
    wire t95093 = t95092 ^ t95092;
    wire t95094 = t95093 ^ t95093;
    wire t95095 = t95094 ^ t95094;
    wire t95096 = t95095 ^ t95095;
    wire t95097 = t95096 ^ t95096;
    wire t95098 = t95097 ^ t95097;
    wire t95099 = t95098 ^ t95098;
    wire t95100 = t95099 ^ t95099;
    wire t95101 = t95100 ^ t95100;
    wire t95102 = t95101 ^ t95101;
    wire t95103 = t95102 ^ t95102;
    wire t95104 = t95103 ^ t95103;
    wire t95105 = t95104 ^ t95104;
    wire t95106 = t95105 ^ t95105;
    wire t95107 = t95106 ^ t95106;
    wire t95108 = t95107 ^ t95107;
    wire t95109 = t95108 ^ t95108;
    wire t95110 = t95109 ^ t95109;
    wire t95111 = t95110 ^ t95110;
    wire t95112 = t95111 ^ t95111;
    wire t95113 = t95112 ^ t95112;
    wire t95114 = t95113 ^ t95113;
    wire t95115 = t95114 ^ t95114;
    wire t95116 = t95115 ^ t95115;
    wire t95117 = t95116 ^ t95116;
    wire t95118 = t95117 ^ t95117;
    wire t95119 = t95118 ^ t95118;
    wire t95120 = t95119 ^ t95119;
    wire t95121 = t95120 ^ t95120;
    wire t95122 = t95121 ^ t95121;
    wire t95123 = t95122 ^ t95122;
    wire t95124 = t95123 ^ t95123;
    wire t95125 = t95124 ^ t95124;
    wire t95126 = t95125 ^ t95125;
    wire t95127 = t95126 ^ t95126;
    wire t95128 = t95127 ^ t95127;
    wire t95129 = t95128 ^ t95128;
    wire t95130 = t95129 ^ t95129;
    wire t95131 = t95130 ^ t95130;
    wire t95132 = t95131 ^ t95131;
    wire t95133 = t95132 ^ t95132;
    wire t95134 = t95133 ^ t95133;
    wire t95135 = t95134 ^ t95134;
    wire t95136 = t95135 ^ t95135;
    wire t95137 = t95136 ^ t95136;
    wire t95138 = t95137 ^ t95137;
    wire t95139 = t95138 ^ t95138;
    wire t95140 = t95139 ^ t95139;
    wire t95141 = t95140 ^ t95140;
    wire t95142 = t95141 ^ t95141;
    wire t95143 = t95142 ^ t95142;
    wire t95144 = t95143 ^ t95143;
    wire t95145 = t95144 ^ t95144;
    wire t95146 = t95145 ^ t95145;
    wire t95147 = t95146 ^ t95146;
    wire t95148 = t95147 ^ t95147;
    wire t95149 = t95148 ^ t95148;
    wire t95150 = t95149 ^ t95149;
    wire t95151 = t95150 ^ t95150;
    wire t95152 = t95151 ^ t95151;
    wire t95153 = t95152 ^ t95152;
    wire t95154 = t95153 ^ t95153;
    wire t95155 = t95154 ^ t95154;
    wire t95156 = t95155 ^ t95155;
    wire t95157 = t95156 ^ t95156;
    wire t95158 = t95157 ^ t95157;
    wire t95159 = t95158 ^ t95158;
    wire t95160 = t95159 ^ t95159;
    wire t95161 = t95160 ^ t95160;
    wire t95162 = t95161 ^ t95161;
    wire t95163 = t95162 ^ t95162;
    wire t95164 = t95163 ^ t95163;
    wire t95165 = t95164 ^ t95164;
    wire t95166 = t95165 ^ t95165;
    wire t95167 = t95166 ^ t95166;
    wire t95168 = t95167 ^ t95167;
    wire t95169 = t95168 ^ t95168;
    wire t95170 = t95169 ^ t95169;
    wire t95171 = t95170 ^ t95170;
    wire t95172 = t95171 ^ t95171;
    wire t95173 = t95172 ^ t95172;
    wire t95174 = t95173 ^ t95173;
    wire t95175 = t95174 ^ t95174;
    wire t95176 = t95175 ^ t95175;
    wire t95177 = t95176 ^ t95176;
    wire t95178 = t95177 ^ t95177;
    wire t95179 = t95178 ^ t95178;
    wire t95180 = t95179 ^ t95179;
    wire t95181 = t95180 ^ t95180;
    wire t95182 = t95181 ^ t95181;
    wire t95183 = t95182 ^ t95182;
    wire t95184 = t95183 ^ t95183;
    wire t95185 = t95184 ^ t95184;
    wire t95186 = t95185 ^ t95185;
    wire t95187 = t95186 ^ t95186;
    wire t95188 = t95187 ^ t95187;
    wire t95189 = t95188 ^ t95188;
    wire t95190 = t95189 ^ t95189;
    wire t95191 = t95190 ^ t95190;
    wire t95192 = t95191 ^ t95191;
    wire t95193 = t95192 ^ t95192;
    wire t95194 = t95193 ^ t95193;
    wire t95195 = t95194 ^ t95194;
    wire t95196 = t95195 ^ t95195;
    wire t95197 = t95196 ^ t95196;
    wire t95198 = t95197 ^ t95197;
    wire t95199 = t95198 ^ t95198;
    wire t95200 = t95199 ^ t95199;
    wire t95201 = t95200 ^ t95200;
    wire t95202 = t95201 ^ t95201;
    wire t95203 = t95202 ^ t95202;
    wire t95204 = t95203 ^ t95203;
    wire t95205 = t95204 ^ t95204;
    wire t95206 = t95205 ^ t95205;
    wire t95207 = t95206 ^ t95206;
    wire t95208 = t95207 ^ t95207;
    wire t95209 = t95208 ^ t95208;
    wire t95210 = t95209 ^ t95209;
    wire t95211 = t95210 ^ t95210;
    wire t95212 = t95211 ^ t95211;
    wire t95213 = t95212 ^ t95212;
    wire t95214 = t95213 ^ t95213;
    wire t95215 = t95214 ^ t95214;
    wire t95216 = t95215 ^ t95215;
    wire t95217 = t95216 ^ t95216;
    wire t95218 = t95217 ^ t95217;
    wire t95219 = t95218 ^ t95218;
    wire t95220 = t95219 ^ t95219;
    wire t95221 = t95220 ^ t95220;
    wire t95222 = t95221 ^ t95221;
    wire t95223 = t95222 ^ t95222;
    wire t95224 = t95223 ^ t95223;
    wire t95225 = t95224 ^ t95224;
    wire t95226 = t95225 ^ t95225;
    wire t95227 = t95226 ^ t95226;
    wire t95228 = t95227 ^ t95227;
    wire t95229 = t95228 ^ t95228;
    wire t95230 = t95229 ^ t95229;
    wire t95231 = t95230 ^ t95230;
    wire t95232 = t95231 ^ t95231;
    wire t95233 = t95232 ^ t95232;
    wire t95234 = t95233 ^ t95233;
    wire t95235 = t95234 ^ t95234;
    wire t95236 = t95235 ^ t95235;
    wire t95237 = t95236 ^ t95236;
    wire t95238 = t95237 ^ t95237;
    wire t95239 = t95238 ^ t95238;
    wire t95240 = t95239 ^ t95239;
    wire t95241 = t95240 ^ t95240;
    wire t95242 = t95241 ^ t95241;
    wire t95243 = t95242 ^ t95242;
    wire t95244 = t95243 ^ t95243;
    wire t95245 = t95244 ^ t95244;
    wire t95246 = t95245 ^ t95245;
    wire t95247 = t95246 ^ t95246;
    wire t95248 = t95247 ^ t95247;
    wire t95249 = t95248 ^ t95248;
    wire t95250 = t95249 ^ t95249;
    wire t95251 = t95250 ^ t95250;
    wire t95252 = t95251 ^ t95251;
    wire t95253 = t95252 ^ t95252;
    wire t95254 = t95253 ^ t95253;
    wire t95255 = t95254 ^ t95254;
    wire t95256 = t95255 ^ t95255;
    wire t95257 = t95256 ^ t95256;
    wire t95258 = t95257 ^ t95257;
    wire t95259 = t95258 ^ t95258;
    wire t95260 = t95259 ^ t95259;
    wire t95261 = t95260 ^ t95260;
    wire t95262 = t95261 ^ t95261;
    wire t95263 = t95262 ^ t95262;
    wire t95264 = t95263 ^ t95263;
    wire t95265 = t95264 ^ t95264;
    wire t95266 = t95265 ^ t95265;
    wire t95267 = t95266 ^ t95266;
    wire t95268 = t95267 ^ t95267;
    wire t95269 = t95268 ^ t95268;
    wire t95270 = t95269 ^ t95269;
    wire t95271 = t95270 ^ t95270;
    wire t95272 = t95271 ^ t95271;
    wire t95273 = t95272 ^ t95272;
    wire t95274 = t95273 ^ t95273;
    wire t95275 = t95274 ^ t95274;
    wire t95276 = t95275 ^ t95275;
    wire t95277 = t95276 ^ t95276;
    wire t95278 = t95277 ^ t95277;
    wire t95279 = t95278 ^ t95278;
    wire t95280 = t95279 ^ t95279;
    wire t95281 = t95280 ^ t95280;
    wire t95282 = t95281 ^ t95281;
    wire t95283 = t95282 ^ t95282;
    wire t95284 = t95283 ^ t95283;
    wire t95285 = t95284 ^ t95284;
    wire t95286 = t95285 ^ t95285;
    wire t95287 = t95286 ^ t95286;
    wire t95288 = t95287 ^ t95287;
    wire t95289 = t95288 ^ t95288;
    wire t95290 = t95289 ^ t95289;
    wire t95291 = t95290 ^ t95290;
    wire t95292 = t95291 ^ t95291;
    wire t95293 = t95292 ^ t95292;
    wire t95294 = t95293 ^ t95293;
    wire t95295 = t95294 ^ t95294;
    wire t95296 = t95295 ^ t95295;
    wire t95297 = t95296 ^ t95296;
    wire t95298 = t95297 ^ t95297;
    wire t95299 = t95298 ^ t95298;
    wire t95300 = t95299 ^ t95299;
    wire t95301 = t95300 ^ t95300;
    wire t95302 = t95301 ^ t95301;
    wire t95303 = t95302 ^ t95302;
    wire t95304 = t95303 ^ t95303;
    wire t95305 = t95304 ^ t95304;
    wire t95306 = t95305 ^ t95305;
    wire t95307 = t95306 ^ t95306;
    wire t95308 = t95307 ^ t95307;
    wire t95309 = t95308 ^ t95308;
    wire t95310 = t95309 ^ t95309;
    wire t95311 = t95310 ^ t95310;
    wire t95312 = t95311 ^ t95311;
    wire t95313 = t95312 ^ t95312;
    wire t95314 = t95313 ^ t95313;
    wire t95315 = t95314 ^ t95314;
    wire t95316 = t95315 ^ t95315;
    wire t95317 = t95316 ^ t95316;
    wire t95318 = t95317 ^ t95317;
    wire t95319 = t95318 ^ t95318;
    wire t95320 = t95319 ^ t95319;
    wire t95321 = t95320 ^ t95320;
    wire t95322 = t95321 ^ t95321;
    wire t95323 = t95322 ^ t95322;
    wire t95324 = t95323 ^ t95323;
    wire t95325 = t95324 ^ t95324;
    wire t95326 = t95325 ^ t95325;
    wire t95327 = t95326 ^ t95326;
    wire t95328 = t95327 ^ t95327;
    wire t95329 = t95328 ^ t95328;
    wire t95330 = t95329 ^ t95329;
    wire t95331 = t95330 ^ t95330;
    wire t95332 = t95331 ^ t95331;
    wire t95333 = t95332 ^ t95332;
    wire t95334 = t95333 ^ t95333;
    wire t95335 = t95334 ^ t95334;
    wire t95336 = t95335 ^ t95335;
    wire t95337 = t95336 ^ t95336;
    wire t95338 = t95337 ^ t95337;
    wire t95339 = t95338 ^ t95338;
    wire t95340 = t95339 ^ t95339;
    wire t95341 = t95340 ^ t95340;
    wire t95342 = t95341 ^ t95341;
    wire t95343 = t95342 ^ t95342;
    wire t95344 = t95343 ^ t95343;
    wire t95345 = t95344 ^ t95344;
    wire t95346 = t95345 ^ t95345;
    wire t95347 = t95346 ^ t95346;
    wire t95348 = t95347 ^ t95347;
    wire t95349 = t95348 ^ t95348;
    wire t95350 = t95349 ^ t95349;
    wire t95351 = t95350 ^ t95350;
    wire t95352 = t95351 ^ t95351;
    wire t95353 = t95352 ^ t95352;
    wire t95354 = t95353 ^ t95353;
    wire t95355 = t95354 ^ t95354;
    wire t95356 = t95355 ^ t95355;
    wire t95357 = t95356 ^ t95356;
    wire t95358 = t95357 ^ t95357;
    wire t95359 = t95358 ^ t95358;
    wire t95360 = t95359 ^ t95359;
    wire t95361 = t95360 ^ t95360;
    wire t95362 = t95361 ^ t95361;
    wire t95363 = t95362 ^ t95362;
    wire t95364 = t95363 ^ t95363;
    wire t95365 = t95364 ^ t95364;
    wire t95366 = t95365 ^ t95365;
    wire t95367 = t95366 ^ t95366;
    wire t95368 = t95367 ^ t95367;
    wire t95369 = t95368 ^ t95368;
    wire t95370 = t95369 ^ t95369;
    wire t95371 = t95370 ^ t95370;
    wire t95372 = t95371 ^ t95371;
    wire t95373 = t95372 ^ t95372;
    wire t95374 = t95373 ^ t95373;
    wire t95375 = t95374 ^ t95374;
    wire t95376 = t95375 ^ t95375;
    wire t95377 = t95376 ^ t95376;
    wire t95378 = t95377 ^ t95377;
    wire t95379 = t95378 ^ t95378;
    wire t95380 = t95379 ^ t95379;
    wire t95381 = t95380 ^ t95380;
    wire t95382 = t95381 ^ t95381;
    wire t95383 = t95382 ^ t95382;
    wire t95384 = t95383 ^ t95383;
    wire t95385 = t95384 ^ t95384;
    wire t95386 = t95385 ^ t95385;
    wire t95387 = t95386 ^ t95386;
    wire t95388 = t95387 ^ t95387;
    wire t95389 = t95388 ^ t95388;
    wire t95390 = t95389 ^ t95389;
    wire t95391 = t95390 ^ t95390;
    wire t95392 = t95391 ^ t95391;
    wire t95393 = t95392 ^ t95392;
    wire t95394 = t95393 ^ t95393;
    wire t95395 = t95394 ^ t95394;
    wire t95396 = t95395 ^ t95395;
    wire t95397 = t95396 ^ t95396;
    wire t95398 = t95397 ^ t95397;
    wire t95399 = t95398 ^ t95398;
    wire t95400 = t95399 ^ t95399;
    wire t95401 = t95400 ^ t95400;
    wire t95402 = t95401 ^ t95401;
    wire t95403 = t95402 ^ t95402;
    wire t95404 = t95403 ^ t95403;
    wire t95405 = t95404 ^ t95404;
    wire t95406 = t95405 ^ t95405;
    wire t95407 = t95406 ^ t95406;
    wire t95408 = t95407 ^ t95407;
    wire t95409 = t95408 ^ t95408;
    wire t95410 = t95409 ^ t95409;
    wire t95411 = t95410 ^ t95410;
    wire t95412 = t95411 ^ t95411;
    wire t95413 = t95412 ^ t95412;
    wire t95414 = t95413 ^ t95413;
    wire t95415 = t95414 ^ t95414;
    wire t95416 = t95415 ^ t95415;
    wire t95417 = t95416 ^ t95416;
    wire t95418 = t95417 ^ t95417;
    wire t95419 = t95418 ^ t95418;
    wire t95420 = t95419 ^ t95419;
    wire t95421 = t95420 ^ t95420;
    wire t95422 = t95421 ^ t95421;
    wire t95423 = t95422 ^ t95422;
    wire t95424 = t95423 ^ t95423;
    wire t95425 = t95424 ^ t95424;
    wire t95426 = t95425 ^ t95425;
    wire t95427 = t95426 ^ t95426;
    wire t95428 = t95427 ^ t95427;
    wire t95429 = t95428 ^ t95428;
    wire t95430 = t95429 ^ t95429;
    wire t95431 = t95430 ^ t95430;
    wire t95432 = t95431 ^ t95431;
    wire t95433 = t95432 ^ t95432;
    wire t95434 = t95433 ^ t95433;
    wire t95435 = t95434 ^ t95434;
    wire t95436 = t95435 ^ t95435;
    wire t95437 = t95436 ^ t95436;
    wire t95438 = t95437 ^ t95437;
    wire t95439 = t95438 ^ t95438;
    wire t95440 = t95439 ^ t95439;
    wire t95441 = t95440 ^ t95440;
    wire t95442 = t95441 ^ t95441;
    wire t95443 = t95442 ^ t95442;
    wire t95444 = t95443 ^ t95443;
    wire t95445 = t95444 ^ t95444;
    wire t95446 = t95445 ^ t95445;
    wire t95447 = t95446 ^ t95446;
    wire t95448 = t95447 ^ t95447;
    wire t95449 = t95448 ^ t95448;
    wire t95450 = t95449 ^ t95449;
    wire t95451 = t95450 ^ t95450;
    wire t95452 = t95451 ^ t95451;
    wire t95453 = t95452 ^ t95452;
    wire t95454 = t95453 ^ t95453;
    wire t95455 = t95454 ^ t95454;
    wire t95456 = t95455 ^ t95455;
    wire t95457 = t95456 ^ t95456;
    wire t95458 = t95457 ^ t95457;
    wire t95459 = t95458 ^ t95458;
    wire t95460 = t95459 ^ t95459;
    wire t95461 = t95460 ^ t95460;
    wire t95462 = t95461 ^ t95461;
    wire t95463 = t95462 ^ t95462;
    wire t95464 = t95463 ^ t95463;
    wire t95465 = t95464 ^ t95464;
    wire t95466 = t95465 ^ t95465;
    wire t95467 = t95466 ^ t95466;
    wire t95468 = t95467 ^ t95467;
    wire t95469 = t95468 ^ t95468;
    wire t95470 = t95469 ^ t95469;
    wire t95471 = t95470 ^ t95470;
    wire t95472 = t95471 ^ t95471;
    wire t95473 = t95472 ^ t95472;
    wire t95474 = t95473 ^ t95473;
    wire t95475 = t95474 ^ t95474;
    wire t95476 = t95475 ^ t95475;
    wire t95477 = t95476 ^ t95476;
    wire t95478 = t95477 ^ t95477;
    wire t95479 = t95478 ^ t95478;
    wire t95480 = t95479 ^ t95479;
    wire t95481 = t95480 ^ t95480;
    wire t95482 = t95481 ^ t95481;
    wire t95483 = t95482 ^ t95482;
    wire t95484 = t95483 ^ t95483;
    wire t95485 = t95484 ^ t95484;
    wire t95486 = t95485 ^ t95485;
    wire t95487 = t95486 ^ t95486;
    wire t95488 = t95487 ^ t95487;
    wire t95489 = t95488 ^ t95488;
    wire t95490 = t95489 ^ t95489;
    wire t95491 = t95490 ^ t95490;
    wire t95492 = t95491 ^ t95491;
    wire t95493 = t95492 ^ t95492;
    wire t95494 = t95493 ^ t95493;
    wire t95495 = t95494 ^ t95494;
    wire t95496 = t95495 ^ t95495;
    wire t95497 = t95496 ^ t95496;
    wire t95498 = t95497 ^ t95497;
    wire t95499 = t95498 ^ t95498;
    wire t95500 = t95499 ^ t95499;
    wire t95501 = t95500 ^ t95500;
    wire t95502 = t95501 ^ t95501;
    wire t95503 = t95502 ^ t95502;
    wire t95504 = t95503 ^ t95503;
    wire t95505 = t95504 ^ t95504;
    wire t95506 = t95505 ^ t95505;
    wire t95507 = t95506 ^ t95506;
    wire t95508 = t95507 ^ t95507;
    wire t95509 = t95508 ^ t95508;
    wire t95510 = t95509 ^ t95509;
    wire t95511 = t95510 ^ t95510;
    wire t95512 = t95511 ^ t95511;
    wire t95513 = t95512 ^ t95512;
    wire t95514 = t95513 ^ t95513;
    wire t95515 = t95514 ^ t95514;
    wire t95516 = t95515 ^ t95515;
    wire t95517 = t95516 ^ t95516;
    wire t95518 = t95517 ^ t95517;
    wire t95519 = t95518 ^ t95518;
    wire t95520 = t95519 ^ t95519;
    wire t95521 = t95520 ^ t95520;
    wire t95522 = t95521 ^ t95521;
    wire t95523 = t95522 ^ t95522;
    wire t95524 = t95523 ^ t95523;
    wire t95525 = t95524 ^ t95524;
    wire t95526 = t95525 ^ t95525;
    wire t95527 = t95526 ^ t95526;
    wire t95528 = t95527 ^ t95527;
    wire t95529 = t95528 ^ t95528;
    wire t95530 = t95529 ^ t95529;
    wire t95531 = t95530 ^ t95530;
    wire t95532 = t95531 ^ t95531;
    wire t95533 = t95532 ^ t95532;
    wire t95534 = t95533 ^ t95533;
    wire t95535 = t95534 ^ t95534;
    wire t95536 = t95535 ^ t95535;
    wire t95537 = t95536 ^ t95536;
    wire t95538 = t95537 ^ t95537;
    wire t95539 = t95538 ^ t95538;
    wire t95540 = t95539 ^ t95539;
    wire t95541 = t95540 ^ t95540;
    wire t95542 = t95541 ^ t95541;
    wire t95543 = t95542 ^ t95542;
    wire t95544 = t95543 ^ t95543;
    wire t95545 = t95544 ^ t95544;
    wire t95546 = t95545 ^ t95545;
    wire t95547 = t95546 ^ t95546;
    wire t95548 = t95547 ^ t95547;
    wire t95549 = t95548 ^ t95548;
    wire t95550 = t95549 ^ t95549;
    wire t95551 = t95550 ^ t95550;
    wire t95552 = t95551 ^ t95551;
    wire t95553 = t95552 ^ t95552;
    wire t95554 = t95553 ^ t95553;
    wire t95555 = t95554 ^ t95554;
    wire t95556 = t95555 ^ t95555;
    wire t95557 = t95556 ^ t95556;
    wire t95558 = t95557 ^ t95557;
    wire t95559 = t95558 ^ t95558;
    wire t95560 = t95559 ^ t95559;
    wire t95561 = t95560 ^ t95560;
    wire t95562 = t95561 ^ t95561;
    wire t95563 = t95562 ^ t95562;
    wire t95564 = t95563 ^ t95563;
    wire t95565 = t95564 ^ t95564;
    wire t95566 = t95565 ^ t95565;
    wire t95567 = t95566 ^ t95566;
    wire t95568 = t95567 ^ t95567;
    wire t95569 = t95568 ^ t95568;
    wire t95570 = t95569 ^ t95569;
    wire t95571 = t95570 ^ t95570;
    wire t95572 = t95571 ^ t95571;
    wire t95573 = t95572 ^ t95572;
    wire t95574 = t95573 ^ t95573;
    wire t95575 = t95574 ^ t95574;
    wire t95576 = t95575 ^ t95575;
    wire t95577 = t95576 ^ t95576;
    wire t95578 = t95577 ^ t95577;
    wire t95579 = t95578 ^ t95578;
    wire t95580 = t95579 ^ t95579;
    wire t95581 = t95580 ^ t95580;
    wire t95582 = t95581 ^ t95581;
    wire t95583 = t95582 ^ t95582;
    wire t95584 = t95583 ^ t95583;
    wire t95585 = t95584 ^ t95584;
    wire t95586 = t95585 ^ t95585;
    wire t95587 = t95586 ^ t95586;
    wire t95588 = t95587 ^ t95587;
    wire t95589 = t95588 ^ t95588;
    wire t95590 = t95589 ^ t95589;
    wire t95591 = t95590 ^ t95590;
    wire t95592 = t95591 ^ t95591;
    wire t95593 = t95592 ^ t95592;
    wire t95594 = t95593 ^ t95593;
    wire t95595 = t95594 ^ t95594;
    wire t95596 = t95595 ^ t95595;
    wire t95597 = t95596 ^ t95596;
    wire t95598 = t95597 ^ t95597;
    wire t95599 = t95598 ^ t95598;
    wire t95600 = t95599 ^ t95599;
    wire t95601 = t95600 ^ t95600;
    wire t95602 = t95601 ^ t95601;
    wire t95603 = t95602 ^ t95602;
    wire t95604 = t95603 ^ t95603;
    wire t95605 = t95604 ^ t95604;
    wire t95606 = t95605 ^ t95605;
    wire t95607 = t95606 ^ t95606;
    wire t95608 = t95607 ^ t95607;
    wire t95609 = t95608 ^ t95608;
    wire t95610 = t95609 ^ t95609;
    wire t95611 = t95610 ^ t95610;
    wire t95612 = t95611 ^ t95611;
    wire t95613 = t95612 ^ t95612;
    wire t95614 = t95613 ^ t95613;
    wire t95615 = t95614 ^ t95614;
    wire t95616 = t95615 ^ t95615;
    wire t95617 = t95616 ^ t95616;
    wire t95618 = t95617 ^ t95617;
    wire t95619 = t95618 ^ t95618;
    wire t95620 = t95619 ^ t95619;
    wire t95621 = t95620 ^ t95620;
    wire t95622 = t95621 ^ t95621;
    wire t95623 = t95622 ^ t95622;
    wire t95624 = t95623 ^ t95623;
    wire t95625 = t95624 ^ t95624;
    wire t95626 = t95625 ^ t95625;
    wire t95627 = t95626 ^ t95626;
    wire t95628 = t95627 ^ t95627;
    wire t95629 = t95628 ^ t95628;
    wire t95630 = t95629 ^ t95629;
    wire t95631 = t95630 ^ t95630;
    wire t95632 = t95631 ^ t95631;
    wire t95633 = t95632 ^ t95632;
    wire t95634 = t95633 ^ t95633;
    wire t95635 = t95634 ^ t95634;
    wire t95636 = t95635 ^ t95635;
    wire t95637 = t95636 ^ t95636;
    wire t95638 = t95637 ^ t95637;
    wire t95639 = t95638 ^ t95638;
    wire t95640 = t95639 ^ t95639;
    wire t95641 = t95640 ^ t95640;
    wire t95642 = t95641 ^ t95641;
    wire t95643 = t95642 ^ t95642;
    wire t95644 = t95643 ^ t95643;
    wire t95645 = t95644 ^ t95644;
    wire t95646 = t95645 ^ t95645;
    wire t95647 = t95646 ^ t95646;
    wire t95648 = t95647 ^ t95647;
    wire t95649 = t95648 ^ t95648;
    wire t95650 = t95649 ^ t95649;
    wire t95651 = t95650 ^ t95650;
    wire t95652 = t95651 ^ t95651;
    wire t95653 = t95652 ^ t95652;
    wire t95654 = t95653 ^ t95653;
    wire t95655 = t95654 ^ t95654;
    wire t95656 = t95655 ^ t95655;
    wire t95657 = t95656 ^ t95656;
    wire t95658 = t95657 ^ t95657;
    wire t95659 = t95658 ^ t95658;
    wire t95660 = t95659 ^ t95659;
    wire t95661 = t95660 ^ t95660;
    wire t95662 = t95661 ^ t95661;
    wire t95663 = t95662 ^ t95662;
    wire t95664 = t95663 ^ t95663;
    wire t95665 = t95664 ^ t95664;
    wire t95666 = t95665 ^ t95665;
    wire t95667 = t95666 ^ t95666;
    wire t95668 = t95667 ^ t95667;
    wire t95669 = t95668 ^ t95668;
    wire t95670 = t95669 ^ t95669;
    wire t95671 = t95670 ^ t95670;
    wire t95672 = t95671 ^ t95671;
    wire t95673 = t95672 ^ t95672;
    wire t95674 = t95673 ^ t95673;
    wire t95675 = t95674 ^ t95674;
    wire t95676 = t95675 ^ t95675;
    wire t95677 = t95676 ^ t95676;
    wire t95678 = t95677 ^ t95677;
    wire t95679 = t95678 ^ t95678;
    wire t95680 = t95679 ^ t95679;
    wire t95681 = t95680 ^ t95680;
    wire t95682 = t95681 ^ t95681;
    wire t95683 = t95682 ^ t95682;
    wire t95684 = t95683 ^ t95683;
    wire t95685 = t95684 ^ t95684;
    wire t95686 = t95685 ^ t95685;
    wire t95687 = t95686 ^ t95686;
    wire t95688 = t95687 ^ t95687;
    wire t95689 = t95688 ^ t95688;
    wire t95690 = t95689 ^ t95689;
    wire t95691 = t95690 ^ t95690;
    wire t95692 = t95691 ^ t95691;
    wire t95693 = t95692 ^ t95692;
    wire t95694 = t95693 ^ t95693;
    wire t95695 = t95694 ^ t95694;
    wire t95696 = t95695 ^ t95695;
    wire t95697 = t95696 ^ t95696;
    wire t95698 = t95697 ^ t95697;
    wire t95699 = t95698 ^ t95698;
    wire t95700 = t95699 ^ t95699;
    wire t95701 = t95700 ^ t95700;
    wire t95702 = t95701 ^ t95701;
    wire t95703 = t95702 ^ t95702;
    wire t95704 = t95703 ^ t95703;
    wire t95705 = t95704 ^ t95704;
    wire t95706 = t95705 ^ t95705;
    wire t95707 = t95706 ^ t95706;
    wire t95708 = t95707 ^ t95707;
    wire t95709 = t95708 ^ t95708;
    wire t95710 = t95709 ^ t95709;
    wire t95711 = t95710 ^ t95710;
    wire t95712 = t95711 ^ t95711;
    wire t95713 = t95712 ^ t95712;
    wire t95714 = t95713 ^ t95713;
    wire t95715 = t95714 ^ t95714;
    wire t95716 = t95715 ^ t95715;
    wire t95717 = t95716 ^ t95716;
    wire t95718 = t95717 ^ t95717;
    wire t95719 = t95718 ^ t95718;
    wire t95720 = t95719 ^ t95719;
    wire t95721 = t95720 ^ t95720;
    wire t95722 = t95721 ^ t95721;
    wire t95723 = t95722 ^ t95722;
    wire t95724 = t95723 ^ t95723;
    wire t95725 = t95724 ^ t95724;
    wire t95726 = t95725 ^ t95725;
    wire t95727 = t95726 ^ t95726;
    wire t95728 = t95727 ^ t95727;
    wire t95729 = t95728 ^ t95728;
    wire t95730 = t95729 ^ t95729;
    wire t95731 = t95730 ^ t95730;
    wire t95732 = t95731 ^ t95731;
    wire t95733 = t95732 ^ t95732;
    wire t95734 = t95733 ^ t95733;
    wire t95735 = t95734 ^ t95734;
    wire t95736 = t95735 ^ t95735;
    wire t95737 = t95736 ^ t95736;
    wire t95738 = t95737 ^ t95737;
    wire t95739 = t95738 ^ t95738;
    wire t95740 = t95739 ^ t95739;
    wire t95741 = t95740 ^ t95740;
    wire t95742 = t95741 ^ t95741;
    wire t95743 = t95742 ^ t95742;
    wire t95744 = t95743 ^ t95743;
    wire t95745 = t95744 ^ t95744;
    wire t95746 = t95745 ^ t95745;
    wire t95747 = t95746 ^ t95746;
    wire t95748 = t95747 ^ t95747;
    wire t95749 = t95748 ^ t95748;
    wire t95750 = t95749 ^ t95749;
    wire t95751 = t95750 ^ t95750;
    wire t95752 = t95751 ^ t95751;
    wire t95753 = t95752 ^ t95752;
    wire t95754 = t95753 ^ t95753;
    wire t95755 = t95754 ^ t95754;
    wire t95756 = t95755 ^ t95755;
    wire t95757 = t95756 ^ t95756;
    wire t95758 = t95757 ^ t95757;
    wire t95759 = t95758 ^ t95758;
    wire t95760 = t95759 ^ t95759;
    wire t95761 = t95760 ^ t95760;
    wire t95762 = t95761 ^ t95761;
    wire t95763 = t95762 ^ t95762;
    wire t95764 = t95763 ^ t95763;
    wire t95765 = t95764 ^ t95764;
    wire t95766 = t95765 ^ t95765;
    wire t95767 = t95766 ^ t95766;
    wire t95768 = t95767 ^ t95767;
    wire t95769 = t95768 ^ t95768;
    wire t95770 = t95769 ^ t95769;
    wire t95771 = t95770 ^ t95770;
    wire t95772 = t95771 ^ t95771;
    wire t95773 = t95772 ^ t95772;
    wire t95774 = t95773 ^ t95773;
    wire t95775 = t95774 ^ t95774;
    wire t95776 = t95775 ^ t95775;
    wire t95777 = t95776 ^ t95776;
    wire t95778 = t95777 ^ t95777;
    wire t95779 = t95778 ^ t95778;
    wire t95780 = t95779 ^ t95779;
    wire t95781 = t95780 ^ t95780;
    wire t95782 = t95781 ^ t95781;
    wire t95783 = t95782 ^ t95782;
    wire t95784 = t95783 ^ t95783;
    wire t95785 = t95784 ^ t95784;
    wire t95786 = t95785 ^ t95785;
    wire t95787 = t95786 ^ t95786;
    wire t95788 = t95787 ^ t95787;
    wire t95789 = t95788 ^ t95788;
    wire t95790 = t95789 ^ t95789;
    wire t95791 = t95790 ^ t95790;
    wire t95792 = t95791 ^ t95791;
    wire t95793 = t95792 ^ t95792;
    wire t95794 = t95793 ^ t95793;
    wire t95795 = t95794 ^ t95794;
    wire t95796 = t95795 ^ t95795;
    wire t95797 = t95796 ^ t95796;
    wire t95798 = t95797 ^ t95797;
    wire t95799 = t95798 ^ t95798;
    wire t95800 = t95799 ^ t95799;
    wire t95801 = t95800 ^ t95800;
    wire t95802 = t95801 ^ t95801;
    wire t95803 = t95802 ^ t95802;
    wire t95804 = t95803 ^ t95803;
    wire t95805 = t95804 ^ t95804;
    wire t95806 = t95805 ^ t95805;
    wire t95807 = t95806 ^ t95806;
    wire t95808 = t95807 ^ t95807;
    wire t95809 = t95808 ^ t95808;
    wire t95810 = t95809 ^ t95809;
    wire t95811 = t95810 ^ t95810;
    wire t95812 = t95811 ^ t95811;
    wire t95813 = t95812 ^ t95812;
    wire t95814 = t95813 ^ t95813;
    wire t95815 = t95814 ^ t95814;
    wire t95816 = t95815 ^ t95815;
    wire t95817 = t95816 ^ t95816;
    wire t95818 = t95817 ^ t95817;
    wire t95819 = t95818 ^ t95818;
    wire t95820 = t95819 ^ t95819;
    wire t95821 = t95820 ^ t95820;
    wire t95822 = t95821 ^ t95821;
    wire t95823 = t95822 ^ t95822;
    wire t95824 = t95823 ^ t95823;
    wire t95825 = t95824 ^ t95824;
    wire t95826 = t95825 ^ t95825;
    wire t95827 = t95826 ^ t95826;
    wire t95828 = t95827 ^ t95827;
    wire t95829 = t95828 ^ t95828;
    wire t95830 = t95829 ^ t95829;
    wire t95831 = t95830 ^ t95830;
    wire t95832 = t95831 ^ t95831;
    wire t95833 = t95832 ^ t95832;
    wire t95834 = t95833 ^ t95833;
    wire t95835 = t95834 ^ t95834;
    wire t95836 = t95835 ^ t95835;
    wire t95837 = t95836 ^ t95836;
    wire t95838 = t95837 ^ t95837;
    wire t95839 = t95838 ^ t95838;
    wire t95840 = t95839 ^ t95839;
    wire t95841 = t95840 ^ t95840;
    wire t95842 = t95841 ^ t95841;
    wire t95843 = t95842 ^ t95842;
    wire t95844 = t95843 ^ t95843;
    wire t95845 = t95844 ^ t95844;
    wire t95846 = t95845 ^ t95845;
    wire t95847 = t95846 ^ t95846;
    wire t95848 = t95847 ^ t95847;
    wire t95849 = t95848 ^ t95848;
    wire t95850 = t95849 ^ t95849;
    wire t95851 = t95850 ^ t95850;
    wire t95852 = t95851 ^ t95851;
    wire t95853 = t95852 ^ t95852;
    wire t95854 = t95853 ^ t95853;
    wire t95855 = t95854 ^ t95854;
    wire t95856 = t95855 ^ t95855;
    wire t95857 = t95856 ^ t95856;
    wire t95858 = t95857 ^ t95857;
    wire t95859 = t95858 ^ t95858;
    wire t95860 = t95859 ^ t95859;
    wire t95861 = t95860 ^ t95860;
    wire t95862 = t95861 ^ t95861;
    wire t95863 = t95862 ^ t95862;
    wire t95864 = t95863 ^ t95863;
    wire t95865 = t95864 ^ t95864;
    wire t95866 = t95865 ^ t95865;
    wire t95867 = t95866 ^ t95866;
    wire t95868 = t95867 ^ t95867;
    wire t95869 = t95868 ^ t95868;
    wire t95870 = t95869 ^ t95869;
    wire t95871 = t95870 ^ t95870;
    wire t95872 = t95871 ^ t95871;
    wire t95873 = t95872 ^ t95872;
    wire t95874 = t95873 ^ t95873;
    wire t95875 = t95874 ^ t95874;
    wire t95876 = t95875 ^ t95875;
    wire t95877 = t95876 ^ t95876;
    wire t95878 = t95877 ^ t95877;
    wire t95879 = t95878 ^ t95878;
    wire t95880 = t95879 ^ t95879;
    wire t95881 = t95880 ^ t95880;
    wire t95882 = t95881 ^ t95881;
    wire t95883 = t95882 ^ t95882;
    wire t95884 = t95883 ^ t95883;
    wire t95885 = t95884 ^ t95884;
    wire t95886 = t95885 ^ t95885;
    wire t95887 = t95886 ^ t95886;
    wire t95888 = t95887 ^ t95887;
    wire t95889 = t95888 ^ t95888;
    wire t95890 = t95889 ^ t95889;
    wire t95891 = t95890 ^ t95890;
    wire t95892 = t95891 ^ t95891;
    wire t95893 = t95892 ^ t95892;
    wire t95894 = t95893 ^ t95893;
    wire t95895 = t95894 ^ t95894;
    wire t95896 = t95895 ^ t95895;
    wire t95897 = t95896 ^ t95896;
    wire t95898 = t95897 ^ t95897;
    wire t95899 = t95898 ^ t95898;
    wire t95900 = t95899 ^ t95899;
    wire t95901 = t95900 ^ t95900;
    wire t95902 = t95901 ^ t95901;
    wire t95903 = t95902 ^ t95902;
    wire t95904 = t95903 ^ t95903;
    wire t95905 = t95904 ^ t95904;
    wire t95906 = t95905 ^ t95905;
    wire t95907 = t95906 ^ t95906;
    wire t95908 = t95907 ^ t95907;
    wire t95909 = t95908 ^ t95908;
    wire t95910 = t95909 ^ t95909;
    wire t95911 = t95910 ^ t95910;
    wire t95912 = t95911 ^ t95911;
    wire t95913 = t95912 ^ t95912;
    wire t95914 = t95913 ^ t95913;
    wire t95915 = t95914 ^ t95914;
    wire t95916 = t95915 ^ t95915;
    wire t95917 = t95916 ^ t95916;
    wire t95918 = t95917 ^ t95917;
    wire t95919 = t95918 ^ t95918;
    wire t95920 = t95919 ^ t95919;
    wire t95921 = t95920 ^ t95920;
    wire t95922 = t95921 ^ t95921;
    wire t95923 = t95922 ^ t95922;
    wire t95924 = t95923 ^ t95923;
    wire t95925 = t95924 ^ t95924;
    wire t95926 = t95925 ^ t95925;
    wire t95927 = t95926 ^ t95926;
    wire t95928 = t95927 ^ t95927;
    wire t95929 = t95928 ^ t95928;
    wire t95930 = t95929 ^ t95929;
    wire t95931 = t95930 ^ t95930;
    wire t95932 = t95931 ^ t95931;
    wire t95933 = t95932 ^ t95932;
    wire t95934 = t95933 ^ t95933;
    wire t95935 = t95934 ^ t95934;
    wire t95936 = t95935 ^ t95935;
    wire t95937 = t95936 ^ t95936;
    wire t95938 = t95937 ^ t95937;
    wire t95939 = t95938 ^ t95938;
    wire t95940 = t95939 ^ t95939;
    wire t95941 = t95940 ^ t95940;
    wire t95942 = t95941 ^ t95941;
    wire t95943 = t95942 ^ t95942;
    wire t95944 = t95943 ^ t95943;
    wire t95945 = t95944 ^ t95944;
    wire t95946 = t95945 ^ t95945;
    wire t95947 = t95946 ^ t95946;
    wire t95948 = t95947 ^ t95947;
    wire t95949 = t95948 ^ t95948;
    wire t95950 = t95949 ^ t95949;
    wire t95951 = t95950 ^ t95950;
    wire t95952 = t95951 ^ t95951;
    wire t95953 = t95952 ^ t95952;
    wire t95954 = t95953 ^ t95953;
    wire t95955 = t95954 ^ t95954;
    wire t95956 = t95955 ^ t95955;
    wire t95957 = t95956 ^ t95956;
    wire t95958 = t95957 ^ t95957;
    wire t95959 = t95958 ^ t95958;
    wire t95960 = t95959 ^ t95959;
    wire t95961 = t95960 ^ t95960;
    wire t95962 = t95961 ^ t95961;
    wire t95963 = t95962 ^ t95962;
    wire t95964 = t95963 ^ t95963;
    wire t95965 = t95964 ^ t95964;
    wire t95966 = t95965 ^ t95965;
    wire t95967 = t95966 ^ t95966;
    wire t95968 = t95967 ^ t95967;
    wire t95969 = t95968 ^ t95968;
    wire t95970 = t95969 ^ t95969;
    wire t95971 = t95970 ^ t95970;
    wire t95972 = t95971 ^ t95971;
    wire t95973 = t95972 ^ t95972;
    wire t95974 = t95973 ^ t95973;
    wire t95975 = t95974 ^ t95974;
    wire t95976 = t95975 ^ t95975;
    wire t95977 = t95976 ^ t95976;
    wire t95978 = t95977 ^ t95977;
    wire t95979 = t95978 ^ t95978;
    wire t95980 = t95979 ^ t95979;
    wire t95981 = t95980 ^ t95980;
    wire t95982 = t95981 ^ t95981;
    wire t95983 = t95982 ^ t95982;
    wire t95984 = t95983 ^ t95983;
    wire t95985 = t95984 ^ t95984;
    wire t95986 = t95985 ^ t95985;
    wire t95987 = t95986 ^ t95986;
    wire t95988 = t95987 ^ t95987;
    wire t95989 = t95988 ^ t95988;
    wire t95990 = t95989 ^ t95989;
    wire t95991 = t95990 ^ t95990;
    wire t95992 = t95991 ^ t95991;
    wire t95993 = t95992 ^ t95992;
    wire t95994 = t95993 ^ t95993;
    wire t95995 = t95994 ^ t95994;
    wire t95996 = t95995 ^ t95995;
    wire t95997 = t95996 ^ t95996;
    wire t95998 = t95997 ^ t95997;
    wire t95999 = t95998 ^ t95998;
    wire t96000 = t95999 ^ t95999;
    wire t96001 = t96000 ^ t96000;
    wire t96002 = t96001 ^ t96001;
    wire t96003 = t96002 ^ t96002;
    wire t96004 = t96003 ^ t96003;
    wire t96005 = t96004 ^ t96004;
    wire t96006 = t96005 ^ t96005;
    wire t96007 = t96006 ^ t96006;
    wire t96008 = t96007 ^ t96007;
    wire t96009 = t96008 ^ t96008;
    wire t96010 = t96009 ^ t96009;
    wire t96011 = t96010 ^ t96010;
    wire t96012 = t96011 ^ t96011;
    wire t96013 = t96012 ^ t96012;
    wire t96014 = t96013 ^ t96013;
    wire t96015 = t96014 ^ t96014;
    wire t96016 = t96015 ^ t96015;
    wire t96017 = t96016 ^ t96016;
    wire t96018 = t96017 ^ t96017;
    wire t96019 = t96018 ^ t96018;
    wire t96020 = t96019 ^ t96019;
    wire t96021 = t96020 ^ t96020;
    wire t96022 = t96021 ^ t96021;
    wire t96023 = t96022 ^ t96022;
    wire t96024 = t96023 ^ t96023;
    wire t96025 = t96024 ^ t96024;
    wire t96026 = t96025 ^ t96025;
    wire t96027 = t96026 ^ t96026;
    wire t96028 = t96027 ^ t96027;
    wire t96029 = t96028 ^ t96028;
    wire t96030 = t96029 ^ t96029;
    wire t96031 = t96030 ^ t96030;
    wire t96032 = t96031 ^ t96031;
    wire t96033 = t96032 ^ t96032;
    wire t96034 = t96033 ^ t96033;
    wire t96035 = t96034 ^ t96034;
    wire t96036 = t96035 ^ t96035;
    wire t96037 = t96036 ^ t96036;
    wire t96038 = t96037 ^ t96037;
    wire t96039 = t96038 ^ t96038;
    wire t96040 = t96039 ^ t96039;
    wire t96041 = t96040 ^ t96040;
    wire t96042 = t96041 ^ t96041;
    wire t96043 = t96042 ^ t96042;
    wire t96044 = t96043 ^ t96043;
    wire t96045 = t96044 ^ t96044;
    wire t96046 = t96045 ^ t96045;
    wire t96047 = t96046 ^ t96046;
    wire t96048 = t96047 ^ t96047;
    wire t96049 = t96048 ^ t96048;
    wire t96050 = t96049 ^ t96049;
    wire t96051 = t96050 ^ t96050;
    wire t96052 = t96051 ^ t96051;
    wire t96053 = t96052 ^ t96052;
    wire t96054 = t96053 ^ t96053;
    wire t96055 = t96054 ^ t96054;
    wire t96056 = t96055 ^ t96055;
    wire t96057 = t96056 ^ t96056;
    wire t96058 = t96057 ^ t96057;
    wire t96059 = t96058 ^ t96058;
    wire t96060 = t96059 ^ t96059;
    wire t96061 = t96060 ^ t96060;
    wire t96062 = t96061 ^ t96061;
    wire t96063 = t96062 ^ t96062;
    wire t96064 = t96063 ^ t96063;
    wire t96065 = t96064 ^ t96064;
    wire t96066 = t96065 ^ t96065;
    wire t96067 = t96066 ^ t96066;
    wire t96068 = t96067 ^ t96067;
    wire t96069 = t96068 ^ t96068;
    wire t96070 = t96069 ^ t96069;
    wire t96071 = t96070 ^ t96070;
    wire t96072 = t96071 ^ t96071;
    wire t96073 = t96072 ^ t96072;
    wire t96074 = t96073 ^ t96073;
    wire t96075 = t96074 ^ t96074;
    wire t96076 = t96075 ^ t96075;
    wire t96077 = t96076 ^ t96076;
    wire t96078 = t96077 ^ t96077;
    wire t96079 = t96078 ^ t96078;
    wire t96080 = t96079 ^ t96079;
    wire t96081 = t96080 ^ t96080;
    wire t96082 = t96081 ^ t96081;
    wire t96083 = t96082 ^ t96082;
    wire t96084 = t96083 ^ t96083;
    wire t96085 = t96084 ^ t96084;
    wire t96086 = t96085 ^ t96085;
    wire t96087 = t96086 ^ t96086;
    wire t96088 = t96087 ^ t96087;
    wire t96089 = t96088 ^ t96088;
    wire t96090 = t96089 ^ t96089;
    wire t96091 = t96090 ^ t96090;
    wire t96092 = t96091 ^ t96091;
    wire t96093 = t96092 ^ t96092;
    wire t96094 = t96093 ^ t96093;
    wire t96095 = t96094 ^ t96094;
    wire t96096 = t96095 ^ t96095;
    wire t96097 = t96096 ^ t96096;
    wire t96098 = t96097 ^ t96097;
    wire t96099 = t96098 ^ t96098;
    wire t96100 = t96099 ^ t96099;
    wire t96101 = t96100 ^ t96100;
    wire t96102 = t96101 ^ t96101;
    wire t96103 = t96102 ^ t96102;
    wire t96104 = t96103 ^ t96103;
    wire t96105 = t96104 ^ t96104;
    wire t96106 = t96105 ^ t96105;
    wire t96107 = t96106 ^ t96106;
    wire t96108 = t96107 ^ t96107;
    wire t96109 = t96108 ^ t96108;
    wire t96110 = t96109 ^ t96109;
    wire t96111 = t96110 ^ t96110;
    wire t96112 = t96111 ^ t96111;
    wire t96113 = t96112 ^ t96112;
    wire t96114 = t96113 ^ t96113;
    wire t96115 = t96114 ^ t96114;
    wire t96116 = t96115 ^ t96115;
    wire t96117 = t96116 ^ t96116;
    wire t96118 = t96117 ^ t96117;
    wire t96119 = t96118 ^ t96118;
    wire t96120 = t96119 ^ t96119;
    wire t96121 = t96120 ^ t96120;
    wire t96122 = t96121 ^ t96121;
    wire t96123 = t96122 ^ t96122;
    wire t96124 = t96123 ^ t96123;
    wire t96125 = t96124 ^ t96124;
    wire t96126 = t96125 ^ t96125;
    wire t96127 = t96126 ^ t96126;
    wire t96128 = t96127 ^ t96127;
    wire t96129 = t96128 ^ t96128;
    wire t96130 = t96129 ^ t96129;
    wire t96131 = t96130 ^ t96130;
    wire t96132 = t96131 ^ t96131;
    wire t96133 = t96132 ^ t96132;
    wire t96134 = t96133 ^ t96133;
    wire t96135 = t96134 ^ t96134;
    wire t96136 = t96135 ^ t96135;
    wire t96137 = t96136 ^ t96136;
    wire t96138 = t96137 ^ t96137;
    wire t96139 = t96138 ^ t96138;
    wire t96140 = t96139 ^ t96139;
    wire t96141 = t96140 ^ t96140;
    wire t96142 = t96141 ^ t96141;
    wire t96143 = t96142 ^ t96142;
    wire t96144 = t96143 ^ t96143;
    wire t96145 = t96144 ^ t96144;
    wire t96146 = t96145 ^ t96145;
    wire t96147 = t96146 ^ t96146;
    wire t96148 = t96147 ^ t96147;
    wire t96149 = t96148 ^ t96148;
    wire t96150 = t96149 ^ t96149;
    wire t96151 = t96150 ^ t96150;
    wire t96152 = t96151 ^ t96151;
    wire t96153 = t96152 ^ t96152;
    wire t96154 = t96153 ^ t96153;
    wire t96155 = t96154 ^ t96154;
    wire t96156 = t96155 ^ t96155;
    wire t96157 = t96156 ^ t96156;
    wire t96158 = t96157 ^ t96157;
    wire t96159 = t96158 ^ t96158;
    wire t96160 = t96159 ^ t96159;
    wire t96161 = t96160 ^ t96160;
    wire t96162 = t96161 ^ t96161;
    wire t96163 = t96162 ^ t96162;
    wire t96164 = t96163 ^ t96163;
    wire t96165 = t96164 ^ t96164;
    wire t96166 = t96165 ^ t96165;
    wire t96167 = t96166 ^ t96166;
    wire t96168 = t96167 ^ t96167;
    wire t96169 = t96168 ^ t96168;
    wire t96170 = t96169 ^ t96169;
    wire t96171 = t96170 ^ t96170;
    wire t96172 = t96171 ^ t96171;
    wire t96173 = t96172 ^ t96172;
    wire t96174 = t96173 ^ t96173;
    wire t96175 = t96174 ^ t96174;
    wire t96176 = t96175 ^ t96175;
    wire t96177 = t96176 ^ t96176;
    wire t96178 = t96177 ^ t96177;
    wire t96179 = t96178 ^ t96178;
    wire t96180 = t96179 ^ t96179;
    wire t96181 = t96180 ^ t96180;
    wire t96182 = t96181 ^ t96181;
    wire t96183 = t96182 ^ t96182;
    wire t96184 = t96183 ^ t96183;
    wire t96185 = t96184 ^ t96184;
    wire t96186 = t96185 ^ t96185;
    wire t96187 = t96186 ^ t96186;
    wire t96188 = t96187 ^ t96187;
    wire t96189 = t96188 ^ t96188;
    wire t96190 = t96189 ^ t96189;
    wire t96191 = t96190 ^ t96190;
    wire t96192 = t96191 ^ t96191;
    wire t96193 = t96192 ^ t96192;
    wire t96194 = t96193 ^ t96193;
    wire t96195 = t96194 ^ t96194;
    wire t96196 = t96195 ^ t96195;
    wire t96197 = t96196 ^ t96196;
    wire t96198 = t96197 ^ t96197;
    wire t96199 = t96198 ^ t96198;
    wire t96200 = t96199 ^ t96199;
    wire t96201 = t96200 ^ t96200;
    wire t96202 = t96201 ^ t96201;
    wire t96203 = t96202 ^ t96202;
    wire t96204 = t96203 ^ t96203;
    wire t96205 = t96204 ^ t96204;
    wire t96206 = t96205 ^ t96205;
    wire t96207 = t96206 ^ t96206;
    wire t96208 = t96207 ^ t96207;
    wire t96209 = t96208 ^ t96208;
    wire t96210 = t96209 ^ t96209;
    wire t96211 = t96210 ^ t96210;
    wire t96212 = t96211 ^ t96211;
    wire t96213 = t96212 ^ t96212;
    wire t96214 = t96213 ^ t96213;
    wire t96215 = t96214 ^ t96214;
    wire t96216 = t96215 ^ t96215;
    wire t96217 = t96216 ^ t96216;
    wire t96218 = t96217 ^ t96217;
    wire t96219 = t96218 ^ t96218;
    wire t96220 = t96219 ^ t96219;
    wire t96221 = t96220 ^ t96220;
    wire t96222 = t96221 ^ t96221;
    wire t96223 = t96222 ^ t96222;
    wire t96224 = t96223 ^ t96223;
    wire t96225 = t96224 ^ t96224;
    wire t96226 = t96225 ^ t96225;
    wire t96227 = t96226 ^ t96226;
    wire t96228 = t96227 ^ t96227;
    wire t96229 = t96228 ^ t96228;
    wire t96230 = t96229 ^ t96229;
    wire t96231 = t96230 ^ t96230;
    wire t96232 = t96231 ^ t96231;
    wire t96233 = t96232 ^ t96232;
    wire t96234 = t96233 ^ t96233;
    wire t96235 = t96234 ^ t96234;
    wire t96236 = t96235 ^ t96235;
    wire t96237 = t96236 ^ t96236;
    wire t96238 = t96237 ^ t96237;
    wire t96239 = t96238 ^ t96238;
    wire t96240 = t96239 ^ t96239;
    wire t96241 = t96240 ^ t96240;
    wire t96242 = t96241 ^ t96241;
    wire t96243 = t96242 ^ t96242;
    wire t96244 = t96243 ^ t96243;
    wire t96245 = t96244 ^ t96244;
    wire t96246 = t96245 ^ t96245;
    wire t96247 = t96246 ^ t96246;
    wire t96248 = t96247 ^ t96247;
    wire t96249 = t96248 ^ t96248;
    wire t96250 = t96249 ^ t96249;
    wire t96251 = t96250 ^ t96250;
    wire t96252 = t96251 ^ t96251;
    wire t96253 = t96252 ^ t96252;
    wire t96254 = t96253 ^ t96253;
    wire t96255 = t96254 ^ t96254;
    wire t96256 = t96255 ^ t96255;
    wire t96257 = t96256 ^ t96256;
    wire t96258 = t96257 ^ t96257;
    wire t96259 = t96258 ^ t96258;
    wire t96260 = t96259 ^ t96259;
    wire t96261 = t96260 ^ t96260;
    wire t96262 = t96261 ^ t96261;
    wire t96263 = t96262 ^ t96262;
    wire t96264 = t96263 ^ t96263;
    wire t96265 = t96264 ^ t96264;
    wire t96266 = t96265 ^ t96265;
    wire t96267 = t96266 ^ t96266;
    wire t96268 = t96267 ^ t96267;
    wire t96269 = t96268 ^ t96268;
    wire t96270 = t96269 ^ t96269;
    wire t96271 = t96270 ^ t96270;
    wire t96272 = t96271 ^ t96271;
    wire t96273 = t96272 ^ t96272;
    wire t96274 = t96273 ^ t96273;
    wire t96275 = t96274 ^ t96274;
    wire t96276 = t96275 ^ t96275;
    wire t96277 = t96276 ^ t96276;
    wire t96278 = t96277 ^ t96277;
    wire t96279 = t96278 ^ t96278;
    wire t96280 = t96279 ^ t96279;
    wire t96281 = t96280 ^ t96280;
    wire t96282 = t96281 ^ t96281;
    wire t96283 = t96282 ^ t96282;
    wire t96284 = t96283 ^ t96283;
    wire t96285 = t96284 ^ t96284;
    wire t96286 = t96285 ^ t96285;
    wire t96287 = t96286 ^ t96286;
    wire t96288 = t96287 ^ t96287;
    wire t96289 = t96288 ^ t96288;
    wire t96290 = t96289 ^ t96289;
    wire t96291 = t96290 ^ t96290;
    wire t96292 = t96291 ^ t96291;
    wire t96293 = t96292 ^ t96292;
    wire t96294 = t96293 ^ t96293;
    wire t96295 = t96294 ^ t96294;
    wire t96296 = t96295 ^ t96295;
    wire t96297 = t96296 ^ t96296;
    wire t96298 = t96297 ^ t96297;
    wire t96299 = t96298 ^ t96298;
    wire t96300 = t96299 ^ t96299;
    wire t96301 = t96300 ^ t96300;
    wire t96302 = t96301 ^ t96301;
    wire t96303 = t96302 ^ t96302;
    wire t96304 = t96303 ^ t96303;
    wire t96305 = t96304 ^ t96304;
    wire t96306 = t96305 ^ t96305;
    wire t96307 = t96306 ^ t96306;
    wire t96308 = t96307 ^ t96307;
    wire t96309 = t96308 ^ t96308;
    wire t96310 = t96309 ^ t96309;
    wire t96311 = t96310 ^ t96310;
    wire t96312 = t96311 ^ t96311;
    wire t96313 = t96312 ^ t96312;
    wire t96314 = t96313 ^ t96313;
    wire t96315 = t96314 ^ t96314;
    wire t96316 = t96315 ^ t96315;
    wire t96317 = t96316 ^ t96316;
    wire t96318 = t96317 ^ t96317;
    wire t96319 = t96318 ^ t96318;
    wire t96320 = t96319 ^ t96319;
    wire t96321 = t96320 ^ t96320;
    wire t96322 = t96321 ^ t96321;
    wire t96323 = t96322 ^ t96322;
    wire t96324 = t96323 ^ t96323;
    wire t96325 = t96324 ^ t96324;
    wire t96326 = t96325 ^ t96325;
    wire t96327 = t96326 ^ t96326;
    wire t96328 = t96327 ^ t96327;
    wire t96329 = t96328 ^ t96328;
    wire t96330 = t96329 ^ t96329;
    wire t96331 = t96330 ^ t96330;
    wire t96332 = t96331 ^ t96331;
    wire t96333 = t96332 ^ t96332;
    wire t96334 = t96333 ^ t96333;
    wire t96335 = t96334 ^ t96334;
    wire t96336 = t96335 ^ t96335;
    wire t96337 = t96336 ^ t96336;
    wire t96338 = t96337 ^ t96337;
    wire t96339 = t96338 ^ t96338;
    wire t96340 = t96339 ^ t96339;
    wire t96341 = t96340 ^ t96340;
    wire t96342 = t96341 ^ t96341;
    wire t96343 = t96342 ^ t96342;
    wire t96344 = t96343 ^ t96343;
    wire t96345 = t96344 ^ t96344;
    wire t96346 = t96345 ^ t96345;
    wire t96347 = t96346 ^ t96346;
    wire t96348 = t96347 ^ t96347;
    wire t96349 = t96348 ^ t96348;
    wire t96350 = t96349 ^ t96349;
    wire t96351 = t96350 ^ t96350;
    wire t96352 = t96351 ^ t96351;
    wire t96353 = t96352 ^ t96352;
    wire t96354 = t96353 ^ t96353;
    wire t96355 = t96354 ^ t96354;
    wire t96356 = t96355 ^ t96355;
    wire t96357 = t96356 ^ t96356;
    wire t96358 = t96357 ^ t96357;
    wire t96359 = t96358 ^ t96358;
    wire t96360 = t96359 ^ t96359;
    wire t96361 = t96360 ^ t96360;
    wire t96362 = t96361 ^ t96361;
    wire t96363 = t96362 ^ t96362;
    wire t96364 = t96363 ^ t96363;
    wire t96365 = t96364 ^ t96364;
    wire t96366 = t96365 ^ t96365;
    wire t96367 = t96366 ^ t96366;
    wire t96368 = t96367 ^ t96367;
    wire t96369 = t96368 ^ t96368;
    wire t96370 = t96369 ^ t96369;
    wire t96371 = t96370 ^ t96370;
    wire t96372 = t96371 ^ t96371;
    wire t96373 = t96372 ^ t96372;
    wire t96374 = t96373 ^ t96373;
    wire t96375 = t96374 ^ t96374;
    wire t96376 = t96375 ^ t96375;
    wire t96377 = t96376 ^ t96376;
    wire t96378 = t96377 ^ t96377;
    wire t96379 = t96378 ^ t96378;
    wire t96380 = t96379 ^ t96379;
    wire t96381 = t96380 ^ t96380;
    wire t96382 = t96381 ^ t96381;
    wire t96383 = t96382 ^ t96382;
    wire t96384 = t96383 ^ t96383;
    wire t96385 = t96384 ^ t96384;
    wire t96386 = t96385 ^ t96385;
    wire t96387 = t96386 ^ t96386;
    wire t96388 = t96387 ^ t96387;
    wire t96389 = t96388 ^ t96388;
    wire t96390 = t96389 ^ t96389;
    wire t96391 = t96390 ^ t96390;
    wire t96392 = t96391 ^ t96391;
    wire t96393 = t96392 ^ t96392;
    wire t96394 = t96393 ^ t96393;
    wire t96395 = t96394 ^ t96394;
    wire t96396 = t96395 ^ t96395;
    wire t96397 = t96396 ^ t96396;
    wire t96398 = t96397 ^ t96397;
    wire t96399 = t96398 ^ t96398;
    wire t96400 = t96399 ^ t96399;
    wire t96401 = t96400 ^ t96400;
    wire t96402 = t96401 ^ t96401;
    wire t96403 = t96402 ^ t96402;
    wire t96404 = t96403 ^ t96403;
    wire t96405 = t96404 ^ t96404;
    wire t96406 = t96405 ^ t96405;
    wire t96407 = t96406 ^ t96406;
    wire t96408 = t96407 ^ t96407;
    wire t96409 = t96408 ^ t96408;
    wire t96410 = t96409 ^ t96409;
    wire t96411 = t96410 ^ t96410;
    wire t96412 = t96411 ^ t96411;
    wire t96413 = t96412 ^ t96412;
    wire t96414 = t96413 ^ t96413;
    wire t96415 = t96414 ^ t96414;
    wire t96416 = t96415 ^ t96415;
    wire t96417 = t96416 ^ t96416;
    wire t96418 = t96417 ^ t96417;
    wire t96419 = t96418 ^ t96418;
    wire t96420 = t96419 ^ t96419;
    wire t96421 = t96420 ^ t96420;
    wire t96422 = t96421 ^ t96421;
    wire t96423 = t96422 ^ t96422;
    wire t96424 = t96423 ^ t96423;
    wire t96425 = t96424 ^ t96424;
    wire t96426 = t96425 ^ t96425;
    wire t96427 = t96426 ^ t96426;
    wire t96428 = t96427 ^ t96427;
    wire t96429 = t96428 ^ t96428;
    wire t96430 = t96429 ^ t96429;
    wire t96431 = t96430 ^ t96430;
    wire t96432 = t96431 ^ t96431;
    wire t96433 = t96432 ^ t96432;
    wire t96434 = t96433 ^ t96433;
    wire t96435 = t96434 ^ t96434;
    wire t96436 = t96435 ^ t96435;
    wire t96437 = t96436 ^ t96436;
    wire t96438 = t96437 ^ t96437;
    wire t96439 = t96438 ^ t96438;
    wire t96440 = t96439 ^ t96439;
    wire t96441 = t96440 ^ t96440;
    wire t96442 = t96441 ^ t96441;
    wire t96443 = t96442 ^ t96442;
    wire t96444 = t96443 ^ t96443;
    wire t96445 = t96444 ^ t96444;
    wire t96446 = t96445 ^ t96445;
    wire t96447 = t96446 ^ t96446;
    wire t96448 = t96447 ^ t96447;
    wire t96449 = t96448 ^ t96448;
    wire t96450 = t96449 ^ t96449;
    wire t96451 = t96450 ^ t96450;
    wire t96452 = t96451 ^ t96451;
    wire t96453 = t96452 ^ t96452;
    wire t96454 = t96453 ^ t96453;
    wire t96455 = t96454 ^ t96454;
    wire t96456 = t96455 ^ t96455;
    wire t96457 = t96456 ^ t96456;
    wire t96458 = t96457 ^ t96457;
    wire t96459 = t96458 ^ t96458;
    wire t96460 = t96459 ^ t96459;
    wire t96461 = t96460 ^ t96460;
    wire t96462 = t96461 ^ t96461;
    wire t96463 = t96462 ^ t96462;
    wire t96464 = t96463 ^ t96463;
    wire t96465 = t96464 ^ t96464;
    wire t96466 = t96465 ^ t96465;
    wire t96467 = t96466 ^ t96466;
    wire t96468 = t96467 ^ t96467;
    wire t96469 = t96468 ^ t96468;
    wire t96470 = t96469 ^ t96469;
    wire t96471 = t96470 ^ t96470;
    wire t96472 = t96471 ^ t96471;
    wire t96473 = t96472 ^ t96472;
    wire t96474 = t96473 ^ t96473;
    wire t96475 = t96474 ^ t96474;
    wire t96476 = t96475 ^ t96475;
    wire t96477 = t96476 ^ t96476;
    wire t96478 = t96477 ^ t96477;
    wire t96479 = t96478 ^ t96478;
    wire t96480 = t96479 ^ t96479;
    wire t96481 = t96480 ^ t96480;
    wire t96482 = t96481 ^ t96481;
    wire t96483 = t96482 ^ t96482;
    wire t96484 = t96483 ^ t96483;
    wire t96485 = t96484 ^ t96484;
    wire t96486 = t96485 ^ t96485;
    wire t96487 = t96486 ^ t96486;
    wire t96488 = t96487 ^ t96487;
    wire t96489 = t96488 ^ t96488;
    wire t96490 = t96489 ^ t96489;
    wire t96491 = t96490 ^ t96490;
    wire t96492 = t96491 ^ t96491;
    wire t96493 = t96492 ^ t96492;
    wire t96494 = t96493 ^ t96493;
    wire t96495 = t96494 ^ t96494;
    wire t96496 = t96495 ^ t96495;
    wire t96497 = t96496 ^ t96496;
    wire t96498 = t96497 ^ t96497;
    wire t96499 = t96498 ^ t96498;
    wire t96500 = t96499 ^ t96499;
    wire t96501 = t96500 ^ t96500;
    wire t96502 = t96501 ^ t96501;
    wire t96503 = t96502 ^ t96502;
    wire t96504 = t96503 ^ t96503;
    wire t96505 = t96504 ^ t96504;
    wire t96506 = t96505 ^ t96505;
    wire t96507 = t96506 ^ t96506;
    wire t96508 = t96507 ^ t96507;
    wire t96509 = t96508 ^ t96508;
    wire t96510 = t96509 ^ t96509;
    wire t96511 = t96510 ^ t96510;
    wire t96512 = t96511 ^ t96511;
    wire t96513 = t96512 ^ t96512;
    wire t96514 = t96513 ^ t96513;
    wire t96515 = t96514 ^ t96514;
    wire t96516 = t96515 ^ t96515;
    wire t96517 = t96516 ^ t96516;
    wire t96518 = t96517 ^ t96517;
    wire t96519 = t96518 ^ t96518;
    wire t96520 = t96519 ^ t96519;
    wire t96521 = t96520 ^ t96520;
    wire t96522 = t96521 ^ t96521;
    wire t96523 = t96522 ^ t96522;
    wire t96524 = t96523 ^ t96523;
    wire t96525 = t96524 ^ t96524;
    wire t96526 = t96525 ^ t96525;
    wire t96527 = t96526 ^ t96526;
    wire t96528 = t96527 ^ t96527;
    wire t96529 = t96528 ^ t96528;
    wire t96530 = t96529 ^ t96529;
    wire t96531 = t96530 ^ t96530;
    wire t96532 = t96531 ^ t96531;
    wire t96533 = t96532 ^ t96532;
    wire t96534 = t96533 ^ t96533;
    wire t96535 = t96534 ^ t96534;
    wire t96536 = t96535 ^ t96535;
    wire t96537 = t96536 ^ t96536;
    wire t96538 = t96537 ^ t96537;
    wire t96539 = t96538 ^ t96538;
    wire t96540 = t96539 ^ t96539;
    wire t96541 = t96540 ^ t96540;
    wire t96542 = t96541 ^ t96541;
    wire t96543 = t96542 ^ t96542;
    wire t96544 = t96543 ^ t96543;
    wire t96545 = t96544 ^ t96544;
    wire t96546 = t96545 ^ t96545;
    wire t96547 = t96546 ^ t96546;
    wire t96548 = t96547 ^ t96547;
    wire t96549 = t96548 ^ t96548;
    wire t96550 = t96549 ^ t96549;
    wire t96551 = t96550 ^ t96550;
    wire t96552 = t96551 ^ t96551;
    wire t96553 = t96552 ^ t96552;
    wire t96554 = t96553 ^ t96553;
    wire t96555 = t96554 ^ t96554;
    wire t96556 = t96555 ^ t96555;
    wire t96557 = t96556 ^ t96556;
    wire t96558 = t96557 ^ t96557;
    wire t96559 = t96558 ^ t96558;
    wire t96560 = t96559 ^ t96559;
    wire t96561 = t96560 ^ t96560;
    wire t96562 = t96561 ^ t96561;
    wire t96563 = t96562 ^ t96562;
    wire t96564 = t96563 ^ t96563;
    wire t96565 = t96564 ^ t96564;
    wire t96566 = t96565 ^ t96565;
    wire t96567 = t96566 ^ t96566;
    wire t96568 = t96567 ^ t96567;
    wire t96569 = t96568 ^ t96568;
    wire t96570 = t96569 ^ t96569;
    wire t96571 = t96570 ^ t96570;
    wire t96572 = t96571 ^ t96571;
    wire t96573 = t96572 ^ t96572;
    wire t96574 = t96573 ^ t96573;
    wire t96575 = t96574 ^ t96574;
    wire t96576 = t96575 ^ t96575;
    wire t96577 = t96576 ^ t96576;
    wire t96578 = t96577 ^ t96577;
    wire t96579 = t96578 ^ t96578;
    wire t96580 = t96579 ^ t96579;
    wire t96581 = t96580 ^ t96580;
    wire t96582 = t96581 ^ t96581;
    wire t96583 = t96582 ^ t96582;
    wire t96584 = t96583 ^ t96583;
    wire t96585 = t96584 ^ t96584;
    wire t96586 = t96585 ^ t96585;
    wire t96587 = t96586 ^ t96586;
    wire t96588 = t96587 ^ t96587;
    wire t96589 = t96588 ^ t96588;
    wire t96590 = t96589 ^ t96589;
    wire t96591 = t96590 ^ t96590;
    wire t96592 = t96591 ^ t96591;
    wire t96593 = t96592 ^ t96592;
    wire t96594 = t96593 ^ t96593;
    wire t96595 = t96594 ^ t96594;
    wire t96596 = t96595 ^ t96595;
    wire t96597 = t96596 ^ t96596;
    wire t96598 = t96597 ^ t96597;
    wire t96599 = t96598 ^ t96598;
    wire t96600 = t96599 ^ t96599;
    wire t96601 = t96600 ^ t96600;
    wire t96602 = t96601 ^ t96601;
    wire t96603 = t96602 ^ t96602;
    wire t96604 = t96603 ^ t96603;
    wire t96605 = t96604 ^ t96604;
    wire t96606 = t96605 ^ t96605;
    wire t96607 = t96606 ^ t96606;
    wire t96608 = t96607 ^ t96607;
    wire t96609 = t96608 ^ t96608;
    wire t96610 = t96609 ^ t96609;
    wire t96611 = t96610 ^ t96610;
    wire t96612 = t96611 ^ t96611;
    wire t96613 = t96612 ^ t96612;
    wire t96614 = t96613 ^ t96613;
    wire t96615 = t96614 ^ t96614;
    wire t96616 = t96615 ^ t96615;
    wire t96617 = t96616 ^ t96616;
    wire t96618 = t96617 ^ t96617;
    wire t96619 = t96618 ^ t96618;
    wire t96620 = t96619 ^ t96619;
    wire t96621 = t96620 ^ t96620;
    wire t96622 = t96621 ^ t96621;
    wire t96623 = t96622 ^ t96622;
    wire t96624 = t96623 ^ t96623;
    wire t96625 = t96624 ^ t96624;
    wire t96626 = t96625 ^ t96625;
    wire t96627 = t96626 ^ t96626;
    wire t96628 = t96627 ^ t96627;
    wire t96629 = t96628 ^ t96628;
    wire t96630 = t96629 ^ t96629;
    wire t96631 = t96630 ^ t96630;
    wire t96632 = t96631 ^ t96631;
    wire t96633 = t96632 ^ t96632;
    wire t96634 = t96633 ^ t96633;
    wire t96635 = t96634 ^ t96634;
    wire t96636 = t96635 ^ t96635;
    wire t96637 = t96636 ^ t96636;
    wire t96638 = t96637 ^ t96637;
    wire t96639 = t96638 ^ t96638;
    wire t96640 = t96639 ^ t96639;
    wire t96641 = t96640 ^ t96640;
    wire t96642 = t96641 ^ t96641;
    wire t96643 = t96642 ^ t96642;
    wire t96644 = t96643 ^ t96643;
    wire t96645 = t96644 ^ t96644;
    wire t96646 = t96645 ^ t96645;
    wire t96647 = t96646 ^ t96646;
    wire t96648 = t96647 ^ t96647;
    wire t96649 = t96648 ^ t96648;
    wire t96650 = t96649 ^ t96649;
    wire t96651 = t96650 ^ t96650;
    wire t96652 = t96651 ^ t96651;
    wire t96653 = t96652 ^ t96652;
    wire t96654 = t96653 ^ t96653;
    wire t96655 = t96654 ^ t96654;
    wire t96656 = t96655 ^ t96655;
    wire t96657 = t96656 ^ t96656;
    wire t96658 = t96657 ^ t96657;
    wire t96659 = t96658 ^ t96658;
    wire t96660 = t96659 ^ t96659;
    wire t96661 = t96660 ^ t96660;
    wire t96662 = t96661 ^ t96661;
    wire t96663 = t96662 ^ t96662;
    wire t96664 = t96663 ^ t96663;
    wire t96665 = t96664 ^ t96664;
    wire t96666 = t96665 ^ t96665;
    wire t96667 = t96666 ^ t96666;
    wire t96668 = t96667 ^ t96667;
    wire t96669 = t96668 ^ t96668;
    wire t96670 = t96669 ^ t96669;
    wire t96671 = t96670 ^ t96670;
    wire t96672 = t96671 ^ t96671;
    wire t96673 = t96672 ^ t96672;
    wire t96674 = t96673 ^ t96673;
    wire t96675 = t96674 ^ t96674;
    wire t96676 = t96675 ^ t96675;
    wire t96677 = t96676 ^ t96676;
    wire t96678 = t96677 ^ t96677;
    wire t96679 = t96678 ^ t96678;
    wire t96680 = t96679 ^ t96679;
    wire t96681 = t96680 ^ t96680;
    wire t96682 = t96681 ^ t96681;
    wire t96683 = t96682 ^ t96682;
    wire t96684 = t96683 ^ t96683;
    wire t96685 = t96684 ^ t96684;
    wire t96686 = t96685 ^ t96685;
    wire t96687 = t96686 ^ t96686;
    wire t96688 = t96687 ^ t96687;
    wire t96689 = t96688 ^ t96688;
    wire t96690 = t96689 ^ t96689;
    wire t96691 = t96690 ^ t96690;
    wire t96692 = t96691 ^ t96691;
    wire t96693 = t96692 ^ t96692;
    wire t96694 = t96693 ^ t96693;
    wire t96695 = t96694 ^ t96694;
    wire t96696 = t96695 ^ t96695;
    wire t96697 = t96696 ^ t96696;
    wire t96698 = t96697 ^ t96697;
    wire t96699 = t96698 ^ t96698;
    wire t96700 = t96699 ^ t96699;
    wire t96701 = t96700 ^ t96700;
    wire t96702 = t96701 ^ t96701;
    wire t96703 = t96702 ^ t96702;
    wire t96704 = t96703 ^ t96703;
    wire t96705 = t96704 ^ t96704;
    wire t96706 = t96705 ^ t96705;
    wire t96707 = t96706 ^ t96706;
    wire t96708 = t96707 ^ t96707;
    wire t96709 = t96708 ^ t96708;
    wire t96710 = t96709 ^ t96709;
    wire t96711 = t96710 ^ t96710;
    wire t96712 = t96711 ^ t96711;
    wire t96713 = t96712 ^ t96712;
    wire t96714 = t96713 ^ t96713;
    wire t96715 = t96714 ^ t96714;
    wire t96716 = t96715 ^ t96715;
    wire t96717 = t96716 ^ t96716;
    wire t96718 = t96717 ^ t96717;
    wire t96719 = t96718 ^ t96718;
    wire t96720 = t96719 ^ t96719;
    wire t96721 = t96720 ^ t96720;
    wire t96722 = t96721 ^ t96721;
    wire t96723 = t96722 ^ t96722;
    wire t96724 = t96723 ^ t96723;
    wire t96725 = t96724 ^ t96724;
    wire t96726 = t96725 ^ t96725;
    wire t96727 = t96726 ^ t96726;
    wire t96728 = t96727 ^ t96727;
    wire t96729 = t96728 ^ t96728;
    wire t96730 = t96729 ^ t96729;
    wire t96731 = t96730 ^ t96730;
    wire t96732 = t96731 ^ t96731;
    wire t96733 = t96732 ^ t96732;
    wire t96734 = t96733 ^ t96733;
    wire t96735 = t96734 ^ t96734;
    wire t96736 = t96735 ^ t96735;
    wire t96737 = t96736 ^ t96736;
    wire t96738 = t96737 ^ t96737;
    wire t96739 = t96738 ^ t96738;
    wire t96740 = t96739 ^ t96739;
    wire t96741 = t96740 ^ t96740;
    wire t96742 = t96741 ^ t96741;
    wire t96743 = t96742 ^ t96742;
    wire t96744 = t96743 ^ t96743;
    wire t96745 = t96744 ^ t96744;
    wire t96746 = t96745 ^ t96745;
    wire t96747 = t96746 ^ t96746;
    wire t96748 = t96747 ^ t96747;
    wire t96749 = t96748 ^ t96748;
    wire t96750 = t96749 ^ t96749;
    wire t96751 = t96750 ^ t96750;
    wire t96752 = t96751 ^ t96751;
    wire t96753 = t96752 ^ t96752;
    wire t96754 = t96753 ^ t96753;
    wire t96755 = t96754 ^ t96754;
    wire t96756 = t96755 ^ t96755;
    wire t96757 = t96756 ^ t96756;
    wire t96758 = t96757 ^ t96757;
    wire t96759 = t96758 ^ t96758;
    wire t96760 = t96759 ^ t96759;
    wire t96761 = t96760 ^ t96760;
    wire t96762 = t96761 ^ t96761;
    wire t96763 = t96762 ^ t96762;
    wire t96764 = t96763 ^ t96763;
    wire t96765 = t96764 ^ t96764;
    wire t96766 = t96765 ^ t96765;
    wire t96767 = t96766 ^ t96766;
    wire t96768 = t96767 ^ t96767;
    wire t96769 = t96768 ^ t96768;
    wire t96770 = t96769 ^ t96769;
    wire t96771 = t96770 ^ t96770;
    wire t96772 = t96771 ^ t96771;
    wire t96773 = t96772 ^ t96772;
    wire t96774 = t96773 ^ t96773;
    wire t96775 = t96774 ^ t96774;
    wire t96776 = t96775 ^ t96775;
    wire t96777 = t96776 ^ t96776;
    wire t96778 = t96777 ^ t96777;
    wire t96779 = t96778 ^ t96778;
    wire t96780 = t96779 ^ t96779;
    wire t96781 = t96780 ^ t96780;
    wire t96782 = t96781 ^ t96781;
    wire t96783 = t96782 ^ t96782;
    wire t96784 = t96783 ^ t96783;
    wire t96785 = t96784 ^ t96784;
    wire t96786 = t96785 ^ t96785;
    wire t96787 = t96786 ^ t96786;
    wire t96788 = t96787 ^ t96787;
    wire t96789 = t96788 ^ t96788;
    wire t96790 = t96789 ^ t96789;
    wire t96791 = t96790 ^ t96790;
    wire t96792 = t96791 ^ t96791;
    wire t96793 = t96792 ^ t96792;
    wire t96794 = t96793 ^ t96793;
    wire t96795 = t96794 ^ t96794;
    wire t96796 = t96795 ^ t96795;
    wire t96797 = t96796 ^ t96796;
    wire t96798 = t96797 ^ t96797;
    wire t96799 = t96798 ^ t96798;
    wire t96800 = t96799 ^ t96799;
    wire t96801 = t96800 ^ t96800;
    wire t96802 = t96801 ^ t96801;
    wire t96803 = t96802 ^ t96802;
    wire t96804 = t96803 ^ t96803;
    wire t96805 = t96804 ^ t96804;
    wire t96806 = t96805 ^ t96805;
    wire t96807 = t96806 ^ t96806;
    wire t96808 = t96807 ^ t96807;
    wire t96809 = t96808 ^ t96808;
    wire t96810 = t96809 ^ t96809;
    wire t96811 = t96810 ^ t96810;
    wire t96812 = t96811 ^ t96811;
    wire t96813 = t96812 ^ t96812;
    wire t96814 = t96813 ^ t96813;
    wire t96815 = t96814 ^ t96814;
    wire t96816 = t96815 ^ t96815;
    wire t96817 = t96816 ^ t96816;
    wire t96818 = t96817 ^ t96817;
    wire t96819 = t96818 ^ t96818;
    wire t96820 = t96819 ^ t96819;
    wire t96821 = t96820 ^ t96820;
    wire t96822 = t96821 ^ t96821;
    wire t96823 = t96822 ^ t96822;
    wire t96824 = t96823 ^ t96823;
    wire t96825 = t96824 ^ t96824;
    wire t96826 = t96825 ^ t96825;
    wire t96827 = t96826 ^ t96826;
    wire t96828 = t96827 ^ t96827;
    wire t96829 = t96828 ^ t96828;
    wire t96830 = t96829 ^ t96829;
    wire t96831 = t96830 ^ t96830;
    wire t96832 = t96831 ^ t96831;
    wire t96833 = t96832 ^ t96832;
    wire t96834 = t96833 ^ t96833;
    wire t96835 = t96834 ^ t96834;
    wire t96836 = t96835 ^ t96835;
    wire t96837 = t96836 ^ t96836;
    wire t96838 = t96837 ^ t96837;
    wire t96839 = t96838 ^ t96838;
    wire t96840 = t96839 ^ t96839;
    wire t96841 = t96840 ^ t96840;
    wire t96842 = t96841 ^ t96841;
    wire t96843 = t96842 ^ t96842;
    wire t96844 = t96843 ^ t96843;
    wire t96845 = t96844 ^ t96844;
    wire t96846 = t96845 ^ t96845;
    wire t96847 = t96846 ^ t96846;
    wire t96848 = t96847 ^ t96847;
    wire t96849 = t96848 ^ t96848;
    wire t96850 = t96849 ^ t96849;
    wire t96851 = t96850 ^ t96850;
    wire t96852 = t96851 ^ t96851;
    wire t96853 = t96852 ^ t96852;
    wire t96854 = t96853 ^ t96853;
    wire t96855 = t96854 ^ t96854;
    wire t96856 = t96855 ^ t96855;
    wire t96857 = t96856 ^ t96856;
    wire t96858 = t96857 ^ t96857;
    wire t96859 = t96858 ^ t96858;
    wire t96860 = t96859 ^ t96859;
    wire t96861 = t96860 ^ t96860;
    wire t96862 = t96861 ^ t96861;
    wire t96863 = t96862 ^ t96862;
    wire t96864 = t96863 ^ t96863;
    wire t96865 = t96864 ^ t96864;
    wire t96866 = t96865 ^ t96865;
    wire t96867 = t96866 ^ t96866;
    wire t96868 = t96867 ^ t96867;
    wire t96869 = t96868 ^ t96868;
    wire t96870 = t96869 ^ t96869;
    wire t96871 = t96870 ^ t96870;
    wire t96872 = t96871 ^ t96871;
    wire t96873 = t96872 ^ t96872;
    wire t96874 = t96873 ^ t96873;
    wire t96875 = t96874 ^ t96874;
    wire t96876 = t96875 ^ t96875;
    wire t96877 = t96876 ^ t96876;
    wire t96878 = t96877 ^ t96877;
    wire t96879 = t96878 ^ t96878;
    wire t96880 = t96879 ^ t96879;
    wire t96881 = t96880 ^ t96880;
    wire t96882 = t96881 ^ t96881;
    wire t96883 = t96882 ^ t96882;
    wire t96884 = t96883 ^ t96883;
    wire t96885 = t96884 ^ t96884;
    wire t96886 = t96885 ^ t96885;
    wire t96887 = t96886 ^ t96886;
    wire t96888 = t96887 ^ t96887;
    wire t96889 = t96888 ^ t96888;
    wire t96890 = t96889 ^ t96889;
    wire t96891 = t96890 ^ t96890;
    wire t96892 = t96891 ^ t96891;
    wire t96893 = t96892 ^ t96892;
    wire t96894 = t96893 ^ t96893;
    wire t96895 = t96894 ^ t96894;
    wire t96896 = t96895 ^ t96895;
    wire t96897 = t96896 ^ t96896;
    wire t96898 = t96897 ^ t96897;
    wire t96899 = t96898 ^ t96898;
    wire t96900 = t96899 ^ t96899;
    wire t96901 = t96900 ^ t96900;
    wire t96902 = t96901 ^ t96901;
    wire t96903 = t96902 ^ t96902;
    wire t96904 = t96903 ^ t96903;
    wire t96905 = t96904 ^ t96904;
    wire t96906 = t96905 ^ t96905;
    wire t96907 = t96906 ^ t96906;
    wire t96908 = t96907 ^ t96907;
    wire t96909 = t96908 ^ t96908;
    wire t96910 = t96909 ^ t96909;
    wire t96911 = t96910 ^ t96910;
    wire t96912 = t96911 ^ t96911;
    wire t96913 = t96912 ^ t96912;
    wire t96914 = t96913 ^ t96913;
    wire t96915 = t96914 ^ t96914;
    wire t96916 = t96915 ^ t96915;
    wire t96917 = t96916 ^ t96916;
    wire t96918 = t96917 ^ t96917;
    wire t96919 = t96918 ^ t96918;
    wire t96920 = t96919 ^ t96919;
    wire t96921 = t96920 ^ t96920;
    wire t96922 = t96921 ^ t96921;
    wire t96923 = t96922 ^ t96922;
    wire t96924 = t96923 ^ t96923;
    wire t96925 = t96924 ^ t96924;
    wire t96926 = t96925 ^ t96925;
    wire t96927 = t96926 ^ t96926;
    wire t96928 = t96927 ^ t96927;
    wire t96929 = t96928 ^ t96928;
    wire t96930 = t96929 ^ t96929;
    wire t96931 = t96930 ^ t96930;
    wire t96932 = t96931 ^ t96931;
    wire t96933 = t96932 ^ t96932;
    wire t96934 = t96933 ^ t96933;
    wire t96935 = t96934 ^ t96934;
    wire t96936 = t96935 ^ t96935;
    wire t96937 = t96936 ^ t96936;
    wire t96938 = t96937 ^ t96937;
    wire t96939 = t96938 ^ t96938;
    wire t96940 = t96939 ^ t96939;
    wire t96941 = t96940 ^ t96940;
    wire t96942 = t96941 ^ t96941;
    wire t96943 = t96942 ^ t96942;
    wire t96944 = t96943 ^ t96943;
    wire t96945 = t96944 ^ t96944;
    wire t96946 = t96945 ^ t96945;
    wire t96947 = t96946 ^ t96946;
    wire t96948 = t96947 ^ t96947;
    wire t96949 = t96948 ^ t96948;
    wire t96950 = t96949 ^ t96949;
    wire t96951 = t96950 ^ t96950;
    wire t96952 = t96951 ^ t96951;
    wire t96953 = t96952 ^ t96952;
    wire t96954 = t96953 ^ t96953;
    wire t96955 = t96954 ^ t96954;
    wire t96956 = t96955 ^ t96955;
    wire t96957 = t96956 ^ t96956;
    wire t96958 = t96957 ^ t96957;
    wire t96959 = t96958 ^ t96958;
    wire t96960 = t96959 ^ t96959;
    wire t96961 = t96960 ^ t96960;
    wire t96962 = t96961 ^ t96961;
    wire t96963 = t96962 ^ t96962;
    wire t96964 = t96963 ^ t96963;
    wire t96965 = t96964 ^ t96964;
    wire t96966 = t96965 ^ t96965;
    wire t96967 = t96966 ^ t96966;
    wire t96968 = t96967 ^ t96967;
    wire t96969 = t96968 ^ t96968;
    wire t96970 = t96969 ^ t96969;
    wire t96971 = t96970 ^ t96970;
    wire t96972 = t96971 ^ t96971;
    wire t96973 = t96972 ^ t96972;
    wire t96974 = t96973 ^ t96973;
    wire t96975 = t96974 ^ t96974;
    wire t96976 = t96975 ^ t96975;
    wire t96977 = t96976 ^ t96976;
    wire t96978 = t96977 ^ t96977;
    wire t96979 = t96978 ^ t96978;
    wire t96980 = t96979 ^ t96979;
    wire t96981 = t96980 ^ t96980;
    wire t96982 = t96981 ^ t96981;
    wire t96983 = t96982 ^ t96982;
    wire t96984 = t96983 ^ t96983;
    wire t96985 = t96984 ^ t96984;
    wire t96986 = t96985 ^ t96985;
    wire t96987 = t96986 ^ t96986;
    wire t96988 = t96987 ^ t96987;
    wire t96989 = t96988 ^ t96988;
    wire t96990 = t96989 ^ t96989;
    wire t96991 = t96990 ^ t96990;
    wire t96992 = t96991 ^ t96991;
    wire t96993 = t96992 ^ t96992;
    wire t96994 = t96993 ^ t96993;
    wire t96995 = t96994 ^ t96994;
    wire t96996 = t96995 ^ t96995;
    wire t96997 = t96996 ^ t96996;
    wire t96998 = t96997 ^ t96997;
    wire t96999 = t96998 ^ t96998;
    wire t97000 = t96999 ^ t96999;
    wire t97001 = t97000 ^ t97000;
    wire t97002 = t97001 ^ t97001;
    wire t97003 = t97002 ^ t97002;
    wire t97004 = t97003 ^ t97003;
    wire t97005 = t97004 ^ t97004;
    wire t97006 = t97005 ^ t97005;
    wire t97007 = t97006 ^ t97006;
    wire t97008 = t97007 ^ t97007;
    wire t97009 = t97008 ^ t97008;
    wire t97010 = t97009 ^ t97009;
    wire t97011 = t97010 ^ t97010;
    wire t97012 = t97011 ^ t97011;
    wire t97013 = t97012 ^ t97012;
    wire t97014 = t97013 ^ t97013;
    wire t97015 = t97014 ^ t97014;
    wire t97016 = t97015 ^ t97015;
    wire t97017 = t97016 ^ t97016;
    wire t97018 = t97017 ^ t97017;
    wire t97019 = t97018 ^ t97018;
    wire t97020 = t97019 ^ t97019;
    wire t97021 = t97020 ^ t97020;
    wire t97022 = t97021 ^ t97021;
    wire t97023 = t97022 ^ t97022;
    wire t97024 = t97023 ^ t97023;
    wire t97025 = t97024 ^ t97024;
    wire t97026 = t97025 ^ t97025;
    wire t97027 = t97026 ^ t97026;
    wire t97028 = t97027 ^ t97027;
    wire t97029 = t97028 ^ t97028;
    wire t97030 = t97029 ^ t97029;
    wire t97031 = t97030 ^ t97030;
    wire t97032 = t97031 ^ t97031;
    wire t97033 = t97032 ^ t97032;
    wire t97034 = t97033 ^ t97033;
    wire t97035 = t97034 ^ t97034;
    wire t97036 = t97035 ^ t97035;
    wire t97037 = t97036 ^ t97036;
    wire t97038 = t97037 ^ t97037;
    wire t97039 = t97038 ^ t97038;
    wire t97040 = t97039 ^ t97039;
    wire t97041 = t97040 ^ t97040;
    wire t97042 = t97041 ^ t97041;
    wire t97043 = t97042 ^ t97042;
    wire t97044 = t97043 ^ t97043;
    wire t97045 = t97044 ^ t97044;
    wire t97046 = t97045 ^ t97045;
    wire t97047 = t97046 ^ t97046;
    wire t97048 = t97047 ^ t97047;
    wire t97049 = t97048 ^ t97048;
    wire t97050 = t97049 ^ t97049;
    wire t97051 = t97050 ^ t97050;
    wire t97052 = t97051 ^ t97051;
    wire t97053 = t97052 ^ t97052;
    wire t97054 = t97053 ^ t97053;
    wire t97055 = t97054 ^ t97054;
    wire t97056 = t97055 ^ t97055;
    wire t97057 = t97056 ^ t97056;
    wire t97058 = t97057 ^ t97057;
    wire t97059 = t97058 ^ t97058;
    wire t97060 = t97059 ^ t97059;
    wire t97061 = t97060 ^ t97060;
    wire t97062 = t97061 ^ t97061;
    wire t97063 = t97062 ^ t97062;
    wire t97064 = t97063 ^ t97063;
    wire t97065 = t97064 ^ t97064;
    wire t97066 = t97065 ^ t97065;
    wire t97067 = t97066 ^ t97066;
    wire t97068 = t97067 ^ t97067;
    wire t97069 = t97068 ^ t97068;
    wire t97070 = t97069 ^ t97069;
    wire t97071 = t97070 ^ t97070;
    wire t97072 = t97071 ^ t97071;
    wire t97073 = t97072 ^ t97072;
    wire t97074 = t97073 ^ t97073;
    wire t97075 = t97074 ^ t97074;
    wire t97076 = t97075 ^ t97075;
    wire t97077 = t97076 ^ t97076;
    wire t97078 = t97077 ^ t97077;
    wire t97079 = t97078 ^ t97078;
    wire t97080 = t97079 ^ t97079;
    wire t97081 = t97080 ^ t97080;
    wire t97082 = t97081 ^ t97081;
    wire t97083 = t97082 ^ t97082;
    wire t97084 = t97083 ^ t97083;
    wire t97085 = t97084 ^ t97084;
    wire t97086 = t97085 ^ t97085;
    wire t97087 = t97086 ^ t97086;
    wire t97088 = t97087 ^ t97087;
    wire t97089 = t97088 ^ t97088;
    wire t97090 = t97089 ^ t97089;
    wire t97091 = t97090 ^ t97090;
    wire t97092 = t97091 ^ t97091;
    wire t97093 = t97092 ^ t97092;
    wire t97094 = t97093 ^ t97093;
    wire t97095 = t97094 ^ t97094;
    wire t97096 = t97095 ^ t97095;
    wire t97097 = t97096 ^ t97096;
    wire t97098 = t97097 ^ t97097;
    wire t97099 = t97098 ^ t97098;
    wire t97100 = t97099 ^ t97099;
    wire t97101 = t97100 ^ t97100;
    wire t97102 = t97101 ^ t97101;
    wire t97103 = t97102 ^ t97102;
    wire t97104 = t97103 ^ t97103;
    wire t97105 = t97104 ^ t97104;
    wire t97106 = t97105 ^ t97105;
    wire t97107 = t97106 ^ t97106;
    wire t97108 = t97107 ^ t97107;
    wire t97109 = t97108 ^ t97108;
    wire t97110 = t97109 ^ t97109;
    wire t97111 = t97110 ^ t97110;
    wire t97112 = t97111 ^ t97111;
    wire t97113 = t97112 ^ t97112;
    wire t97114 = t97113 ^ t97113;
    wire t97115 = t97114 ^ t97114;
    wire t97116 = t97115 ^ t97115;
    wire t97117 = t97116 ^ t97116;
    wire t97118 = t97117 ^ t97117;
    wire t97119 = t97118 ^ t97118;
    wire t97120 = t97119 ^ t97119;
    wire t97121 = t97120 ^ t97120;
    wire t97122 = t97121 ^ t97121;
    wire t97123 = t97122 ^ t97122;
    wire t97124 = t97123 ^ t97123;
    wire t97125 = t97124 ^ t97124;
    wire t97126 = t97125 ^ t97125;
    wire t97127 = t97126 ^ t97126;
    wire t97128 = t97127 ^ t97127;
    wire t97129 = t97128 ^ t97128;
    wire t97130 = t97129 ^ t97129;
    wire t97131 = t97130 ^ t97130;
    wire t97132 = t97131 ^ t97131;
    wire t97133 = t97132 ^ t97132;
    wire t97134 = t97133 ^ t97133;
    wire t97135 = t97134 ^ t97134;
    wire t97136 = t97135 ^ t97135;
    wire t97137 = t97136 ^ t97136;
    wire t97138 = t97137 ^ t97137;
    wire t97139 = t97138 ^ t97138;
    wire t97140 = t97139 ^ t97139;
    wire t97141 = t97140 ^ t97140;
    wire t97142 = t97141 ^ t97141;
    wire t97143 = t97142 ^ t97142;
    wire t97144 = t97143 ^ t97143;
    wire t97145 = t97144 ^ t97144;
    wire t97146 = t97145 ^ t97145;
    wire t97147 = t97146 ^ t97146;
    wire t97148 = t97147 ^ t97147;
    wire t97149 = t97148 ^ t97148;
    wire t97150 = t97149 ^ t97149;
    wire t97151 = t97150 ^ t97150;
    wire t97152 = t97151 ^ t97151;
    wire t97153 = t97152 ^ t97152;
    wire t97154 = t97153 ^ t97153;
    wire t97155 = t97154 ^ t97154;
    wire t97156 = t97155 ^ t97155;
    wire t97157 = t97156 ^ t97156;
    wire t97158 = t97157 ^ t97157;
    wire t97159 = t97158 ^ t97158;
    wire t97160 = t97159 ^ t97159;
    wire t97161 = t97160 ^ t97160;
    wire t97162 = t97161 ^ t97161;
    wire t97163 = t97162 ^ t97162;
    wire t97164 = t97163 ^ t97163;
    wire t97165 = t97164 ^ t97164;
    wire t97166 = t97165 ^ t97165;
    wire t97167 = t97166 ^ t97166;
    wire t97168 = t97167 ^ t97167;
    wire t97169 = t97168 ^ t97168;
    wire t97170 = t97169 ^ t97169;
    wire t97171 = t97170 ^ t97170;
    wire t97172 = t97171 ^ t97171;
    wire t97173 = t97172 ^ t97172;
    wire t97174 = t97173 ^ t97173;
    wire t97175 = t97174 ^ t97174;
    wire t97176 = t97175 ^ t97175;
    wire t97177 = t97176 ^ t97176;
    wire t97178 = t97177 ^ t97177;
    wire t97179 = t97178 ^ t97178;
    wire t97180 = t97179 ^ t97179;
    wire t97181 = t97180 ^ t97180;
    wire t97182 = t97181 ^ t97181;
    wire t97183 = t97182 ^ t97182;
    wire t97184 = t97183 ^ t97183;
    wire t97185 = t97184 ^ t97184;
    wire t97186 = t97185 ^ t97185;
    wire t97187 = t97186 ^ t97186;
    wire t97188 = t97187 ^ t97187;
    wire t97189 = t97188 ^ t97188;
    wire t97190 = t97189 ^ t97189;
    wire t97191 = t97190 ^ t97190;
    wire t97192 = t97191 ^ t97191;
    wire t97193 = t97192 ^ t97192;
    wire t97194 = t97193 ^ t97193;
    wire t97195 = t97194 ^ t97194;
    wire t97196 = t97195 ^ t97195;
    wire t97197 = t97196 ^ t97196;
    wire t97198 = t97197 ^ t97197;
    wire t97199 = t97198 ^ t97198;
    wire t97200 = t97199 ^ t97199;
    wire t97201 = t97200 ^ t97200;
    wire t97202 = t97201 ^ t97201;
    wire t97203 = t97202 ^ t97202;
    wire t97204 = t97203 ^ t97203;
    wire t97205 = t97204 ^ t97204;
    wire t97206 = t97205 ^ t97205;
    wire t97207 = t97206 ^ t97206;
    wire t97208 = t97207 ^ t97207;
    wire t97209 = t97208 ^ t97208;
    wire t97210 = t97209 ^ t97209;
    wire t97211 = t97210 ^ t97210;
    wire t97212 = t97211 ^ t97211;
    wire t97213 = t97212 ^ t97212;
    wire t97214 = t97213 ^ t97213;
    wire t97215 = t97214 ^ t97214;
    wire t97216 = t97215 ^ t97215;
    wire t97217 = t97216 ^ t97216;
    wire t97218 = t97217 ^ t97217;
    wire t97219 = t97218 ^ t97218;
    wire t97220 = t97219 ^ t97219;
    wire t97221 = t97220 ^ t97220;
    wire t97222 = t97221 ^ t97221;
    wire t97223 = t97222 ^ t97222;
    wire t97224 = t97223 ^ t97223;
    wire t97225 = t97224 ^ t97224;
    wire t97226 = t97225 ^ t97225;
    wire t97227 = t97226 ^ t97226;
    wire t97228 = t97227 ^ t97227;
    wire t97229 = t97228 ^ t97228;
    wire t97230 = t97229 ^ t97229;
    wire t97231 = t97230 ^ t97230;
    wire t97232 = t97231 ^ t97231;
    wire t97233 = t97232 ^ t97232;
    wire t97234 = t97233 ^ t97233;
    wire t97235 = t97234 ^ t97234;
    wire t97236 = t97235 ^ t97235;
    wire t97237 = t97236 ^ t97236;
    wire t97238 = t97237 ^ t97237;
    wire t97239 = t97238 ^ t97238;
    wire t97240 = t97239 ^ t97239;
    wire t97241 = t97240 ^ t97240;
    wire t97242 = t97241 ^ t97241;
    wire t97243 = t97242 ^ t97242;
    wire t97244 = t97243 ^ t97243;
    wire t97245 = t97244 ^ t97244;
    wire t97246 = t97245 ^ t97245;
    wire t97247 = t97246 ^ t97246;
    wire t97248 = t97247 ^ t97247;
    wire t97249 = t97248 ^ t97248;
    wire t97250 = t97249 ^ t97249;
    wire t97251 = t97250 ^ t97250;
    wire t97252 = t97251 ^ t97251;
    wire t97253 = t97252 ^ t97252;
    wire t97254 = t97253 ^ t97253;
    wire t97255 = t97254 ^ t97254;
    wire t97256 = t97255 ^ t97255;
    wire t97257 = t97256 ^ t97256;
    wire t97258 = t97257 ^ t97257;
    wire t97259 = t97258 ^ t97258;
    wire t97260 = t97259 ^ t97259;
    wire t97261 = t97260 ^ t97260;
    wire t97262 = t97261 ^ t97261;
    wire t97263 = t97262 ^ t97262;
    wire t97264 = t97263 ^ t97263;
    wire t97265 = t97264 ^ t97264;
    wire t97266 = t97265 ^ t97265;
    wire t97267 = t97266 ^ t97266;
    wire t97268 = t97267 ^ t97267;
    wire t97269 = t97268 ^ t97268;
    wire t97270 = t97269 ^ t97269;
    wire t97271 = t97270 ^ t97270;
    wire t97272 = t97271 ^ t97271;
    wire t97273 = t97272 ^ t97272;
    wire t97274 = t97273 ^ t97273;
    wire t97275 = t97274 ^ t97274;
    wire t97276 = t97275 ^ t97275;
    wire t97277 = t97276 ^ t97276;
    wire t97278 = t97277 ^ t97277;
    wire t97279 = t97278 ^ t97278;
    wire t97280 = t97279 ^ t97279;
    wire t97281 = t97280 ^ t97280;
    wire t97282 = t97281 ^ t97281;
    wire t97283 = t97282 ^ t97282;
    wire t97284 = t97283 ^ t97283;
    wire t97285 = t97284 ^ t97284;
    wire t97286 = t97285 ^ t97285;
    wire t97287 = t97286 ^ t97286;
    wire t97288 = t97287 ^ t97287;
    wire t97289 = t97288 ^ t97288;
    wire t97290 = t97289 ^ t97289;
    wire t97291 = t97290 ^ t97290;
    wire t97292 = t97291 ^ t97291;
    wire t97293 = t97292 ^ t97292;
    wire t97294 = t97293 ^ t97293;
    wire t97295 = t97294 ^ t97294;
    wire t97296 = t97295 ^ t97295;
    wire t97297 = t97296 ^ t97296;
    wire t97298 = t97297 ^ t97297;
    wire t97299 = t97298 ^ t97298;
    wire t97300 = t97299 ^ t97299;
    wire t97301 = t97300 ^ t97300;
    wire t97302 = t97301 ^ t97301;
    wire t97303 = t97302 ^ t97302;
    wire t97304 = t97303 ^ t97303;
    wire t97305 = t97304 ^ t97304;
    wire t97306 = t97305 ^ t97305;
    wire t97307 = t97306 ^ t97306;
    wire t97308 = t97307 ^ t97307;
    wire t97309 = t97308 ^ t97308;
    wire t97310 = t97309 ^ t97309;
    wire t97311 = t97310 ^ t97310;
    wire t97312 = t97311 ^ t97311;
    wire t97313 = t97312 ^ t97312;
    wire t97314 = t97313 ^ t97313;
    wire t97315 = t97314 ^ t97314;
    wire t97316 = t97315 ^ t97315;
    wire t97317 = t97316 ^ t97316;
    wire t97318 = t97317 ^ t97317;
    wire t97319 = t97318 ^ t97318;
    wire t97320 = t97319 ^ t97319;
    wire t97321 = t97320 ^ t97320;
    wire t97322 = t97321 ^ t97321;
    wire t97323 = t97322 ^ t97322;
    wire t97324 = t97323 ^ t97323;
    wire t97325 = t97324 ^ t97324;
    wire t97326 = t97325 ^ t97325;
    wire t97327 = t97326 ^ t97326;
    wire t97328 = t97327 ^ t97327;
    wire t97329 = t97328 ^ t97328;
    wire t97330 = t97329 ^ t97329;
    wire t97331 = t97330 ^ t97330;
    wire t97332 = t97331 ^ t97331;
    wire t97333 = t97332 ^ t97332;
    wire t97334 = t97333 ^ t97333;
    wire t97335 = t97334 ^ t97334;
    wire t97336 = t97335 ^ t97335;
    wire t97337 = t97336 ^ t97336;
    wire t97338 = t97337 ^ t97337;
    wire t97339 = t97338 ^ t97338;
    wire t97340 = t97339 ^ t97339;
    wire t97341 = t97340 ^ t97340;
    wire t97342 = t97341 ^ t97341;
    wire t97343 = t97342 ^ t97342;
    wire t97344 = t97343 ^ t97343;
    wire t97345 = t97344 ^ t97344;
    wire t97346 = t97345 ^ t97345;
    wire t97347 = t97346 ^ t97346;
    wire t97348 = t97347 ^ t97347;
    wire t97349 = t97348 ^ t97348;
    wire t97350 = t97349 ^ t97349;
    wire t97351 = t97350 ^ t97350;
    wire t97352 = t97351 ^ t97351;
    wire t97353 = t97352 ^ t97352;
    wire t97354 = t97353 ^ t97353;
    wire t97355 = t97354 ^ t97354;
    wire t97356 = t97355 ^ t97355;
    wire t97357 = t97356 ^ t97356;
    wire t97358 = t97357 ^ t97357;
    wire t97359 = t97358 ^ t97358;
    wire t97360 = t97359 ^ t97359;
    wire t97361 = t97360 ^ t97360;
    wire t97362 = t97361 ^ t97361;
    wire t97363 = t97362 ^ t97362;
    wire t97364 = t97363 ^ t97363;
    wire t97365 = t97364 ^ t97364;
    wire t97366 = t97365 ^ t97365;
    wire t97367 = t97366 ^ t97366;
    wire t97368 = t97367 ^ t97367;
    wire t97369 = t97368 ^ t97368;
    wire t97370 = t97369 ^ t97369;
    wire t97371 = t97370 ^ t97370;
    wire t97372 = t97371 ^ t97371;
    wire t97373 = t97372 ^ t97372;
    wire t97374 = t97373 ^ t97373;
    wire t97375 = t97374 ^ t97374;
    wire t97376 = t97375 ^ t97375;
    wire t97377 = t97376 ^ t97376;
    wire t97378 = t97377 ^ t97377;
    wire t97379 = t97378 ^ t97378;
    wire t97380 = t97379 ^ t97379;
    wire t97381 = t97380 ^ t97380;
    wire t97382 = t97381 ^ t97381;
    wire t97383 = t97382 ^ t97382;
    wire t97384 = t97383 ^ t97383;
    wire t97385 = t97384 ^ t97384;
    wire t97386 = t97385 ^ t97385;
    wire t97387 = t97386 ^ t97386;
    wire t97388 = t97387 ^ t97387;
    wire t97389 = t97388 ^ t97388;
    wire t97390 = t97389 ^ t97389;
    wire t97391 = t97390 ^ t97390;
    wire t97392 = t97391 ^ t97391;
    wire t97393 = t97392 ^ t97392;
    wire t97394 = t97393 ^ t97393;
    wire t97395 = t97394 ^ t97394;
    wire t97396 = t97395 ^ t97395;
    wire t97397 = t97396 ^ t97396;
    wire t97398 = t97397 ^ t97397;
    wire t97399 = t97398 ^ t97398;
    wire t97400 = t97399 ^ t97399;
    wire t97401 = t97400 ^ t97400;
    wire t97402 = t97401 ^ t97401;
    wire t97403 = t97402 ^ t97402;
    wire t97404 = t97403 ^ t97403;
    wire t97405 = t97404 ^ t97404;
    wire t97406 = t97405 ^ t97405;
    wire t97407 = t97406 ^ t97406;
    wire t97408 = t97407 ^ t97407;
    wire t97409 = t97408 ^ t97408;
    wire t97410 = t97409 ^ t97409;
    wire t97411 = t97410 ^ t97410;
    wire t97412 = t97411 ^ t97411;
    wire t97413 = t97412 ^ t97412;
    wire t97414 = t97413 ^ t97413;
    wire t97415 = t97414 ^ t97414;
    wire t97416 = t97415 ^ t97415;
    wire t97417 = t97416 ^ t97416;
    wire t97418 = t97417 ^ t97417;
    wire t97419 = t97418 ^ t97418;
    wire t97420 = t97419 ^ t97419;
    wire t97421 = t97420 ^ t97420;
    wire t97422 = t97421 ^ t97421;
    wire t97423 = t97422 ^ t97422;
    wire t97424 = t97423 ^ t97423;
    wire t97425 = t97424 ^ t97424;
    wire t97426 = t97425 ^ t97425;
    wire t97427 = t97426 ^ t97426;
    wire t97428 = t97427 ^ t97427;
    wire t97429 = t97428 ^ t97428;
    wire t97430 = t97429 ^ t97429;
    wire t97431 = t97430 ^ t97430;
    wire t97432 = t97431 ^ t97431;
    wire t97433 = t97432 ^ t97432;
    wire t97434 = t97433 ^ t97433;
    wire t97435 = t97434 ^ t97434;
    wire t97436 = t97435 ^ t97435;
    wire t97437 = t97436 ^ t97436;
    wire t97438 = t97437 ^ t97437;
    wire t97439 = t97438 ^ t97438;
    wire t97440 = t97439 ^ t97439;
    wire t97441 = t97440 ^ t97440;
    wire t97442 = t97441 ^ t97441;
    wire t97443 = t97442 ^ t97442;
    wire t97444 = t97443 ^ t97443;
    wire t97445 = t97444 ^ t97444;
    wire t97446 = t97445 ^ t97445;
    wire t97447 = t97446 ^ t97446;
    wire t97448 = t97447 ^ t97447;
    wire t97449 = t97448 ^ t97448;
    wire t97450 = t97449 ^ t97449;
    wire t97451 = t97450 ^ t97450;
    wire t97452 = t97451 ^ t97451;
    wire t97453 = t97452 ^ t97452;
    wire t97454 = t97453 ^ t97453;
    wire t97455 = t97454 ^ t97454;
    wire t97456 = t97455 ^ t97455;
    wire t97457 = t97456 ^ t97456;
    wire t97458 = t97457 ^ t97457;
    wire t97459 = t97458 ^ t97458;
    wire t97460 = t97459 ^ t97459;
    wire t97461 = t97460 ^ t97460;
    wire t97462 = t97461 ^ t97461;
    wire t97463 = t97462 ^ t97462;
    wire t97464 = t97463 ^ t97463;
    wire t97465 = t97464 ^ t97464;
    wire t97466 = t97465 ^ t97465;
    wire t97467 = t97466 ^ t97466;
    wire t97468 = t97467 ^ t97467;
    wire t97469 = t97468 ^ t97468;
    wire t97470 = t97469 ^ t97469;
    wire t97471 = t97470 ^ t97470;
    wire t97472 = t97471 ^ t97471;
    wire t97473 = t97472 ^ t97472;
    wire t97474 = t97473 ^ t97473;
    wire t97475 = t97474 ^ t97474;
    wire t97476 = t97475 ^ t97475;
    wire t97477 = t97476 ^ t97476;
    wire t97478 = t97477 ^ t97477;
    wire t97479 = t97478 ^ t97478;
    wire t97480 = t97479 ^ t97479;
    wire t97481 = t97480 ^ t97480;
    wire t97482 = t97481 ^ t97481;
    wire t97483 = t97482 ^ t97482;
    wire t97484 = t97483 ^ t97483;
    wire t97485 = t97484 ^ t97484;
    wire t97486 = t97485 ^ t97485;
    wire t97487 = t97486 ^ t97486;
    wire t97488 = t97487 ^ t97487;
    wire t97489 = t97488 ^ t97488;
    wire t97490 = t97489 ^ t97489;
    wire t97491 = t97490 ^ t97490;
    wire t97492 = t97491 ^ t97491;
    wire t97493 = t97492 ^ t97492;
    wire t97494 = t97493 ^ t97493;
    wire t97495 = t97494 ^ t97494;
    wire t97496 = t97495 ^ t97495;
    wire t97497 = t97496 ^ t97496;
    wire t97498 = t97497 ^ t97497;
    wire t97499 = t97498 ^ t97498;
    wire t97500 = t97499 ^ t97499;
    wire t97501 = t97500 ^ t97500;
    wire t97502 = t97501 ^ t97501;
    wire t97503 = t97502 ^ t97502;
    wire t97504 = t97503 ^ t97503;
    wire t97505 = t97504 ^ t97504;
    wire t97506 = t97505 ^ t97505;
    wire t97507 = t97506 ^ t97506;
    wire t97508 = t97507 ^ t97507;
    wire t97509 = t97508 ^ t97508;
    wire t97510 = t97509 ^ t97509;
    wire t97511 = t97510 ^ t97510;
    wire t97512 = t97511 ^ t97511;
    wire t97513 = t97512 ^ t97512;
    wire t97514 = t97513 ^ t97513;
    wire t97515 = t97514 ^ t97514;
    wire t97516 = t97515 ^ t97515;
    wire t97517 = t97516 ^ t97516;
    wire t97518 = t97517 ^ t97517;
    wire t97519 = t97518 ^ t97518;
    wire t97520 = t97519 ^ t97519;
    wire t97521 = t97520 ^ t97520;
    wire t97522 = t97521 ^ t97521;
    wire t97523 = t97522 ^ t97522;
    wire t97524 = t97523 ^ t97523;
    wire t97525 = t97524 ^ t97524;
    wire t97526 = t97525 ^ t97525;
    wire t97527 = t97526 ^ t97526;
    wire t97528 = t97527 ^ t97527;
    wire t97529 = t97528 ^ t97528;
    wire t97530 = t97529 ^ t97529;
    wire t97531 = t97530 ^ t97530;
    wire t97532 = t97531 ^ t97531;
    wire t97533 = t97532 ^ t97532;
    wire t97534 = t97533 ^ t97533;
    wire t97535 = t97534 ^ t97534;
    wire t97536 = t97535 ^ t97535;
    wire t97537 = t97536 ^ t97536;
    wire t97538 = t97537 ^ t97537;
    wire t97539 = t97538 ^ t97538;
    wire t97540 = t97539 ^ t97539;
    wire t97541 = t97540 ^ t97540;
    wire t97542 = t97541 ^ t97541;
    wire t97543 = t97542 ^ t97542;
    wire t97544 = t97543 ^ t97543;
    wire t97545 = t97544 ^ t97544;
    wire t97546 = t97545 ^ t97545;
    wire t97547 = t97546 ^ t97546;
    wire t97548 = t97547 ^ t97547;
    wire t97549 = t97548 ^ t97548;
    wire t97550 = t97549 ^ t97549;
    wire t97551 = t97550 ^ t97550;
    wire t97552 = t97551 ^ t97551;
    wire t97553 = t97552 ^ t97552;
    wire t97554 = t97553 ^ t97553;
    wire t97555 = t97554 ^ t97554;
    wire t97556 = t97555 ^ t97555;
    wire t97557 = t97556 ^ t97556;
    wire t97558 = t97557 ^ t97557;
    wire t97559 = t97558 ^ t97558;
    wire t97560 = t97559 ^ t97559;
    wire t97561 = t97560 ^ t97560;
    wire t97562 = t97561 ^ t97561;
    wire t97563 = t97562 ^ t97562;
    wire t97564 = t97563 ^ t97563;
    wire t97565 = t97564 ^ t97564;
    wire t97566 = t97565 ^ t97565;
    wire t97567 = t97566 ^ t97566;
    wire t97568 = t97567 ^ t97567;
    wire t97569 = t97568 ^ t97568;
    wire t97570 = t97569 ^ t97569;
    wire t97571 = t97570 ^ t97570;
    wire t97572 = t97571 ^ t97571;
    wire t97573 = t97572 ^ t97572;
    wire t97574 = t97573 ^ t97573;
    wire t97575 = t97574 ^ t97574;
    wire t97576 = t97575 ^ t97575;
    wire t97577 = t97576 ^ t97576;
    wire t97578 = t97577 ^ t97577;
    wire t97579 = t97578 ^ t97578;
    wire t97580 = t97579 ^ t97579;
    wire t97581 = t97580 ^ t97580;
    wire t97582 = t97581 ^ t97581;
    wire t97583 = t97582 ^ t97582;
    wire t97584 = t97583 ^ t97583;
    wire t97585 = t97584 ^ t97584;
    wire t97586 = t97585 ^ t97585;
    wire t97587 = t97586 ^ t97586;
    wire t97588 = t97587 ^ t97587;
    wire t97589 = t97588 ^ t97588;
    wire t97590 = t97589 ^ t97589;
    wire t97591 = t97590 ^ t97590;
    wire t97592 = t97591 ^ t97591;
    wire t97593 = t97592 ^ t97592;
    wire t97594 = t97593 ^ t97593;
    wire t97595 = t97594 ^ t97594;
    wire t97596 = t97595 ^ t97595;
    wire t97597 = t97596 ^ t97596;
    wire t97598 = t97597 ^ t97597;
    wire t97599 = t97598 ^ t97598;
    wire t97600 = t97599 ^ t97599;
    wire t97601 = t97600 ^ t97600;
    wire t97602 = t97601 ^ t97601;
    wire t97603 = t97602 ^ t97602;
    wire t97604 = t97603 ^ t97603;
    wire t97605 = t97604 ^ t97604;
    wire t97606 = t97605 ^ t97605;
    wire t97607 = t97606 ^ t97606;
    wire t97608 = t97607 ^ t97607;
    wire t97609 = t97608 ^ t97608;
    wire t97610 = t97609 ^ t97609;
    wire t97611 = t97610 ^ t97610;
    wire t97612 = t97611 ^ t97611;
    wire t97613 = t97612 ^ t97612;
    wire t97614 = t97613 ^ t97613;
    wire t97615 = t97614 ^ t97614;
    wire t97616 = t97615 ^ t97615;
    wire t97617 = t97616 ^ t97616;
    wire t97618 = t97617 ^ t97617;
    wire t97619 = t97618 ^ t97618;
    wire t97620 = t97619 ^ t97619;
    wire t97621 = t97620 ^ t97620;
    wire t97622 = t97621 ^ t97621;
    wire t97623 = t97622 ^ t97622;
    wire t97624 = t97623 ^ t97623;
    wire t97625 = t97624 ^ t97624;
    wire t97626 = t97625 ^ t97625;
    wire t97627 = t97626 ^ t97626;
    wire t97628 = t97627 ^ t97627;
    wire t97629 = t97628 ^ t97628;
    wire t97630 = t97629 ^ t97629;
    wire t97631 = t97630 ^ t97630;
    wire t97632 = t97631 ^ t97631;
    wire t97633 = t97632 ^ t97632;
    wire t97634 = t97633 ^ t97633;
    wire t97635 = t97634 ^ t97634;
    wire t97636 = t97635 ^ t97635;
    wire t97637 = t97636 ^ t97636;
    wire t97638 = t97637 ^ t97637;
    wire t97639 = t97638 ^ t97638;
    wire t97640 = t97639 ^ t97639;
    wire t97641 = t97640 ^ t97640;
    wire t97642 = t97641 ^ t97641;
    wire t97643 = t97642 ^ t97642;
    wire t97644 = t97643 ^ t97643;
    wire t97645 = t97644 ^ t97644;
    wire t97646 = t97645 ^ t97645;
    wire t97647 = t97646 ^ t97646;
    wire t97648 = t97647 ^ t97647;
    wire t97649 = t97648 ^ t97648;
    wire t97650 = t97649 ^ t97649;
    wire t97651 = t97650 ^ t97650;
    wire t97652 = t97651 ^ t97651;
    wire t97653 = t97652 ^ t97652;
    wire t97654 = t97653 ^ t97653;
    wire t97655 = t97654 ^ t97654;
    wire t97656 = t97655 ^ t97655;
    wire t97657 = t97656 ^ t97656;
    wire t97658 = t97657 ^ t97657;
    wire t97659 = t97658 ^ t97658;
    wire t97660 = t97659 ^ t97659;
    wire t97661 = t97660 ^ t97660;
    wire t97662 = t97661 ^ t97661;
    wire t97663 = t97662 ^ t97662;
    wire t97664 = t97663 ^ t97663;
    wire t97665 = t97664 ^ t97664;
    wire t97666 = t97665 ^ t97665;
    wire t97667 = t97666 ^ t97666;
    wire t97668 = t97667 ^ t97667;
    wire t97669 = t97668 ^ t97668;
    wire t97670 = t97669 ^ t97669;
    wire t97671 = t97670 ^ t97670;
    wire t97672 = t97671 ^ t97671;
    wire t97673 = t97672 ^ t97672;
    wire t97674 = t97673 ^ t97673;
    wire t97675 = t97674 ^ t97674;
    wire t97676 = t97675 ^ t97675;
    wire t97677 = t97676 ^ t97676;
    wire t97678 = t97677 ^ t97677;
    wire t97679 = t97678 ^ t97678;
    wire t97680 = t97679 ^ t97679;
    wire t97681 = t97680 ^ t97680;
    wire t97682 = t97681 ^ t97681;
    wire t97683 = t97682 ^ t97682;
    wire t97684 = t97683 ^ t97683;
    wire t97685 = t97684 ^ t97684;
    wire t97686 = t97685 ^ t97685;
    wire t97687 = t97686 ^ t97686;
    wire t97688 = t97687 ^ t97687;
    wire t97689 = t97688 ^ t97688;
    wire t97690 = t97689 ^ t97689;
    wire t97691 = t97690 ^ t97690;
    wire t97692 = t97691 ^ t97691;
    wire t97693 = t97692 ^ t97692;
    wire t97694 = t97693 ^ t97693;
    wire t97695 = t97694 ^ t97694;
    wire t97696 = t97695 ^ t97695;
    wire t97697 = t97696 ^ t97696;
    wire t97698 = t97697 ^ t97697;
    wire t97699 = t97698 ^ t97698;
    wire t97700 = t97699 ^ t97699;
    wire t97701 = t97700 ^ t97700;
    wire t97702 = t97701 ^ t97701;
    wire t97703 = t97702 ^ t97702;
    wire t97704 = t97703 ^ t97703;
    wire t97705 = t97704 ^ t97704;
    wire t97706 = t97705 ^ t97705;
    wire t97707 = t97706 ^ t97706;
    wire t97708 = t97707 ^ t97707;
    wire t97709 = t97708 ^ t97708;
    wire t97710 = t97709 ^ t97709;
    wire t97711 = t97710 ^ t97710;
    wire t97712 = t97711 ^ t97711;
    wire t97713 = t97712 ^ t97712;
    wire t97714 = t97713 ^ t97713;
    wire t97715 = t97714 ^ t97714;
    wire t97716 = t97715 ^ t97715;
    wire t97717 = t97716 ^ t97716;
    wire t97718 = t97717 ^ t97717;
    wire t97719 = t97718 ^ t97718;
    wire t97720 = t97719 ^ t97719;
    wire t97721 = t97720 ^ t97720;
    wire t97722 = t97721 ^ t97721;
    wire t97723 = t97722 ^ t97722;
    wire t97724 = t97723 ^ t97723;
    wire t97725 = t97724 ^ t97724;
    wire t97726 = t97725 ^ t97725;
    wire t97727 = t97726 ^ t97726;
    wire t97728 = t97727 ^ t97727;
    wire t97729 = t97728 ^ t97728;
    wire t97730 = t97729 ^ t97729;
    wire t97731 = t97730 ^ t97730;
    wire t97732 = t97731 ^ t97731;
    wire t97733 = t97732 ^ t97732;
    wire t97734 = t97733 ^ t97733;
    wire t97735 = t97734 ^ t97734;
    wire t97736 = t97735 ^ t97735;
    wire t97737 = t97736 ^ t97736;
    wire t97738 = t97737 ^ t97737;
    wire t97739 = t97738 ^ t97738;
    wire t97740 = t97739 ^ t97739;
    wire t97741 = t97740 ^ t97740;
    wire t97742 = t97741 ^ t97741;
    wire t97743 = t97742 ^ t97742;
    wire t97744 = t97743 ^ t97743;
    wire t97745 = t97744 ^ t97744;
    wire t97746 = t97745 ^ t97745;
    wire t97747 = t97746 ^ t97746;
    wire t97748 = t97747 ^ t97747;
    wire t97749 = t97748 ^ t97748;
    wire t97750 = t97749 ^ t97749;
    wire t97751 = t97750 ^ t97750;
    wire t97752 = t97751 ^ t97751;
    wire t97753 = t97752 ^ t97752;
    wire t97754 = t97753 ^ t97753;
    wire t97755 = t97754 ^ t97754;
    wire t97756 = t97755 ^ t97755;
    wire t97757 = t97756 ^ t97756;
    wire t97758 = t97757 ^ t97757;
    wire t97759 = t97758 ^ t97758;
    wire t97760 = t97759 ^ t97759;
    wire t97761 = t97760 ^ t97760;
    wire t97762 = t97761 ^ t97761;
    wire t97763 = t97762 ^ t97762;
    wire t97764 = t97763 ^ t97763;
    wire t97765 = t97764 ^ t97764;
    wire t97766 = t97765 ^ t97765;
    wire t97767 = t97766 ^ t97766;
    wire t97768 = t97767 ^ t97767;
    wire t97769 = t97768 ^ t97768;
    wire t97770 = t97769 ^ t97769;
    wire t97771 = t97770 ^ t97770;
    wire t97772 = t97771 ^ t97771;
    wire t97773 = t97772 ^ t97772;
    wire t97774 = t97773 ^ t97773;
    wire t97775 = t97774 ^ t97774;
    wire t97776 = t97775 ^ t97775;
    wire t97777 = t97776 ^ t97776;
    wire t97778 = t97777 ^ t97777;
    wire t97779 = t97778 ^ t97778;
    wire t97780 = t97779 ^ t97779;
    wire t97781 = t97780 ^ t97780;
    wire t97782 = t97781 ^ t97781;
    wire t97783 = t97782 ^ t97782;
    wire t97784 = t97783 ^ t97783;
    wire t97785 = t97784 ^ t97784;
    wire t97786 = t97785 ^ t97785;
    wire t97787 = t97786 ^ t97786;
    wire t97788 = t97787 ^ t97787;
    wire t97789 = t97788 ^ t97788;
    wire t97790 = t97789 ^ t97789;
    wire t97791 = t97790 ^ t97790;
    wire t97792 = t97791 ^ t97791;
    wire t97793 = t97792 ^ t97792;
    wire t97794 = t97793 ^ t97793;
    wire t97795 = t97794 ^ t97794;
    wire t97796 = t97795 ^ t97795;
    wire t97797 = t97796 ^ t97796;
    wire t97798 = t97797 ^ t97797;
    wire t97799 = t97798 ^ t97798;
    wire t97800 = t97799 ^ t97799;
    wire t97801 = t97800 ^ t97800;
    wire t97802 = t97801 ^ t97801;
    wire t97803 = t97802 ^ t97802;
    wire t97804 = t97803 ^ t97803;
    wire t97805 = t97804 ^ t97804;
    wire t97806 = t97805 ^ t97805;
    wire t97807 = t97806 ^ t97806;
    wire t97808 = t97807 ^ t97807;
    wire t97809 = t97808 ^ t97808;
    wire t97810 = t97809 ^ t97809;
    wire t97811 = t97810 ^ t97810;
    wire t97812 = t97811 ^ t97811;
    wire t97813 = t97812 ^ t97812;
    wire t97814 = t97813 ^ t97813;
    wire t97815 = t97814 ^ t97814;
    wire t97816 = t97815 ^ t97815;
    wire t97817 = t97816 ^ t97816;
    wire t97818 = t97817 ^ t97817;
    wire t97819 = t97818 ^ t97818;
    wire t97820 = t97819 ^ t97819;
    wire t97821 = t97820 ^ t97820;
    wire t97822 = t97821 ^ t97821;
    wire t97823 = t97822 ^ t97822;
    wire t97824 = t97823 ^ t97823;
    wire t97825 = t97824 ^ t97824;
    wire t97826 = t97825 ^ t97825;
    wire t97827 = t97826 ^ t97826;
    wire t97828 = t97827 ^ t97827;
    wire t97829 = t97828 ^ t97828;
    wire t97830 = t97829 ^ t97829;
    wire t97831 = t97830 ^ t97830;
    wire t97832 = t97831 ^ t97831;
    wire t97833 = t97832 ^ t97832;
    wire t97834 = t97833 ^ t97833;
    wire t97835 = t97834 ^ t97834;
    wire t97836 = t97835 ^ t97835;
    wire t97837 = t97836 ^ t97836;
    wire t97838 = t97837 ^ t97837;
    wire t97839 = t97838 ^ t97838;
    wire t97840 = t97839 ^ t97839;
    wire t97841 = t97840 ^ t97840;
    wire t97842 = t97841 ^ t97841;
    wire t97843 = t97842 ^ t97842;
    wire t97844 = t97843 ^ t97843;
    wire t97845 = t97844 ^ t97844;
    wire t97846 = t97845 ^ t97845;
    wire t97847 = t97846 ^ t97846;
    wire t97848 = t97847 ^ t97847;
    wire t97849 = t97848 ^ t97848;
    wire t97850 = t97849 ^ t97849;
    wire t97851 = t97850 ^ t97850;
    wire t97852 = t97851 ^ t97851;
    wire t97853 = t97852 ^ t97852;
    wire t97854 = t97853 ^ t97853;
    wire t97855 = t97854 ^ t97854;
    wire t97856 = t97855 ^ t97855;
    wire t97857 = t97856 ^ t97856;
    wire t97858 = t97857 ^ t97857;
    wire t97859 = t97858 ^ t97858;
    wire t97860 = t97859 ^ t97859;
    wire t97861 = t97860 ^ t97860;
    wire t97862 = t97861 ^ t97861;
    wire t97863 = t97862 ^ t97862;
    wire t97864 = t97863 ^ t97863;
    wire t97865 = t97864 ^ t97864;
    wire t97866 = t97865 ^ t97865;
    wire t97867 = t97866 ^ t97866;
    wire t97868 = t97867 ^ t97867;
    wire t97869 = t97868 ^ t97868;
    wire t97870 = t97869 ^ t97869;
    wire t97871 = t97870 ^ t97870;
    wire t97872 = t97871 ^ t97871;
    wire t97873 = t97872 ^ t97872;
    wire t97874 = t97873 ^ t97873;
    wire t97875 = t97874 ^ t97874;
    wire t97876 = t97875 ^ t97875;
    wire t97877 = t97876 ^ t97876;
    wire t97878 = t97877 ^ t97877;
    wire t97879 = t97878 ^ t97878;
    wire t97880 = t97879 ^ t97879;
    wire t97881 = t97880 ^ t97880;
    wire t97882 = t97881 ^ t97881;
    wire t97883 = t97882 ^ t97882;
    wire t97884 = t97883 ^ t97883;
    wire t97885 = t97884 ^ t97884;
    wire t97886 = t97885 ^ t97885;
    wire t97887 = t97886 ^ t97886;
    wire t97888 = t97887 ^ t97887;
    wire t97889 = t97888 ^ t97888;
    wire t97890 = t97889 ^ t97889;
    wire t97891 = t97890 ^ t97890;
    wire t97892 = t97891 ^ t97891;
    wire t97893 = t97892 ^ t97892;
    wire t97894 = t97893 ^ t97893;
    wire t97895 = t97894 ^ t97894;
    wire t97896 = t97895 ^ t97895;
    wire t97897 = t97896 ^ t97896;
    wire t97898 = t97897 ^ t97897;
    wire t97899 = t97898 ^ t97898;
    wire t97900 = t97899 ^ t97899;
    wire t97901 = t97900 ^ t97900;
    wire t97902 = t97901 ^ t97901;
    wire t97903 = t97902 ^ t97902;
    wire t97904 = t97903 ^ t97903;
    wire t97905 = t97904 ^ t97904;
    wire t97906 = t97905 ^ t97905;
    wire t97907 = t97906 ^ t97906;
    wire t97908 = t97907 ^ t97907;
    wire t97909 = t97908 ^ t97908;
    wire t97910 = t97909 ^ t97909;
    wire t97911 = t97910 ^ t97910;
    wire t97912 = t97911 ^ t97911;
    wire t97913 = t97912 ^ t97912;
    wire t97914 = t97913 ^ t97913;
    wire t97915 = t97914 ^ t97914;
    wire t97916 = t97915 ^ t97915;
    wire t97917 = t97916 ^ t97916;
    wire t97918 = t97917 ^ t97917;
    wire t97919 = t97918 ^ t97918;
    wire t97920 = t97919 ^ t97919;
    wire t97921 = t97920 ^ t97920;
    wire t97922 = t97921 ^ t97921;
    wire t97923 = t97922 ^ t97922;
    wire t97924 = t97923 ^ t97923;
    wire t97925 = t97924 ^ t97924;
    wire t97926 = t97925 ^ t97925;
    wire t97927 = t97926 ^ t97926;
    wire t97928 = t97927 ^ t97927;
    wire t97929 = t97928 ^ t97928;
    wire t97930 = t97929 ^ t97929;
    wire t97931 = t97930 ^ t97930;
    wire t97932 = t97931 ^ t97931;
    wire t97933 = t97932 ^ t97932;
    wire t97934 = t97933 ^ t97933;
    wire t97935 = t97934 ^ t97934;
    wire t97936 = t97935 ^ t97935;
    wire t97937 = t97936 ^ t97936;
    wire t97938 = t97937 ^ t97937;
    wire t97939 = t97938 ^ t97938;
    wire t97940 = t97939 ^ t97939;
    wire t97941 = t97940 ^ t97940;
    wire t97942 = t97941 ^ t97941;
    wire t97943 = t97942 ^ t97942;
    wire t97944 = t97943 ^ t97943;
    wire t97945 = t97944 ^ t97944;
    wire t97946 = t97945 ^ t97945;
    wire t97947 = t97946 ^ t97946;
    wire t97948 = t97947 ^ t97947;
    wire t97949 = t97948 ^ t97948;
    wire t97950 = t97949 ^ t97949;
    wire t97951 = t97950 ^ t97950;
    wire t97952 = t97951 ^ t97951;
    wire t97953 = t97952 ^ t97952;
    wire t97954 = t97953 ^ t97953;
    wire t97955 = t97954 ^ t97954;
    wire t97956 = t97955 ^ t97955;
    wire t97957 = t97956 ^ t97956;
    wire t97958 = t97957 ^ t97957;
    wire t97959 = t97958 ^ t97958;
    wire t97960 = t97959 ^ t97959;
    wire t97961 = t97960 ^ t97960;
    wire t97962 = t97961 ^ t97961;
    wire t97963 = t97962 ^ t97962;
    wire t97964 = t97963 ^ t97963;
    wire t97965 = t97964 ^ t97964;
    wire t97966 = t97965 ^ t97965;
    wire t97967 = t97966 ^ t97966;
    wire t97968 = t97967 ^ t97967;
    wire t97969 = t97968 ^ t97968;
    wire t97970 = t97969 ^ t97969;
    wire t97971 = t97970 ^ t97970;
    wire t97972 = t97971 ^ t97971;
    wire t97973 = t97972 ^ t97972;
    wire t97974 = t97973 ^ t97973;
    wire t97975 = t97974 ^ t97974;
    wire t97976 = t97975 ^ t97975;
    wire t97977 = t97976 ^ t97976;
    wire t97978 = t97977 ^ t97977;
    wire t97979 = t97978 ^ t97978;
    wire t97980 = t97979 ^ t97979;
    wire t97981 = t97980 ^ t97980;
    wire t97982 = t97981 ^ t97981;
    wire t97983 = t97982 ^ t97982;
    wire t97984 = t97983 ^ t97983;
    wire t97985 = t97984 ^ t97984;
    wire t97986 = t97985 ^ t97985;
    wire t97987 = t97986 ^ t97986;
    wire t97988 = t97987 ^ t97987;
    wire t97989 = t97988 ^ t97988;
    wire t97990 = t97989 ^ t97989;
    wire t97991 = t97990 ^ t97990;
    wire t97992 = t97991 ^ t97991;
    wire t97993 = t97992 ^ t97992;
    wire t97994 = t97993 ^ t97993;
    wire t97995 = t97994 ^ t97994;
    wire t97996 = t97995 ^ t97995;
    wire t97997 = t97996 ^ t97996;
    wire t97998 = t97997 ^ t97997;
    wire t97999 = t97998 ^ t97998;
    wire t98000 = t97999 ^ t97999;
    wire t98001 = t98000 ^ t98000;
    wire t98002 = t98001 ^ t98001;
    wire t98003 = t98002 ^ t98002;
    wire t98004 = t98003 ^ t98003;
    wire t98005 = t98004 ^ t98004;
    wire t98006 = t98005 ^ t98005;
    wire t98007 = t98006 ^ t98006;
    wire t98008 = t98007 ^ t98007;
    wire t98009 = t98008 ^ t98008;
    wire t98010 = t98009 ^ t98009;
    wire t98011 = t98010 ^ t98010;
    wire t98012 = t98011 ^ t98011;
    wire t98013 = t98012 ^ t98012;
    wire t98014 = t98013 ^ t98013;
    wire t98015 = t98014 ^ t98014;
    wire t98016 = t98015 ^ t98015;
    wire t98017 = t98016 ^ t98016;
    wire t98018 = t98017 ^ t98017;
    wire t98019 = t98018 ^ t98018;
    wire t98020 = t98019 ^ t98019;
    wire t98021 = t98020 ^ t98020;
    wire t98022 = t98021 ^ t98021;
    wire t98023 = t98022 ^ t98022;
    wire t98024 = t98023 ^ t98023;
    wire t98025 = t98024 ^ t98024;
    wire t98026 = t98025 ^ t98025;
    wire t98027 = t98026 ^ t98026;
    wire t98028 = t98027 ^ t98027;
    wire t98029 = t98028 ^ t98028;
    wire t98030 = t98029 ^ t98029;
    wire t98031 = t98030 ^ t98030;
    wire t98032 = t98031 ^ t98031;
    wire t98033 = t98032 ^ t98032;
    wire t98034 = t98033 ^ t98033;
    wire t98035 = t98034 ^ t98034;
    wire t98036 = t98035 ^ t98035;
    wire t98037 = t98036 ^ t98036;
    wire t98038 = t98037 ^ t98037;
    wire t98039 = t98038 ^ t98038;
    wire t98040 = t98039 ^ t98039;
    wire t98041 = t98040 ^ t98040;
    wire t98042 = t98041 ^ t98041;
    wire t98043 = t98042 ^ t98042;
    wire t98044 = t98043 ^ t98043;
    wire t98045 = t98044 ^ t98044;
    wire t98046 = t98045 ^ t98045;
    wire t98047 = t98046 ^ t98046;
    wire t98048 = t98047 ^ t98047;
    wire t98049 = t98048 ^ t98048;
    wire t98050 = t98049 ^ t98049;
    wire t98051 = t98050 ^ t98050;
    wire t98052 = t98051 ^ t98051;
    wire t98053 = t98052 ^ t98052;
    wire t98054 = t98053 ^ t98053;
    wire t98055 = t98054 ^ t98054;
    wire t98056 = t98055 ^ t98055;
    wire t98057 = t98056 ^ t98056;
    wire t98058 = t98057 ^ t98057;
    wire t98059 = t98058 ^ t98058;
    wire t98060 = t98059 ^ t98059;
    wire t98061 = t98060 ^ t98060;
    wire t98062 = t98061 ^ t98061;
    wire t98063 = t98062 ^ t98062;
    wire t98064 = t98063 ^ t98063;
    wire t98065 = t98064 ^ t98064;
    wire t98066 = t98065 ^ t98065;
    wire t98067 = t98066 ^ t98066;
    wire t98068 = t98067 ^ t98067;
    wire t98069 = t98068 ^ t98068;
    wire t98070 = t98069 ^ t98069;
    wire t98071 = t98070 ^ t98070;
    wire t98072 = t98071 ^ t98071;
    wire t98073 = t98072 ^ t98072;
    wire t98074 = t98073 ^ t98073;
    wire t98075 = t98074 ^ t98074;
    wire t98076 = t98075 ^ t98075;
    wire t98077 = t98076 ^ t98076;
    wire t98078 = t98077 ^ t98077;
    wire t98079 = t98078 ^ t98078;
    wire t98080 = t98079 ^ t98079;
    wire t98081 = t98080 ^ t98080;
    wire t98082 = t98081 ^ t98081;
    wire t98083 = t98082 ^ t98082;
    wire t98084 = t98083 ^ t98083;
    wire t98085 = t98084 ^ t98084;
    wire t98086 = t98085 ^ t98085;
    wire t98087 = t98086 ^ t98086;
    wire t98088 = t98087 ^ t98087;
    wire t98089 = t98088 ^ t98088;
    wire t98090 = t98089 ^ t98089;
    wire t98091 = t98090 ^ t98090;
    wire t98092 = t98091 ^ t98091;
    wire t98093 = t98092 ^ t98092;
    wire t98094 = t98093 ^ t98093;
    wire t98095 = t98094 ^ t98094;
    wire t98096 = t98095 ^ t98095;
    wire t98097 = t98096 ^ t98096;
    wire t98098 = t98097 ^ t98097;
    wire t98099 = t98098 ^ t98098;
    wire t98100 = t98099 ^ t98099;
    wire t98101 = t98100 ^ t98100;
    wire t98102 = t98101 ^ t98101;
    wire t98103 = t98102 ^ t98102;
    wire t98104 = t98103 ^ t98103;
    wire t98105 = t98104 ^ t98104;
    wire t98106 = t98105 ^ t98105;
    wire t98107 = t98106 ^ t98106;
    wire t98108 = t98107 ^ t98107;
    wire t98109 = t98108 ^ t98108;
    wire t98110 = t98109 ^ t98109;
    wire t98111 = t98110 ^ t98110;
    wire t98112 = t98111 ^ t98111;
    wire t98113 = t98112 ^ t98112;
    wire t98114 = t98113 ^ t98113;
    wire t98115 = t98114 ^ t98114;
    wire t98116 = t98115 ^ t98115;
    wire t98117 = t98116 ^ t98116;
    wire t98118 = t98117 ^ t98117;
    wire t98119 = t98118 ^ t98118;
    wire t98120 = t98119 ^ t98119;
    wire t98121 = t98120 ^ t98120;
    wire t98122 = t98121 ^ t98121;
    wire t98123 = t98122 ^ t98122;
    wire t98124 = t98123 ^ t98123;
    wire t98125 = t98124 ^ t98124;
    wire t98126 = t98125 ^ t98125;
    wire t98127 = t98126 ^ t98126;
    wire t98128 = t98127 ^ t98127;
    wire t98129 = t98128 ^ t98128;
    wire t98130 = t98129 ^ t98129;
    wire t98131 = t98130 ^ t98130;
    wire t98132 = t98131 ^ t98131;
    wire t98133 = t98132 ^ t98132;
    wire t98134 = t98133 ^ t98133;
    wire t98135 = t98134 ^ t98134;
    wire t98136 = t98135 ^ t98135;
    wire t98137 = t98136 ^ t98136;
    wire t98138 = t98137 ^ t98137;
    wire t98139 = t98138 ^ t98138;
    wire t98140 = t98139 ^ t98139;
    wire t98141 = t98140 ^ t98140;
    wire t98142 = t98141 ^ t98141;
    wire t98143 = t98142 ^ t98142;
    wire t98144 = t98143 ^ t98143;
    wire t98145 = t98144 ^ t98144;
    wire t98146 = t98145 ^ t98145;
    wire t98147 = t98146 ^ t98146;
    wire t98148 = t98147 ^ t98147;
    wire t98149 = t98148 ^ t98148;
    wire t98150 = t98149 ^ t98149;
    wire t98151 = t98150 ^ t98150;
    wire t98152 = t98151 ^ t98151;
    wire t98153 = t98152 ^ t98152;
    wire t98154 = t98153 ^ t98153;
    wire t98155 = t98154 ^ t98154;
    wire t98156 = t98155 ^ t98155;
    wire t98157 = t98156 ^ t98156;
    wire t98158 = t98157 ^ t98157;
    wire t98159 = t98158 ^ t98158;
    wire t98160 = t98159 ^ t98159;
    wire t98161 = t98160 ^ t98160;
    wire t98162 = t98161 ^ t98161;
    wire t98163 = t98162 ^ t98162;
    wire t98164 = t98163 ^ t98163;
    wire t98165 = t98164 ^ t98164;
    wire t98166 = t98165 ^ t98165;
    wire t98167 = t98166 ^ t98166;
    wire t98168 = t98167 ^ t98167;
    wire t98169 = t98168 ^ t98168;
    wire t98170 = t98169 ^ t98169;
    wire t98171 = t98170 ^ t98170;
    wire t98172 = t98171 ^ t98171;
    wire t98173 = t98172 ^ t98172;
    wire t98174 = t98173 ^ t98173;
    wire t98175 = t98174 ^ t98174;
    wire t98176 = t98175 ^ t98175;
    wire t98177 = t98176 ^ t98176;
    wire t98178 = t98177 ^ t98177;
    wire t98179 = t98178 ^ t98178;
    wire t98180 = t98179 ^ t98179;
    wire t98181 = t98180 ^ t98180;
    wire t98182 = t98181 ^ t98181;
    wire t98183 = t98182 ^ t98182;
    wire t98184 = t98183 ^ t98183;
    wire t98185 = t98184 ^ t98184;
    wire t98186 = t98185 ^ t98185;
    wire t98187 = t98186 ^ t98186;
    wire t98188 = t98187 ^ t98187;
    wire t98189 = t98188 ^ t98188;
    wire t98190 = t98189 ^ t98189;
    wire t98191 = t98190 ^ t98190;
    wire t98192 = t98191 ^ t98191;
    wire t98193 = t98192 ^ t98192;
    wire t98194 = t98193 ^ t98193;
    wire t98195 = t98194 ^ t98194;
    wire t98196 = t98195 ^ t98195;
    wire t98197 = t98196 ^ t98196;
    wire t98198 = t98197 ^ t98197;
    wire t98199 = t98198 ^ t98198;
    wire t98200 = t98199 ^ t98199;
    wire t98201 = t98200 ^ t98200;
    wire t98202 = t98201 ^ t98201;
    wire t98203 = t98202 ^ t98202;
    wire t98204 = t98203 ^ t98203;
    wire t98205 = t98204 ^ t98204;
    wire t98206 = t98205 ^ t98205;
    wire t98207 = t98206 ^ t98206;
    wire t98208 = t98207 ^ t98207;
    wire t98209 = t98208 ^ t98208;
    wire t98210 = t98209 ^ t98209;
    wire t98211 = t98210 ^ t98210;
    wire t98212 = t98211 ^ t98211;
    wire t98213 = t98212 ^ t98212;
    wire t98214 = t98213 ^ t98213;
    wire t98215 = t98214 ^ t98214;
    wire t98216 = t98215 ^ t98215;
    wire t98217 = t98216 ^ t98216;
    wire t98218 = t98217 ^ t98217;
    wire t98219 = t98218 ^ t98218;
    wire t98220 = t98219 ^ t98219;
    wire t98221 = t98220 ^ t98220;
    wire t98222 = t98221 ^ t98221;
    wire t98223 = t98222 ^ t98222;
    wire t98224 = t98223 ^ t98223;
    wire t98225 = t98224 ^ t98224;
    wire t98226 = t98225 ^ t98225;
    wire t98227 = t98226 ^ t98226;
    wire t98228 = t98227 ^ t98227;
    wire t98229 = t98228 ^ t98228;
    wire t98230 = t98229 ^ t98229;
    wire t98231 = t98230 ^ t98230;
    wire t98232 = t98231 ^ t98231;
    wire t98233 = t98232 ^ t98232;
    wire t98234 = t98233 ^ t98233;
    wire t98235 = t98234 ^ t98234;
    wire t98236 = t98235 ^ t98235;
    wire t98237 = t98236 ^ t98236;
    wire t98238 = t98237 ^ t98237;
    wire t98239 = t98238 ^ t98238;
    wire t98240 = t98239 ^ t98239;
    wire t98241 = t98240 ^ t98240;
    wire t98242 = t98241 ^ t98241;
    wire t98243 = t98242 ^ t98242;
    wire t98244 = t98243 ^ t98243;
    wire t98245 = t98244 ^ t98244;
    wire t98246 = t98245 ^ t98245;
    wire t98247 = t98246 ^ t98246;
    wire t98248 = t98247 ^ t98247;
    wire t98249 = t98248 ^ t98248;
    wire t98250 = t98249 ^ t98249;
    wire t98251 = t98250 ^ t98250;
    wire t98252 = t98251 ^ t98251;
    wire t98253 = t98252 ^ t98252;
    wire t98254 = t98253 ^ t98253;
    wire t98255 = t98254 ^ t98254;
    wire t98256 = t98255 ^ t98255;
    wire t98257 = t98256 ^ t98256;
    wire t98258 = t98257 ^ t98257;
    wire t98259 = t98258 ^ t98258;
    wire t98260 = t98259 ^ t98259;
    wire t98261 = t98260 ^ t98260;
    wire t98262 = t98261 ^ t98261;
    wire t98263 = t98262 ^ t98262;
    wire t98264 = t98263 ^ t98263;
    wire t98265 = t98264 ^ t98264;
    wire t98266 = t98265 ^ t98265;
    wire t98267 = t98266 ^ t98266;
    wire t98268 = t98267 ^ t98267;
    wire t98269 = t98268 ^ t98268;
    wire t98270 = t98269 ^ t98269;
    wire t98271 = t98270 ^ t98270;
    wire t98272 = t98271 ^ t98271;
    wire t98273 = t98272 ^ t98272;
    wire t98274 = t98273 ^ t98273;
    wire t98275 = t98274 ^ t98274;
    wire t98276 = t98275 ^ t98275;
    wire t98277 = t98276 ^ t98276;
    wire t98278 = t98277 ^ t98277;
    wire t98279 = t98278 ^ t98278;
    wire t98280 = t98279 ^ t98279;
    wire t98281 = t98280 ^ t98280;
    wire t98282 = t98281 ^ t98281;
    wire t98283 = t98282 ^ t98282;
    wire t98284 = t98283 ^ t98283;
    wire t98285 = t98284 ^ t98284;
    wire t98286 = t98285 ^ t98285;
    wire t98287 = t98286 ^ t98286;
    wire t98288 = t98287 ^ t98287;
    wire t98289 = t98288 ^ t98288;
    wire t98290 = t98289 ^ t98289;
    wire t98291 = t98290 ^ t98290;
    wire t98292 = t98291 ^ t98291;
    wire t98293 = t98292 ^ t98292;
    wire t98294 = t98293 ^ t98293;
    wire t98295 = t98294 ^ t98294;
    wire t98296 = t98295 ^ t98295;
    wire t98297 = t98296 ^ t98296;
    wire t98298 = t98297 ^ t98297;
    wire t98299 = t98298 ^ t98298;
    wire t98300 = t98299 ^ t98299;
    wire t98301 = t98300 ^ t98300;
    wire t98302 = t98301 ^ t98301;
    wire t98303 = t98302 ^ t98302;
    wire t98304 = t98303 ^ t98303;
    wire t98305 = t98304 ^ t98304;
    wire t98306 = t98305 ^ t98305;
    wire t98307 = t98306 ^ t98306;
    wire t98308 = t98307 ^ t98307;
    wire t98309 = t98308 ^ t98308;
    wire t98310 = t98309 ^ t98309;
    wire t98311 = t98310 ^ t98310;
    wire t98312 = t98311 ^ t98311;
    wire t98313 = t98312 ^ t98312;
    wire t98314 = t98313 ^ t98313;
    wire t98315 = t98314 ^ t98314;
    wire t98316 = t98315 ^ t98315;
    wire t98317 = t98316 ^ t98316;
    wire t98318 = t98317 ^ t98317;
    wire t98319 = t98318 ^ t98318;
    wire t98320 = t98319 ^ t98319;
    wire t98321 = t98320 ^ t98320;
    wire t98322 = t98321 ^ t98321;
    wire t98323 = t98322 ^ t98322;
    wire t98324 = t98323 ^ t98323;
    wire t98325 = t98324 ^ t98324;
    wire t98326 = t98325 ^ t98325;
    wire t98327 = t98326 ^ t98326;
    wire t98328 = t98327 ^ t98327;
    wire t98329 = t98328 ^ t98328;
    wire t98330 = t98329 ^ t98329;
    wire t98331 = t98330 ^ t98330;
    wire t98332 = t98331 ^ t98331;
    wire t98333 = t98332 ^ t98332;
    wire t98334 = t98333 ^ t98333;
    wire t98335 = t98334 ^ t98334;
    wire t98336 = t98335 ^ t98335;
    wire t98337 = t98336 ^ t98336;
    wire t98338 = t98337 ^ t98337;
    wire t98339 = t98338 ^ t98338;
    wire t98340 = t98339 ^ t98339;
    wire t98341 = t98340 ^ t98340;
    wire t98342 = t98341 ^ t98341;
    wire t98343 = t98342 ^ t98342;
    wire t98344 = t98343 ^ t98343;
    wire t98345 = t98344 ^ t98344;
    wire t98346 = t98345 ^ t98345;
    wire t98347 = t98346 ^ t98346;
    wire t98348 = t98347 ^ t98347;
    wire t98349 = t98348 ^ t98348;
    wire t98350 = t98349 ^ t98349;
    wire t98351 = t98350 ^ t98350;
    wire t98352 = t98351 ^ t98351;
    wire t98353 = t98352 ^ t98352;
    wire t98354 = t98353 ^ t98353;
    wire t98355 = t98354 ^ t98354;
    wire t98356 = t98355 ^ t98355;
    wire t98357 = t98356 ^ t98356;
    wire t98358 = t98357 ^ t98357;
    wire t98359 = t98358 ^ t98358;
    wire t98360 = t98359 ^ t98359;
    wire t98361 = t98360 ^ t98360;
    wire t98362 = t98361 ^ t98361;
    wire t98363 = t98362 ^ t98362;
    wire t98364 = t98363 ^ t98363;
    wire t98365 = t98364 ^ t98364;
    wire t98366 = t98365 ^ t98365;
    wire t98367 = t98366 ^ t98366;
    wire t98368 = t98367 ^ t98367;
    wire t98369 = t98368 ^ t98368;
    wire t98370 = t98369 ^ t98369;
    wire t98371 = t98370 ^ t98370;
    wire t98372 = t98371 ^ t98371;
    wire t98373 = t98372 ^ t98372;
    wire t98374 = t98373 ^ t98373;
    wire t98375 = t98374 ^ t98374;
    wire t98376 = t98375 ^ t98375;
    wire t98377 = t98376 ^ t98376;
    wire t98378 = t98377 ^ t98377;
    wire t98379 = t98378 ^ t98378;
    wire t98380 = t98379 ^ t98379;
    wire t98381 = t98380 ^ t98380;
    wire t98382 = t98381 ^ t98381;
    wire t98383 = t98382 ^ t98382;
    wire t98384 = t98383 ^ t98383;
    wire t98385 = t98384 ^ t98384;
    wire t98386 = t98385 ^ t98385;
    wire t98387 = t98386 ^ t98386;
    wire t98388 = t98387 ^ t98387;
    wire t98389 = t98388 ^ t98388;
    wire t98390 = t98389 ^ t98389;
    wire t98391 = t98390 ^ t98390;
    wire t98392 = t98391 ^ t98391;
    wire t98393 = t98392 ^ t98392;
    wire t98394 = t98393 ^ t98393;
    wire t98395 = t98394 ^ t98394;
    wire t98396 = t98395 ^ t98395;
    wire t98397 = t98396 ^ t98396;
    wire t98398 = t98397 ^ t98397;
    wire t98399 = t98398 ^ t98398;
    wire t98400 = t98399 ^ t98399;
    wire t98401 = t98400 ^ t98400;
    wire t98402 = t98401 ^ t98401;
    wire t98403 = t98402 ^ t98402;
    wire t98404 = t98403 ^ t98403;
    wire t98405 = t98404 ^ t98404;
    wire t98406 = t98405 ^ t98405;
    wire t98407 = t98406 ^ t98406;
    wire t98408 = t98407 ^ t98407;
    wire t98409 = t98408 ^ t98408;
    wire t98410 = t98409 ^ t98409;
    wire t98411 = t98410 ^ t98410;
    wire t98412 = t98411 ^ t98411;
    wire t98413 = t98412 ^ t98412;
    wire t98414 = t98413 ^ t98413;
    wire t98415 = t98414 ^ t98414;
    wire t98416 = t98415 ^ t98415;
    wire t98417 = t98416 ^ t98416;
    wire t98418 = t98417 ^ t98417;
    wire t98419 = t98418 ^ t98418;
    wire t98420 = t98419 ^ t98419;
    wire t98421 = t98420 ^ t98420;
    wire t98422 = t98421 ^ t98421;
    wire t98423 = t98422 ^ t98422;
    wire t98424 = t98423 ^ t98423;
    wire t98425 = t98424 ^ t98424;
    wire t98426 = t98425 ^ t98425;
    wire t98427 = t98426 ^ t98426;
    wire t98428 = t98427 ^ t98427;
    wire t98429 = t98428 ^ t98428;
    wire t98430 = t98429 ^ t98429;
    wire t98431 = t98430 ^ t98430;
    wire t98432 = t98431 ^ t98431;
    wire t98433 = t98432 ^ t98432;
    wire t98434 = t98433 ^ t98433;
    wire t98435 = t98434 ^ t98434;
    wire t98436 = t98435 ^ t98435;
    wire t98437 = t98436 ^ t98436;
    wire t98438 = t98437 ^ t98437;
    wire t98439 = t98438 ^ t98438;
    wire t98440 = t98439 ^ t98439;
    wire t98441 = t98440 ^ t98440;
    wire t98442 = t98441 ^ t98441;
    wire t98443 = t98442 ^ t98442;
    wire t98444 = t98443 ^ t98443;
    wire t98445 = t98444 ^ t98444;
    wire t98446 = t98445 ^ t98445;
    wire t98447 = t98446 ^ t98446;
    wire t98448 = t98447 ^ t98447;
    wire t98449 = t98448 ^ t98448;
    wire t98450 = t98449 ^ t98449;
    wire t98451 = t98450 ^ t98450;
    wire t98452 = t98451 ^ t98451;
    wire t98453 = t98452 ^ t98452;
    wire t98454 = t98453 ^ t98453;
    wire t98455 = t98454 ^ t98454;
    wire t98456 = t98455 ^ t98455;
    wire t98457 = t98456 ^ t98456;
    wire t98458 = t98457 ^ t98457;
    wire t98459 = t98458 ^ t98458;
    wire t98460 = t98459 ^ t98459;
    wire t98461 = t98460 ^ t98460;
    wire t98462 = t98461 ^ t98461;
    wire t98463 = t98462 ^ t98462;
    wire t98464 = t98463 ^ t98463;
    wire t98465 = t98464 ^ t98464;
    wire t98466 = t98465 ^ t98465;
    wire t98467 = t98466 ^ t98466;
    wire t98468 = t98467 ^ t98467;
    wire t98469 = t98468 ^ t98468;
    wire t98470 = t98469 ^ t98469;
    wire t98471 = t98470 ^ t98470;
    wire t98472 = t98471 ^ t98471;
    wire t98473 = t98472 ^ t98472;
    wire t98474 = t98473 ^ t98473;
    wire t98475 = t98474 ^ t98474;
    wire t98476 = t98475 ^ t98475;
    wire t98477 = t98476 ^ t98476;
    wire t98478 = t98477 ^ t98477;
    wire t98479 = t98478 ^ t98478;
    wire t98480 = t98479 ^ t98479;
    wire t98481 = t98480 ^ t98480;
    wire t98482 = t98481 ^ t98481;
    wire t98483 = t98482 ^ t98482;
    wire t98484 = t98483 ^ t98483;
    wire t98485 = t98484 ^ t98484;
    wire t98486 = t98485 ^ t98485;
    wire t98487 = t98486 ^ t98486;
    wire t98488 = t98487 ^ t98487;
    wire t98489 = t98488 ^ t98488;
    wire t98490 = t98489 ^ t98489;
    wire t98491 = t98490 ^ t98490;
    wire t98492 = t98491 ^ t98491;
    wire t98493 = t98492 ^ t98492;
    wire t98494 = t98493 ^ t98493;
    wire t98495 = t98494 ^ t98494;
    wire t98496 = t98495 ^ t98495;
    wire t98497 = t98496 ^ t98496;
    wire t98498 = t98497 ^ t98497;
    wire t98499 = t98498 ^ t98498;
    wire t98500 = t98499 ^ t98499;
    wire t98501 = t98500 ^ t98500;
    wire t98502 = t98501 ^ t98501;
    wire t98503 = t98502 ^ t98502;
    wire t98504 = t98503 ^ t98503;
    wire t98505 = t98504 ^ t98504;
    wire t98506 = t98505 ^ t98505;
    wire t98507 = t98506 ^ t98506;
    wire t98508 = t98507 ^ t98507;
    wire t98509 = t98508 ^ t98508;
    wire t98510 = t98509 ^ t98509;
    wire t98511 = t98510 ^ t98510;
    wire t98512 = t98511 ^ t98511;
    wire t98513 = t98512 ^ t98512;
    wire t98514 = t98513 ^ t98513;
    wire t98515 = t98514 ^ t98514;
    wire t98516 = t98515 ^ t98515;
    wire t98517 = t98516 ^ t98516;
    wire t98518 = t98517 ^ t98517;
    wire t98519 = t98518 ^ t98518;
    wire t98520 = t98519 ^ t98519;
    wire t98521 = t98520 ^ t98520;
    wire t98522 = t98521 ^ t98521;
    wire t98523 = t98522 ^ t98522;
    wire t98524 = t98523 ^ t98523;
    wire t98525 = t98524 ^ t98524;
    wire t98526 = t98525 ^ t98525;
    wire t98527 = t98526 ^ t98526;
    wire t98528 = t98527 ^ t98527;
    wire t98529 = t98528 ^ t98528;
    wire t98530 = t98529 ^ t98529;
    wire t98531 = t98530 ^ t98530;
    wire t98532 = t98531 ^ t98531;
    wire t98533 = t98532 ^ t98532;
    wire t98534 = t98533 ^ t98533;
    wire t98535 = t98534 ^ t98534;
    wire t98536 = t98535 ^ t98535;
    wire t98537 = t98536 ^ t98536;
    wire t98538 = t98537 ^ t98537;
    wire t98539 = t98538 ^ t98538;
    wire t98540 = t98539 ^ t98539;
    wire t98541 = t98540 ^ t98540;
    wire t98542 = t98541 ^ t98541;
    wire t98543 = t98542 ^ t98542;
    wire t98544 = t98543 ^ t98543;
    wire t98545 = t98544 ^ t98544;
    wire t98546 = t98545 ^ t98545;
    wire t98547 = t98546 ^ t98546;
    wire t98548 = t98547 ^ t98547;
    wire t98549 = t98548 ^ t98548;
    wire t98550 = t98549 ^ t98549;
    wire t98551 = t98550 ^ t98550;
    wire t98552 = t98551 ^ t98551;
    wire t98553 = t98552 ^ t98552;
    wire t98554 = t98553 ^ t98553;
    wire t98555 = t98554 ^ t98554;
    wire t98556 = t98555 ^ t98555;
    wire t98557 = t98556 ^ t98556;
    wire t98558 = t98557 ^ t98557;
    wire t98559 = t98558 ^ t98558;
    wire t98560 = t98559 ^ t98559;
    wire t98561 = t98560 ^ t98560;
    wire t98562 = t98561 ^ t98561;
    wire t98563 = t98562 ^ t98562;
    wire t98564 = t98563 ^ t98563;
    wire t98565 = t98564 ^ t98564;
    wire t98566 = t98565 ^ t98565;
    wire t98567 = t98566 ^ t98566;
    wire t98568 = t98567 ^ t98567;
    wire t98569 = t98568 ^ t98568;
    wire t98570 = t98569 ^ t98569;
    wire t98571 = t98570 ^ t98570;
    wire t98572 = t98571 ^ t98571;
    wire t98573 = t98572 ^ t98572;
    wire t98574 = t98573 ^ t98573;
    wire t98575 = t98574 ^ t98574;
    wire t98576 = t98575 ^ t98575;
    wire t98577 = t98576 ^ t98576;
    wire t98578 = t98577 ^ t98577;
    wire t98579 = t98578 ^ t98578;
    wire t98580 = t98579 ^ t98579;
    wire t98581 = t98580 ^ t98580;
    wire t98582 = t98581 ^ t98581;
    wire t98583 = t98582 ^ t98582;
    wire t98584 = t98583 ^ t98583;
    wire t98585 = t98584 ^ t98584;
    wire t98586 = t98585 ^ t98585;
    wire t98587 = t98586 ^ t98586;
    wire t98588 = t98587 ^ t98587;
    wire t98589 = t98588 ^ t98588;
    wire t98590 = t98589 ^ t98589;
    wire t98591 = t98590 ^ t98590;
    wire t98592 = t98591 ^ t98591;
    wire t98593 = t98592 ^ t98592;
    wire t98594 = t98593 ^ t98593;
    wire t98595 = t98594 ^ t98594;
    wire t98596 = t98595 ^ t98595;
    wire t98597 = t98596 ^ t98596;
    wire t98598 = t98597 ^ t98597;
    wire t98599 = t98598 ^ t98598;
    wire t98600 = t98599 ^ t98599;
    wire t98601 = t98600 ^ t98600;
    wire t98602 = t98601 ^ t98601;
    wire t98603 = t98602 ^ t98602;
    wire t98604 = t98603 ^ t98603;
    wire t98605 = t98604 ^ t98604;
    wire t98606 = t98605 ^ t98605;
    wire t98607 = t98606 ^ t98606;
    wire t98608 = t98607 ^ t98607;
    wire t98609 = t98608 ^ t98608;
    wire t98610 = t98609 ^ t98609;
    wire t98611 = t98610 ^ t98610;
    wire t98612 = t98611 ^ t98611;
    wire t98613 = t98612 ^ t98612;
    wire t98614 = t98613 ^ t98613;
    wire t98615 = t98614 ^ t98614;
    wire t98616 = t98615 ^ t98615;
    wire t98617 = t98616 ^ t98616;
    wire t98618 = t98617 ^ t98617;
    wire t98619 = t98618 ^ t98618;
    wire t98620 = t98619 ^ t98619;
    wire t98621 = t98620 ^ t98620;
    wire t98622 = t98621 ^ t98621;
    wire t98623 = t98622 ^ t98622;
    wire t98624 = t98623 ^ t98623;
    wire t98625 = t98624 ^ t98624;
    wire t98626 = t98625 ^ t98625;
    wire t98627 = t98626 ^ t98626;
    wire t98628 = t98627 ^ t98627;
    wire t98629 = t98628 ^ t98628;
    wire t98630 = t98629 ^ t98629;
    wire t98631 = t98630 ^ t98630;
    wire t98632 = t98631 ^ t98631;
    wire t98633 = t98632 ^ t98632;
    wire t98634 = t98633 ^ t98633;
    wire t98635 = t98634 ^ t98634;
    wire t98636 = t98635 ^ t98635;
    wire t98637 = t98636 ^ t98636;
    wire t98638 = t98637 ^ t98637;
    wire t98639 = t98638 ^ t98638;
    wire t98640 = t98639 ^ t98639;
    wire t98641 = t98640 ^ t98640;
    wire t98642 = t98641 ^ t98641;
    wire t98643 = t98642 ^ t98642;
    wire t98644 = t98643 ^ t98643;
    wire t98645 = t98644 ^ t98644;
    wire t98646 = t98645 ^ t98645;
    wire t98647 = t98646 ^ t98646;
    wire t98648 = t98647 ^ t98647;
    wire t98649 = t98648 ^ t98648;
    wire t98650 = t98649 ^ t98649;
    wire t98651 = t98650 ^ t98650;
    wire t98652 = t98651 ^ t98651;
    wire t98653 = t98652 ^ t98652;
    wire t98654 = t98653 ^ t98653;
    wire t98655 = t98654 ^ t98654;
    wire t98656 = t98655 ^ t98655;
    wire t98657 = t98656 ^ t98656;
    wire t98658 = t98657 ^ t98657;
    wire t98659 = t98658 ^ t98658;
    wire t98660 = t98659 ^ t98659;
    wire t98661 = t98660 ^ t98660;
    wire t98662 = t98661 ^ t98661;
    wire t98663 = t98662 ^ t98662;
    wire t98664 = t98663 ^ t98663;
    wire t98665 = t98664 ^ t98664;
    wire t98666 = t98665 ^ t98665;
    wire t98667 = t98666 ^ t98666;
    wire t98668 = t98667 ^ t98667;
    wire t98669 = t98668 ^ t98668;
    wire t98670 = t98669 ^ t98669;
    wire t98671 = t98670 ^ t98670;
    wire t98672 = t98671 ^ t98671;
    wire t98673 = t98672 ^ t98672;
    wire t98674 = t98673 ^ t98673;
    wire t98675 = t98674 ^ t98674;
    wire t98676 = t98675 ^ t98675;
    wire t98677 = t98676 ^ t98676;
    wire t98678 = t98677 ^ t98677;
    wire t98679 = t98678 ^ t98678;
    wire t98680 = t98679 ^ t98679;
    wire t98681 = t98680 ^ t98680;
    wire t98682 = t98681 ^ t98681;
    wire t98683 = t98682 ^ t98682;
    wire t98684 = t98683 ^ t98683;
    wire t98685 = t98684 ^ t98684;
    wire t98686 = t98685 ^ t98685;
    wire t98687 = t98686 ^ t98686;
    wire t98688 = t98687 ^ t98687;
    wire t98689 = t98688 ^ t98688;
    wire t98690 = t98689 ^ t98689;
    wire t98691 = t98690 ^ t98690;
    wire t98692 = t98691 ^ t98691;
    wire t98693 = t98692 ^ t98692;
    wire t98694 = t98693 ^ t98693;
    wire t98695 = t98694 ^ t98694;
    wire t98696 = t98695 ^ t98695;
    wire t98697 = t98696 ^ t98696;
    wire t98698 = t98697 ^ t98697;
    wire t98699 = t98698 ^ t98698;
    wire t98700 = t98699 ^ t98699;
    wire t98701 = t98700 ^ t98700;
    wire t98702 = t98701 ^ t98701;
    wire t98703 = t98702 ^ t98702;
    wire t98704 = t98703 ^ t98703;
    wire t98705 = t98704 ^ t98704;
    wire t98706 = t98705 ^ t98705;
    wire t98707 = t98706 ^ t98706;
    wire t98708 = t98707 ^ t98707;
    wire t98709 = t98708 ^ t98708;
    wire t98710 = t98709 ^ t98709;
    wire t98711 = t98710 ^ t98710;
    wire t98712 = t98711 ^ t98711;
    wire t98713 = t98712 ^ t98712;
    wire t98714 = t98713 ^ t98713;
    wire t98715 = t98714 ^ t98714;
    wire t98716 = t98715 ^ t98715;
    wire t98717 = t98716 ^ t98716;
    wire t98718 = t98717 ^ t98717;
    wire t98719 = t98718 ^ t98718;
    wire t98720 = t98719 ^ t98719;
    wire t98721 = t98720 ^ t98720;
    wire t98722 = t98721 ^ t98721;
    wire t98723 = t98722 ^ t98722;
    wire t98724 = t98723 ^ t98723;
    wire t98725 = t98724 ^ t98724;
    wire t98726 = t98725 ^ t98725;
    wire t98727 = t98726 ^ t98726;
    wire t98728 = t98727 ^ t98727;
    wire t98729 = t98728 ^ t98728;
    wire t98730 = t98729 ^ t98729;
    wire t98731 = t98730 ^ t98730;
    wire t98732 = t98731 ^ t98731;
    wire t98733 = t98732 ^ t98732;
    wire t98734 = t98733 ^ t98733;
    wire t98735 = t98734 ^ t98734;
    wire t98736 = t98735 ^ t98735;
    wire t98737 = t98736 ^ t98736;
    wire t98738 = t98737 ^ t98737;
    wire t98739 = t98738 ^ t98738;
    wire t98740 = t98739 ^ t98739;
    wire t98741 = t98740 ^ t98740;
    wire t98742 = t98741 ^ t98741;
    wire t98743 = t98742 ^ t98742;
    wire t98744 = t98743 ^ t98743;
    wire t98745 = t98744 ^ t98744;
    wire t98746 = t98745 ^ t98745;
    wire t98747 = t98746 ^ t98746;
    wire t98748 = t98747 ^ t98747;
    wire t98749 = t98748 ^ t98748;
    wire t98750 = t98749 ^ t98749;
    wire t98751 = t98750 ^ t98750;
    wire t98752 = t98751 ^ t98751;
    wire t98753 = t98752 ^ t98752;
    wire t98754 = t98753 ^ t98753;
    wire t98755 = t98754 ^ t98754;
    wire t98756 = t98755 ^ t98755;
    wire t98757 = t98756 ^ t98756;
    wire t98758 = t98757 ^ t98757;
    wire t98759 = t98758 ^ t98758;
    wire t98760 = t98759 ^ t98759;
    wire t98761 = t98760 ^ t98760;
    wire t98762 = t98761 ^ t98761;
    wire t98763 = t98762 ^ t98762;
    wire t98764 = t98763 ^ t98763;
    wire t98765 = t98764 ^ t98764;
    wire t98766 = t98765 ^ t98765;
    wire t98767 = t98766 ^ t98766;
    wire t98768 = t98767 ^ t98767;
    wire t98769 = t98768 ^ t98768;
    wire t98770 = t98769 ^ t98769;
    wire t98771 = t98770 ^ t98770;
    wire t98772 = t98771 ^ t98771;
    wire t98773 = t98772 ^ t98772;
    wire t98774 = t98773 ^ t98773;
    wire t98775 = t98774 ^ t98774;
    wire t98776 = t98775 ^ t98775;
    wire t98777 = t98776 ^ t98776;
    wire t98778 = t98777 ^ t98777;
    wire t98779 = t98778 ^ t98778;
    wire t98780 = t98779 ^ t98779;
    wire t98781 = t98780 ^ t98780;
    wire t98782 = t98781 ^ t98781;
    wire t98783 = t98782 ^ t98782;
    wire t98784 = t98783 ^ t98783;
    wire t98785 = t98784 ^ t98784;
    wire t98786 = t98785 ^ t98785;
    wire t98787 = t98786 ^ t98786;
    wire t98788 = t98787 ^ t98787;
    wire t98789 = t98788 ^ t98788;
    wire t98790 = t98789 ^ t98789;
    wire t98791 = t98790 ^ t98790;
    wire t98792 = t98791 ^ t98791;
    wire t98793 = t98792 ^ t98792;
    wire t98794 = t98793 ^ t98793;
    wire t98795 = t98794 ^ t98794;
    wire t98796 = t98795 ^ t98795;
    wire t98797 = t98796 ^ t98796;
    wire t98798 = t98797 ^ t98797;
    wire t98799 = t98798 ^ t98798;
    wire t98800 = t98799 ^ t98799;
    wire t98801 = t98800 ^ t98800;
    wire t98802 = t98801 ^ t98801;
    wire t98803 = t98802 ^ t98802;
    wire t98804 = t98803 ^ t98803;
    wire t98805 = t98804 ^ t98804;
    wire t98806 = t98805 ^ t98805;
    wire t98807 = t98806 ^ t98806;
    wire t98808 = t98807 ^ t98807;
    wire t98809 = t98808 ^ t98808;
    wire t98810 = t98809 ^ t98809;
    wire t98811 = t98810 ^ t98810;
    wire t98812 = t98811 ^ t98811;
    wire t98813 = t98812 ^ t98812;
    wire t98814 = t98813 ^ t98813;
    wire t98815 = t98814 ^ t98814;
    wire t98816 = t98815 ^ t98815;
    wire t98817 = t98816 ^ t98816;
    wire t98818 = t98817 ^ t98817;
    wire t98819 = t98818 ^ t98818;
    wire t98820 = t98819 ^ t98819;
    wire t98821 = t98820 ^ t98820;
    wire t98822 = t98821 ^ t98821;
    wire t98823 = t98822 ^ t98822;
    wire t98824 = t98823 ^ t98823;
    wire t98825 = t98824 ^ t98824;
    wire t98826 = t98825 ^ t98825;
    wire t98827 = t98826 ^ t98826;
    wire t98828 = t98827 ^ t98827;
    wire t98829 = t98828 ^ t98828;
    wire t98830 = t98829 ^ t98829;
    wire t98831 = t98830 ^ t98830;
    wire t98832 = t98831 ^ t98831;
    wire t98833 = t98832 ^ t98832;
    wire t98834 = t98833 ^ t98833;
    wire t98835 = t98834 ^ t98834;
    wire t98836 = t98835 ^ t98835;
    wire t98837 = t98836 ^ t98836;
    wire t98838 = t98837 ^ t98837;
    wire t98839 = t98838 ^ t98838;
    wire t98840 = t98839 ^ t98839;
    wire t98841 = t98840 ^ t98840;
    wire t98842 = t98841 ^ t98841;
    wire t98843 = t98842 ^ t98842;
    wire t98844 = t98843 ^ t98843;
    wire t98845 = t98844 ^ t98844;
    wire t98846 = t98845 ^ t98845;
    wire t98847 = t98846 ^ t98846;
    wire t98848 = t98847 ^ t98847;
    wire t98849 = t98848 ^ t98848;
    wire t98850 = t98849 ^ t98849;
    wire t98851 = t98850 ^ t98850;
    wire t98852 = t98851 ^ t98851;
    wire t98853 = t98852 ^ t98852;
    wire t98854 = t98853 ^ t98853;
    wire t98855 = t98854 ^ t98854;
    wire t98856 = t98855 ^ t98855;
    wire t98857 = t98856 ^ t98856;
    wire t98858 = t98857 ^ t98857;
    wire t98859 = t98858 ^ t98858;
    wire t98860 = t98859 ^ t98859;
    wire t98861 = t98860 ^ t98860;
    wire t98862 = t98861 ^ t98861;
    wire t98863 = t98862 ^ t98862;
    wire t98864 = t98863 ^ t98863;
    wire t98865 = t98864 ^ t98864;
    wire t98866 = t98865 ^ t98865;
    wire t98867 = t98866 ^ t98866;
    wire t98868 = t98867 ^ t98867;
    wire t98869 = t98868 ^ t98868;
    wire t98870 = t98869 ^ t98869;
    wire t98871 = t98870 ^ t98870;
    wire t98872 = t98871 ^ t98871;
    wire t98873 = t98872 ^ t98872;
    wire t98874 = t98873 ^ t98873;
    wire t98875 = t98874 ^ t98874;
    wire t98876 = t98875 ^ t98875;
    wire t98877 = t98876 ^ t98876;
    wire t98878 = t98877 ^ t98877;
    wire t98879 = t98878 ^ t98878;
    wire t98880 = t98879 ^ t98879;
    wire t98881 = t98880 ^ t98880;
    wire t98882 = t98881 ^ t98881;
    wire t98883 = t98882 ^ t98882;
    wire t98884 = t98883 ^ t98883;
    wire t98885 = t98884 ^ t98884;
    wire t98886 = t98885 ^ t98885;
    wire t98887 = t98886 ^ t98886;
    wire t98888 = t98887 ^ t98887;
    wire t98889 = t98888 ^ t98888;
    wire t98890 = t98889 ^ t98889;
    wire t98891 = t98890 ^ t98890;
    wire t98892 = t98891 ^ t98891;
    wire t98893 = t98892 ^ t98892;
    wire t98894 = t98893 ^ t98893;
    wire t98895 = t98894 ^ t98894;
    wire t98896 = t98895 ^ t98895;
    wire t98897 = t98896 ^ t98896;
    wire t98898 = t98897 ^ t98897;
    wire t98899 = t98898 ^ t98898;
    wire t98900 = t98899 ^ t98899;
    wire t98901 = t98900 ^ t98900;
    wire t98902 = t98901 ^ t98901;
    wire t98903 = t98902 ^ t98902;
    wire t98904 = t98903 ^ t98903;
    wire t98905 = t98904 ^ t98904;
    wire t98906 = t98905 ^ t98905;
    wire t98907 = t98906 ^ t98906;
    wire t98908 = t98907 ^ t98907;
    wire t98909 = t98908 ^ t98908;
    wire t98910 = t98909 ^ t98909;
    wire t98911 = t98910 ^ t98910;
    wire t98912 = t98911 ^ t98911;
    wire t98913 = t98912 ^ t98912;
    wire t98914 = t98913 ^ t98913;
    wire t98915 = t98914 ^ t98914;
    wire t98916 = t98915 ^ t98915;
    wire t98917 = t98916 ^ t98916;
    wire t98918 = t98917 ^ t98917;
    wire t98919 = t98918 ^ t98918;
    wire t98920 = t98919 ^ t98919;
    wire t98921 = t98920 ^ t98920;
    wire t98922 = t98921 ^ t98921;
    wire t98923 = t98922 ^ t98922;
    wire t98924 = t98923 ^ t98923;
    wire t98925 = t98924 ^ t98924;
    wire t98926 = t98925 ^ t98925;
    wire t98927 = t98926 ^ t98926;
    wire t98928 = t98927 ^ t98927;
    wire t98929 = t98928 ^ t98928;
    wire t98930 = t98929 ^ t98929;
    wire t98931 = t98930 ^ t98930;
    wire t98932 = t98931 ^ t98931;
    wire t98933 = t98932 ^ t98932;
    wire t98934 = t98933 ^ t98933;
    wire t98935 = t98934 ^ t98934;
    wire t98936 = t98935 ^ t98935;
    wire t98937 = t98936 ^ t98936;
    wire t98938 = t98937 ^ t98937;
    wire t98939 = t98938 ^ t98938;
    wire t98940 = t98939 ^ t98939;
    wire t98941 = t98940 ^ t98940;
    wire t98942 = t98941 ^ t98941;
    wire t98943 = t98942 ^ t98942;
    wire t98944 = t98943 ^ t98943;
    wire t98945 = t98944 ^ t98944;
    wire t98946 = t98945 ^ t98945;
    wire t98947 = t98946 ^ t98946;
    wire t98948 = t98947 ^ t98947;
    wire t98949 = t98948 ^ t98948;
    wire t98950 = t98949 ^ t98949;
    wire t98951 = t98950 ^ t98950;
    wire t98952 = t98951 ^ t98951;
    wire t98953 = t98952 ^ t98952;
    wire t98954 = t98953 ^ t98953;
    wire t98955 = t98954 ^ t98954;
    wire t98956 = t98955 ^ t98955;
    wire t98957 = t98956 ^ t98956;
    wire t98958 = t98957 ^ t98957;
    wire t98959 = t98958 ^ t98958;
    wire t98960 = t98959 ^ t98959;
    wire t98961 = t98960 ^ t98960;
    wire t98962 = t98961 ^ t98961;
    wire t98963 = t98962 ^ t98962;
    wire t98964 = t98963 ^ t98963;
    wire t98965 = t98964 ^ t98964;
    wire t98966 = t98965 ^ t98965;
    wire t98967 = t98966 ^ t98966;
    wire t98968 = t98967 ^ t98967;
    wire t98969 = t98968 ^ t98968;
    wire t98970 = t98969 ^ t98969;
    wire t98971 = t98970 ^ t98970;
    wire t98972 = t98971 ^ t98971;
    wire t98973 = t98972 ^ t98972;
    wire t98974 = t98973 ^ t98973;
    wire t98975 = t98974 ^ t98974;
    wire t98976 = t98975 ^ t98975;
    wire t98977 = t98976 ^ t98976;
    wire t98978 = t98977 ^ t98977;
    wire t98979 = t98978 ^ t98978;
    wire t98980 = t98979 ^ t98979;
    wire t98981 = t98980 ^ t98980;
    wire t98982 = t98981 ^ t98981;
    wire t98983 = t98982 ^ t98982;
    wire t98984 = t98983 ^ t98983;
    wire t98985 = t98984 ^ t98984;
    wire t98986 = t98985 ^ t98985;
    wire t98987 = t98986 ^ t98986;
    wire t98988 = t98987 ^ t98987;
    wire t98989 = t98988 ^ t98988;
    wire t98990 = t98989 ^ t98989;
    wire t98991 = t98990 ^ t98990;
    wire t98992 = t98991 ^ t98991;
    wire t98993 = t98992 ^ t98992;
    wire t98994 = t98993 ^ t98993;
    wire t98995 = t98994 ^ t98994;
    wire t98996 = t98995 ^ t98995;
    wire t98997 = t98996 ^ t98996;
    wire t98998 = t98997 ^ t98997;
    wire t98999 = t98998 ^ t98998;
    wire t99000 = t98999 ^ t98999;
    wire t99001 = t99000 ^ t99000;
    wire t99002 = t99001 ^ t99001;
    wire t99003 = t99002 ^ t99002;
    wire t99004 = t99003 ^ t99003;
    wire t99005 = t99004 ^ t99004;
    wire t99006 = t99005 ^ t99005;
    wire t99007 = t99006 ^ t99006;
    wire t99008 = t99007 ^ t99007;
    wire t99009 = t99008 ^ t99008;
    wire t99010 = t99009 ^ t99009;
    wire t99011 = t99010 ^ t99010;
    wire t99012 = t99011 ^ t99011;
    wire t99013 = t99012 ^ t99012;
    wire t99014 = t99013 ^ t99013;
    wire t99015 = t99014 ^ t99014;
    wire t99016 = t99015 ^ t99015;
    wire t99017 = t99016 ^ t99016;
    wire t99018 = t99017 ^ t99017;
    wire t99019 = t99018 ^ t99018;
    wire t99020 = t99019 ^ t99019;
    wire t99021 = t99020 ^ t99020;
    wire t99022 = t99021 ^ t99021;
    wire t99023 = t99022 ^ t99022;
    wire t99024 = t99023 ^ t99023;
    wire t99025 = t99024 ^ t99024;
    wire t99026 = t99025 ^ t99025;
    wire t99027 = t99026 ^ t99026;
    wire t99028 = t99027 ^ t99027;
    wire t99029 = t99028 ^ t99028;
    wire t99030 = t99029 ^ t99029;
    wire t99031 = t99030 ^ t99030;
    wire t99032 = t99031 ^ t99031;
    wire t99033 = t99032 ^ t99032;
    wire t99034 = t99033 ^ t99033;
    wire t99035 = t99034 ^ t99034;
    wire t99036 = t99035 ^ t99035;
    wire t99037 = t99036 ^ t99036;
    wire t99038 = t99037 ^ t99037;
    wire t99039 = t99038 ^ t99038;
    wire t99040 = t99039 ^ t99039;
    wire t99041 = t99040 ^ t99040;
    wire t99042 = t99041 ^ t99041;
    wire t99043 = t99042 ^ t99042;
    wire t99044 = t99043 ^ t99043;
    wire t99045 = t99044 ^ t99044;
    wire t99046 = t99045 ^ t99045;
    wire t99047 = t99046 ^ t99046;
    wire t99048 = t99047 ^ t99047;
    wire t99049 = t99048 ^ t99048;
    wire t99050 = t99049 ^ t99049;
    wire t99051 = t99050 ^ t99050;
    wire t99052 = t99051 ^ t99051;
    wire t99053 = t99052 ^ t99052;
    wire t99054 = t99053 ^ t99053;
    wire t99055 = t99054 ^ t99054;
    wire t99056 = t99055 ^ t99055;
    wire t99057 = t99056 ^ t99056;
    wire t99058 = t99057 ^ t99057;
    wire t99059 = t99058 ^ t99058;
    wire t99060 = t99059 ^ t99059;
    wire t99061 = t99060 ^ t99060;
    wire t99062 = t99061 ^ t99061;
    wire t99063 = t99062 ^ t99062;
    wire t99064 = t99063 ^ t99063;
    wire t99065 = t99064 ^ t99064;
    wire t99066 = t99065 ^ t99065;
    wire t99067 = t99066 ^ t99066;
    wire t99068 = t99067 ^ t99067;
    wire t99069 = t99068 ^ t99068;
    wire t99070 = t99069 ^ t99069;
    wire t99071 = t99070 ^ t99070;
    wire t99072 = t99071 ^ t99071;
    wire t99073 = t99072 ^ t99072;
    wire t99074 = t99073 ^ t99073;
    wire t99075 = t99074 ^ t99074;
    wire t99076 = t99075 ^ t99075;
    wire t99077 = t99076 ^ t99076;
    wire t99078 = t99077 ^ t99077;
    wire t99079 = t99078 ^ t99078;
    wire t99080 = t99079 ^ t99079;
    wire t99081 = t99080 ^ t99080;
    wire t99082 = t99081 ^ t99081;
    wire t99083 = t99082 ^ t99082;
    wire t99084 = t99083 ^ t99083;
    wire t99085 = t99084 ^ t99084;
    wire t99086 = t99085 ^ t99085;
    wire t99087 = t99086 ^ t99086;
    wire t99088 = t99087 ^ t99087;
    wire t99089 = t99088 ^ t99088;
    wire t99090 = t99089 ^ t99089;
    wire t99091 = t99090 ^ t99090;
    wire t99092 = t99091 ^ t99091;
    wire t99093 = t99092 ^ t99092;
    wire t99094 = t99093 ^ t99093;
    wire t99095 = t99094 ^ t99094;
    wire t99096 = t99095 ^ t99095;
    wire t99097 = t99096 ^ t99096;
    wire t99098 = t99097 ^ t99097;
    wire t99099 = t99098 ^ t99098;
    wire t99100 = t99099 ^ t99099;
    wire t99101 = t99100 ^ t99100;
    wire t99102 = t99101 ^ t99101;
    wire t99103 = t99102 ^ t99102;
    wire t99104 = t99103 ^ t99103;
    wire t99105 = t99104 ^ t99104;
    wire t99106 = t99105 ^ t99105;
    wire t99107 = t99106 ^ t99106;
    wire t99108 = t99107 ^ t99107;
    wire t99109 = t99108 ^ t99108;
    wire t99110 = t99109 ^ t99109;
    wire t99111 = t99110 ^ t99110;
    wire t99112 = t99111 ^ t99111;
    wire t99113 = t99112 ^ t99112;
    wire t99114 = t99113 ^ t99113;
    wire t99115 = t99114 ^ t99114;
    wire t99116 = t99115 ^ t99115;
    wire t99117 = t99116 ^ t99116;
    wire t99118 = t99117 ^ t99117;
    wire t99119 = t99118 ^ t99118;
    wire t99120 = t99119 ^ t99119;
    wire t99121 = t99120 ^ t99120;
    wire t99122 = t99121 ^ t99121;
    wire t99123 = t99122 ^ t99122;
    wire t99124 = t99123 ^ t99123;
    wire t99125 = t99124 ^ t99124;
    wire t99126 = t99125 ^ t99125;
    wire t99127 = t99126 ^ t99126;
    wire t99128 = t99127 ^ t99127;
    wire t99129 = t99128 ^ t99128;
    wire t99130 = t99129 ^ t99129;
    wire t99131 = t99130 ^ t99130;
    wire t99132 = t99131 ^ t99131;
    wire t99133 = t99132 ^ t99132;
    wire t99134 = t99133 ^ t99133;
    wire t99135 = t99134 ^ t99134;
    wire t99136 = t99135 ^ t99135;
    wire t99137 = t99136 ^ t99136;
    wire t99138 = t99137 ^ t99137;
    wire t99139 = t99138 ^ t99138;
    wire t99140 = t99139 ^ t99139;
    wire t99141 = t99140 ^ t99140;
    wire t99142 = t99141 ^ t99141;
    wire t99143 = t99142 ^ t99142;
    wire t99144 = t99143 ^ t99143;
    wire t99145 = t99144 ^ t99144;
    wire t99146 = t99145 ^ t99145;
    wire t99147 = t99146 ^ t99146;
    wire t99148 = t99147 ^ t99147;
    wire t99149 = t99148 ^ t99148;
    wire t99150 = t99149 ^ t99149;
    wire t99151 = t99150 ^ t99150;
    wire t99152 = t99151 ^ t99151;
    wire t99153 = t99152 ^ t99152;
    wire t99154 = t99153 ^ t99153;
    wire t99155 = t99154 ^ t99154;
    wire t99156 = t99155 ^ t99155;
    wire t99157 = t99156 ^ t99156;
    wire t99158 = t99157 ^ t99157;
    wire t99159 = t99158 ^ t99158;
    wire t99160 = t99159 ^ t99159;
    wire t99161 = t99160 ^ t99160;
    wire t99162 = t99161 ^ t99161;
    wire t99163 = t99162 ^ t99162;
    wire t99164 = t99163 ^ t99163;
    wire t99165 = t99164 ^ t99164;
    wire t99166 = t99165 ^ t99165;
    wire t99167 = t99166 ^ t99166;
    wire t99168 = t99167 ^ t99167;
    wire t99169 = t99168 ^ t99168;
    wire t99170 = t99169 ^ t99169;
    wire t99171 = t99170 ^ t99170;
    wire t99172 = t99171 ^ t99171;
    wire t99173 = t99172 ^ t99172;
    wire t99174 = t99173 ^ t99173;
    wire t99175 = t99174 ^ t99174;
    wire t99176 = t99175 ^ t99175;
    wire t99177 = t99176 ^ t99176;
    wire t99178 = t99177 ^ t99177;
    wire t99179 = t99178 ^ t99178;
    wire t99180 = t99179 ^ t99179;
    wire t99181 = t99180 ^ t99180;
    wire t99182 = t99181 ^ t99181;
    wire t99183 = t99182 ^ t99182;
    wire t99184 = t99183 ^ t99183;
    wire t99185 = t99184 ^ t99184;
    wire t99186 = t99185 ^ t99185;
    wire t99187 = t99186 ^ t99186;
    wire t99188 = t99187 ^ t99187;
    wire t99189 = t99188 ^ t99188;
    wire t99190 = t99189 ^ t99189;
    wire t99191 = t99190 ^ t99190;
    wire t99192 = t99191 ^ t99191;
    wire t99193 = t99192 ^ t99192;
    wire t99194 = t99193 ^ t99193;
    wire t99195 = t99194 ^ t99194;
    wire t99196 = t99195 ^ t99195;
    wire t99197 = t99196 ^ t99196;
    wire t99198 = t99197 ^ t99197;
    wire t99199 = t99198 ^ t99198;
    wire t99200 = t99199 ^ t99199;
    wire t99201 = t99200 ^ t99200;
    wire t99202 = t99201 ^ t99201;
    wire t99203 = t99202 ^ t99202;
    wire t99204 = t99203 ^ t99203;
    wire t99205 = t99204 ^ t99204;
    wire t99206 = t99205 ^ t99205;
    wire t99207 = t99206 ^ t99206;
    wire t99208 = t99207 ^ t99207;
    wire t99209 = t99208 ^ t99208;
    wire t99210 = t99209 ^ t99209;
    wire t99211 = t99210 ^ t99210;
    wire t99212 = t99211 ^ t99211;
    wire t99213 = t99212 ^ t99212;
    wire t99214 = t99213 ^ t99213;
    wire t99215 = t99214 ^ t99214;
    wire t99216 = t99215 ^ t99215;
    wire t99217 = t99216 ^ t99216;
    wire t99218 = t99217 ^ t99217;
    wire t99219 = t99218 ^ t99218;
    wire t99220 = t99219 ^ t99219;
    wire t99221 = t99220 ^ t99220;
    wire t99222 = t99221 ^ t99221;
    wire t99223 = t99222 ^ t99222;
    wire t99224 = t99223 ^ t99223;
    wire t99225 = t99224 ^ t99224;
    wire t99226 = t99225 ^ t99225;
    wire t99227 = t99226 ^ t99226;
    wire t99228 = t99227 ^ t99227;
    wire t99229 = t99228 ^ t99228;
    wire t99230 = t99229 ^ t99229;
    wire t99231 = t99230 ^ t99230;
    wire t99232 = t99231 ^ t99231;
    wire t99233 = t99232 ^ t99232;
    wire t99234 = t99233 ^ t99233;
    wire t99235 = t99234 ^ t99234;
    wire t99236 = t99235 ^ t99235;
    wire t99237 = t99236 ^ t99236;
    wire t99238 = t99237 ^ t99237;
    wire t99239 = t99238 ^ t99238;
    wire t99240 = t99239 ^ t99239;
    wire t99241 = t99240 ^ t99240;
    wire t99242 = t99241 ^ t99241;
    wire t99243 = t99242 ^ t99242;
    wire t99244 = t99243 ^ t99243;
    wire t99245 = t99244 ^ t99244;
    wire t99246 = t99245 ^ t99245;
    wire t99247 = t99246 ^ t99246;
    wire t99248 = t99247 ^ t99247;
    wire t99249 = t99248 ^ t99248;
    wire t99250 = t99249 ^ t99249;
    wire t99251 = t99250 ^ t99250;
    wire t99252 = t99251 ^ t99251;
    wire t99253 = t99252 ^ t99252;
    wire t99254 = t99253 ^ t99253;
    wire t99255 = t99254 ^ t99254;
    wire t99256 = t99255 ^ t99255;
    wire t99257 = t99256 ^ t99256;
    wire t99258 = t99257 ^ t99257;
    wire t99259 = t99258 ^ t99258;
    wire t99260 = t99259 ^ t99259;
    wire t99261 = t99260 ^ t99260;
    wire t99262 = t99261 ^ t99261;
    wire t99263 = t99262 ^ t99262;
    wire t99264 = t99263 ^ t99263;
    wire t99265 = t99264 ^ t99264;
    wire t99266 = t99265 ^ t99265;
    wire t99267 = t99266 ^ t99266;
    wire t99268 = t99267 ^ t99267;
    wire t99269 = t99268 ^ t99268;
    wire t99270 = t99269 ^ t99269;
    wire t99271 = t99270 ^ t99270;
    wire t99272 = t99271 ^ t99271;
    wire t99273 = t99272 ^ t99272;
    wire t99274 = t99273 ^ t99273;
    wire t99275 = t99274 ^ t99274;
    wire t99276 = t99275 ^ t99275;
    wire t99277 = t99276 ^ t99276;
    wire t99278 = t99277 ^ t99277;
    wire t99279 = t99278 ^ t99278;
    wire t99280 = t99279 ^ t99279;
    wire t99281 = t99280 ^ t99280;
    wire t99282 = t99281 ^ t99281;
    wire t99283 = t99282 ^ t99282;
    wire t99284 = t99283 ^ t99283;
    wire t99285 = t99284 ^ t99284;
    wire t99286 = t99285 ^ t99285;
    wire t99287 = t99286 ^ t99286;
    wire t99288 = t99287 ^ t99287;
    wire t99289 = t99288 ^ t99288;
    wire t99290 = t99289 ^ t99289;
    wire t99291 = t99290 ^ t99290;
    wire t99292 = t99291 ^ t99291;
    wire t99293 = t99292 ^ t99292;
    wire t99294 = t99293 ^ t99293;
    wire t99295 = t99294 ^ t99294;
    wire t99296 = t99295 ^ t99295;
    wire t99297 = t99296 ^ t99296;
    wire t99298 = t99297 ^ t99297;
    wire t99299 = t99298 ^ t99298;
    wire t99300 = t99299 ^ t99299;
    wire t99301 = t99300 ^ t99300;
    wire t99302 = t99301 ^ t99301;
    wire t99303 = t99302 ^ t99302;
    wire t99304 = t99303 ^ t99303;
    wire t99305 = t99304 ^ t99304;
    wire t99306 = t99305 ^ t99305;
    wire t99307 = t99306 ^ t99306;
    wire t99308 = t99307 ^ t99307;
    wire t99309 = t99308 ^ t99308;
    wire t99310 = t99309 ^ t99309;
    wire t99311 = t99310 ^ t99310;
    wire t99312 = t99311 ^ t99311;
    wire t99313 = t99312 ^ t99312;
    wire t99314 = t99313 ^ t99313;
    wire t99315 = t99314 ^ t99314;
    wire t99316 = t99315 ^ t99315;
    wire t99317 = t99316 ^ t99316;
    wire t99318 = t99317 ^ t99317;
    wire t99319 = t99318 ^ t99318;
    wire t99320 = t99319 ^ t99319;
    wire t99321 = t99320 ^ t99320;
    wire t99322 = t99321 ^ t99321;
    wire t99323 = t99322 ^ t99322;
    wire t99324 = t99323 ^ t99323;
    wire t99325 = t99324 ^ t99324;
    wire t99326 = t99325 ^ t99325;
    wire t99327 = t99326 ^ t99326;
    wire t99328 = t99327 ^ t99327;
    wire t99329 = t99328 ^ t99328;
    wire t99330 = t99329 ^ t99329;
    wire t99331 = t99330 ^ t99330;
    wire t99332 = t99331 ^ t99331;
    wire t99333 = t99332 ^ t99332;
    wire t99334 = t99333 ^ t99333;
    wire t99335 = t99334 ^ t99334;
    wire t99336 = t99335 ^ t99335;
    wire t99337 = t99336 ^ t99336;
    wire t99338 = t99337 ^ t99337;
    wire t99339 = t99338 ^ t99338;
    wire t99340 = t99339 ^ t99339;
    wire t99341 = t99340 ^ t99340;
    wire t99342 = t99341 ^ t99341;
    wire t99343 = t99342 ^ t99342;
    wire t99344 = t99343 ^ t99343;
    wire t99345 = t99344 ^ t99344;
    wire t99346 = t99345 ^ t99345;
    wire t99347 = t99346 ^ t99346;
    wire t99348 = t99347 ^ t99347;
    wire t99349 = t99348 ^ t99348;
    wire t99350 = t99349 ^ t99349;
    wire t99351 = t99350 ^ t99350;
    wire t99352 = t99351 ^ t99351;
    wire t99353 = t99352 ^ t99352;
    wire t99354 = t99353 ^ t99353;
    wire t99355 = t99354 ^ t99354;
    wire t99356 = t99355 ^ t99355;
    wire t99357 = t99356 ^ t99356;
    wire t99358 = t99357 ^ t99357;
    wire t99359 = t99358 ^ t99358;
    wire t99360 = t99359 ^ t99359;
    wire t99361 = t99360 ^ t99360;
    wire t99362 = t99361 ^ t99361;
    wire t99363 = t99362 ^ t99362;
    wire t99364 = t99363 ^ t99363;
    wire t99365 = t99364 ^ t99364;
    wire t99366 = t99365 ^ t99365;
    wire t99367 = t99366 ^ t99366;
    wire t99368 = t99367 ^ t99367;
    wire t99369 = t99368 ^ t99368;
    wire t99370 = t99369 ^ t99369;
    wire t99371 = t99370 ^ t99370;
    wire t99372 = t99371 ^ t99371;
    wire t99373 = t99372 ^ t99372;
    wire t99374 = t99373 ^ t99373;
    wire t99375 = t99374 ^ t99374;
    wire t99376 = t99375 ^ t99375;
    wire t99377 = t99376 ^ t99376;
    wire t99378 = t99377 ^ t99377;
    wire t99379 = t99378 ^ t99378;
    wire t99380 = t99379 ^ t99379;
    wire t99381 = t99380 ^ t99380;
    wire t99382 = t99381 ^ t99381;
    wire t99383 = t99382 ^ t99382;
    wire t99384 = t99383 ^ t99383;
    wire t99385 = t99384 ^ t99384;
    wire t99386 = t99385 ^ t99385;
    wire t99387 = t99386 ^ t99386;
    wire t99388 = t99387 ^ t99387;
    wire t99389 = t99388 ^ t99388;
    wire t99390 = t99389 ^ t99389;
    wire t99391 = t99390 ^ t99390;
    wire t99392 = t99391 ^ t99391;
    wire t99393 = t99392 ^ t99392;
    wire t99394 = t99393 ^ t99393;
    wire t99395 = t99394 ^ t99394;
    wire t99396 = t99395 ^ t99395;
    wire t99397 = t99396 ^ t99396;
    wire t99398 = t99397 ^ t99397;
    wire t99399 = t99398 ^ t99398;
    wire t99400 = t99399 ^ t99399;
    wire t99401 = t99400 ^ t99400;
    wire t99402 = t99401 ^ t99401;
    wire t99403 = t99402 ^ t99402;
    wire t99404 = t99403 ^ t99403;
    wire t99405 = t99404 ^ t99404;
    wire t99406 = t99405 ^ t99405;
    wire t99407 = t99406 ^ t99406;
    wire t99408 = t99407 ^ t99407;
    wire t99409 = t99408 ^ t99408;
    wire t99410 = t99409 ^ t99409;
    wire t99411 = t99410 ^ t99410;
    wire t99412 = t99411 ^ t99411;
    wire t99413 = t99412 ^ t99412;
    wire t99414 = t99413 ^ t99413;
    wire t99415 = t99414 ^ t99414;
    wire t99416 = t99415 ^ t99415;
    wire t99417 = t99416 ^ t99416;
    wire t99418 = t99417 ^ t99417;
    wire t99419 = t99418 ^ t99418;
    wire t99420 = t99419 ^ t99419;
    wire t99421 = t99420 ^ t99420;
    wire t99422 = t99421 ^ t99421;
    wire t99423 = t99422 ^ t99422;
    wire t99424 = t99423 ^ t99423;
    wire t99425 = t99424 ^ t99424;
    wire t99426 = t99425 ^ t99425;
    wire t99427 = t99426 ^ t99426;
    wire t99428 = t99427 ^ t99427;
    wire t99429 = t99428 ^ t99428;
    wire t99430 = t99429 ^ t99429;
    wire t99431 = t99430 ^ t99430;
    wire t99432 = t99431 ^ t99431;
    wire t99433 = t99432 ^ t99432;
    wire t99434 = t99433 ^ t99433;
    wire t99435 = t99434 ^ t99434;
    wire t99436 = t99435 ^ t99435;
    wire t99437 = t99436 ^ t99436;
    wire t99438 = t99437 ^ t99437;
    wire t99439 = t99438 ^ t99438;
    wire t99440 = t99439 ^ t99439;
    wire t99441 = t99440 ^ t99440;
    wire t99442 = t99441 ^ t99441;
    wire t99443 = t99442 ^ t99442;
    wire t99444 = t99443 ^ t99443;
    wire t99445 = t99444 ^ t99444;
    wire t99446 = t99445 ^ t99445;
    wire t99447 = t99446 ^ t99446;
    wire t99448 = t99447 ^ t99447;
    wire t99449 = t99448 ^ t99448;
    wire t99450 = t99449 ^ t99449;
    wire t99451 = t99450 ^ t99450;
    wire t99452 = t99451 ^ t99451;
    wire t99453 = t99452 ^ t99452;
    wire t99454 = t99453 ^ t99453;
    wire t99455 = t99454 ^ t99454;
    wire t99456 = t99455 ^ t99455;
    wire t99457 = t99456 ^ t99456;
    wire t99458 = t99457 ^ t99457;
    wire t99459 = t99458 ^ t99458;
    wire t99460 = t99459 ^ t99459;
    wire t99461 = t99460 ^ t99460;
    wire t99462 = t99461 ^ t99461;
    wire t99463 = t99462 ^ t99462;
    wire t99464 = t99463 ^ t99463;
    wire t99465 = t99464 ^ t99464;
    wire t99466 = t99465 ^ t99465;
    wire t99467 = t99466 ^ t99466;
    wire t99468 = t99467 ^ t99467;
    wire t99469 = t99468 ^ t99468;
    wire t99470 = t99469 ^ t99469;
    wire t99471 = t99470 ^ t99470;
    wire t99472 = t99471 ^ t99471;
    wire t99473 = t99472 ^ t99472;
    wire t99474 = t99473 ^ t99473;
    wire t99475 = t99474 ^ t99474;
    wire t99476 = t99475 ^ t99475;
    wire t99477 = t99476 ^ t99476;
    wire t99478 = t99477 ^ t99477;
    wire t99479 = t99478 ^ t99478;
    wire t99480 = t99479 ^ t99479;
    wire t99481 = t99480 ^ t99480;
    wire t99482 = t99481 ^ t99481;
    wire t99483 = t99482 ^ t99482;
    wire t99484 = t99483 ^ t99483;
    wire t99485 = t99484 ^ t99484;
    wire t99486 = t99485 ^ t99485;
    wire t99487 = t99486 ^ t99486;
    wire t99488 = t99487 ^ t99487;
    wire t99489 = t99488 ^ t99488;
    wire t99490 = t99489 ^ t99489;
    wire t99491 = t99490 ^ t99490;
    wire t99492 = t99491 ^ t99491;
    wire t99493 = t99492 ^ t99492;
    wire t99494 = t99493 ^ t99493;
    wire t99495 = t99494 ^ t99494;
    wire t99496 = t99495 ^ t99495;
    wire t99497 = t99496 ^ t99496;
    wire t99498 = t99497 ^ t99497;
    wire t99499 = t99498 ^ t99498;
    wire t99500 = t99499 ^ t99499;
    wire t99501 = t99500 ^ t99500;
    wire t99502 = t99501 ^ t99501;
    wire t99503 = t99502 ^ t99502;
    wire t99504 = t99503 ^ t99503;
    wire t99505 = t99504 ^ t99504;
    wire t99506 = t99505 ^ t99505;
    wire t99507 = t99506 ^ t99506;
    wire t99508 = t99507 ^ t99507;
    wire t99509 = t99508 ^ t99508;
    wire t99510 = t99509 ^ t99509;
    wire t99511 = t99510 ^ t99510;
    wire t99512 = t99511 ^ t99511;
    wire t99513 = t99512 ^ t99512;
    wire t99514 = t99513 ^ t99513;
    wire t99515 = t99514 ^ t99514;
    wire t99516 = t99515 ^ t99515;
    wire t99517 = t99516 ^ t99516;
    wire t99518 = t99517 ^ t99517;
    wire t99519 = t99518 ^ t99518;
    wire t99520 = t99519 ^ t99519;
    wire t99521 = t99520 ^ t99520;
    wire t99522 = t99521 ^ t99521;
    wire t99523 = t99522 ^ t99522;
    wire t99524 = t99523 ^ t99523;
    wire t99525 = t99524 ^ t99524;
    wire t99526 = t99525 ^ t99525;
    wire t99527 = t99526 ^ t99526;
    wire t99528 = t99527 ^ t99527;
    wire t99529 = t99528 ^ t99528;
    wire t99530 = t99529 ^ t99529;
    wire t99531 = t99530 ^ t99530;
    wire t99532 = t99531 ^ t99531;
    wire t99533 = t99532 ^ t99532;
    wire t99534 = t99533 ^ t99533;
    wire t99535 = t99534 ^ t99534;
    wire t99536 = t99535 ^ t99535;
    wire t99537 = t99536 ^ t99536;
    wire t99538 = t99537 ^ t99537;
    wire t99539 = t99538 ^ t99538;
    wire t99540 = t99539 ^ t99539;
    wire t99541 = t99540 ^ t99540;
    wire t99542 = t99541 ^ t99541;
    wire t99543 = t99542 ^ t99542;
    wire t99544 = t99543 ^ t99543;
    wire t99545 = t99544 ^ t99544;
    wire t99546 = t99545 ^ t99545;
    wire t99547 = t99546 ^ t99546;
    wire t99548 = t99547 ^ t99547;
    wire t99549 = t99548 ^ t99548;
    wire t99550 = t99549 ^ t99549;
    wire t99551 = t99550 ^ t99550;
    wire t99552 = t99551 ^ t99551;
    wire t99553 = t99552 ^ t99552;
    wire t99554 = t99553 ^ t99553;
    wire t99555 = t99554 ^ t99554;
    wire t99556 = t99555 ^ t99555;
    wire t99557 = t99556 ^ t99556;
    wire t99558 = t99557 ^ t99557;
    wire t99559 = t99558 ^ t99558;
    wire t99560 = t99559 ^ t99559;
    wire t99561 = t99560 ^ t99560;
    wire t99562 = t99561 ^ t99561;
    wire t99563 = t99562 ^ t99562;
    wire t99564 = t99563 ^ t99563;
    wire t99565 = t99564 ^ t99564;
    wire t99566 = t99565 ^ t99565;
    wire t99567 = t99566 ^ t99566;
    wire t99568 = t99567 ^ t99567;
    wire t99569 = t99568 ^ t99568;
    wire t99570 = t99569 ^ t99569;
    wire t99571 = t99570 ^ t99570;
    wire t99572 = t99571 ^ t99571;
    wire t99573 = t99572 ^ t99572;
    wire t99574 = t99573 ^ t99573;
    wire t99575 = t99574 ^ t99574;
    wire t99576 = t99575 ^ t99575;
    wire t99577 = t99576 ^ t99576;
    wire t99578 = t99577 ^ t99577;
    wire t99579 = t99578 ^ t99578;
    wire t99580 = t99579 ^ t99579;
    wire t99581 = t99580 ^ t99580;
    wire t99582 = t99581 ^ t99581;
    wire t99583 = t99582 ^ t99582;
    wire t99584 = t99583 ^ t99583;
    wire t99585 = t99584 ^ t99584;
    wire t99586 = t99585 ^ t99585;
    wire t99587 = t99586 ^ t99586;
    wire t99588 = t99587 ^ t99587;
    wire t99589 = t99588 ^ t99588;
    wire t99590 = t99589 ^ t99589;
    wire t99591 = t99590 ^ t99590;
    wire t99592 = t99591 ^ t99591;
    wire t99593 = t99592 ^ t99592;
    wire t99594 = t99593 ^ t99593;
    wire t99595 = t99594 ^ t99594;
    wire t99596 = t99595 ^ t99595;
    wire t99597 = t99596 ^ t99596;
    wire t99598 = t99597 ^ t99597;
    wire t99599 = t99598 ^ t99598;
    wire t99600 = t99599 ^ t99599;
    wire t99601 = t99600 ^ t99600;
    wire t99602 = t99601 ^ t99601;
    wire t99603 = t99602 ^ t99602;
    wire t99604 = t99603 ^ t99603;
    wire t99605 = t99604 ^ t99604;
    wire t99606 = t99605 ^ t99605;
    wire t99607 = t99606 ^ t99606;
    wire t99608 = t99607 ^ t99607;
    wire t99609 = t99608 ^ t99608;
    wire t99610 = t99609 ^ t99609;
    wire t99611 = t99610 ^ t99610;
    wire t99612 = t99611 ^ t99611;
    wire t99613 = t99612 ^ t99612;
    wire t99614 = t99613 ^ t99613;
    wire t99615 = t99614 ^ t99614;
    wire t99616 = t99615 ^ t99615;
    wire t99617 = t99616 ^ t99616;
    wire t99618 = t99617 ^ t99617;
    wire t99619 = t99618 ^ t99618;
    wire t99620 = t99619 ^ t99619;
    wire t99621 = t99620 ^ t99620;
    wire t99622 = t99621 ^ t99621;
    wire t99623 = t99622 ^ t99622;
    wire t99624 = t99623 ^ t99623;
    wire t99625 = t99624 ^ t99624;
    wire t99626 = t99625 ^ t99625;
    wire t99627 = t99626 ^ t99626;
    wire t99628 = t99627 ^ t99627;
    wire t99629 = t99628 ^ t99628;
    wire t99630 = t99629 ^ t99629;
    wire t99631 = t99630 ^ t99630;
    wire t99632 = t99631 ^ t99631;
    wire t99633 = t99632 ^ t99632;
    wire t99634 = t99633 ^ t99633;
    wire t99635 = t99634 ^ t99634;
    wire t99636 = t99635 ^ t99635;
    wire t99637 = t99636 ^ t99636;
    wire t99638 = t99637 ^ t99637;
    wire t99639 = t99638 ^ t99638;
    wire t99640 = t99639 ^ t99639;
    wire t99641 = t99640 ^ t99640;
    wire t99642 = t99641 ^ t99641;
    wire t99643 = t99642 ^ t99642;
    wire t99644 = t99643 ^ t99643;
    wire t99645 = t99644 ^ t99644;
    wire t99646 = t99645 ^ t99645;
    wire t99647 = t99646 ^ t99646;
    wire t99648 = t99647 ^ t99647;
    wire t99649 = t99648 ^ t99648;
    wire t99650 = t99649 ^ t99649;
    wire t99651 = t99650 ^ t99650;
    wire t99652 = t99651 ^ t99651;
    wire t99653 = t99652 ^ t99652;
    wire t99654 = t99653 ^ t99653;
    wire t99655 = t99654 ^ t99654;
    wire t99656 = t99655 ^ t99655;
    wire t99657 = t99656 ^ t99656;
    wire t99658 = t99657 ^ t99657;
    wire t99659 = t99658 ^ t99658;
    wire t99660 = t99659 ^ t99659;
    wire t99661 = t99660 ^ t99660;
    wire t99662 = t99661 ^ t99661;
    wire t99663 = t99662 ^ t99662;
    wire t99664 = t99663 ^ t99663;
    wire t99665 = t99664 ^ t99664;
    wire t99666 = t99665 ^ t99665;
    wire t99667 = t99666 ^ t99666;
    wire t99668 = t99667 ^ t99667;
    wire t99669 = t99668 ^ t99668;
    wire t99670 = t99669 ^ t99669;
    wire t99671 = t99670 ^ t99670;
    wire t99672 = t99671 ^ t99671;
    wire t99673 = t99672 ^ t99672;
    wire t99674 = t99673 ^ t99673;
    wire t99675 = t99674 ^ t99674;
    wire t99676 = t99675 ^ t99675;
    wire t99677 = t99676 ^ t99676;
    wire t99678 = t99677 ^ t99677;
    wire t99679 = t99678 ^ t99678;
    wire t99680 = t99679 ^ t99679;
    wire t99681 = t99680 ^ t99680;
    wire t99682 = t99681 ^ t99681;
    wire t99683 = t99682 ^ t99682;
    wire t99684 = t99683 ^ t99683;
    wire t99685 = t99684 ^ t99684;
    wire t99686 = t99685 ^ t99685;
    wire t99687 = t99686 ^ t99686;
    wire t99688 = t99687 ^ t99687;
    wire t99689 = t99688 ^ t99688;
    wire t99690 = t99689 ^ t99689;
    wire t99691 = t99690 ^ t99690;
    wire t99692 = t99691 ^ t99691;
    wire t99693 = t99692 ^ t99692;
    wire t99694 = t99693 ^ t99693;
    wire t99695 = t99694 ^ t99694;
    wire t99696 = t99695 ^ t99695;
    wire t99697 = t99696 ^ t99696;
    wire t99698 = t99697 ^ t99697;
    wire t99699 = t99698 ^ t99698;
    wire t99700 = t99699 ^ t99699;
    wire t99701 = t99700 ^ t99700;
    wire t99702 = t99701 ^ t99701;
    wire t99703 = t99702 ^ t99702;
    wire t99704 = t99703 ^ t99703;
    wire t99705 = t99704 ^ t99704;
    wire t99706 = t99705 ^ t99705;
    wire t99707 = t99706 ^ t99706;
    wire t99708 = t99707 ^ t99707;
    wire t99709 = t99708 ^ t99708;
    wire t99710 = t99709 ^ t99709;
    wire t99711 = t99710 ^ t99710;
    wire t99712 = t99711 ^ t99711;
    wire t99713 = t99712 ^ t99712;
    wire t99714 = t99713 ^ t99713;
    wire t99715 = t99714 ^ t99714;
    wire t99716 = t99715 ^ t99715;
    wire t99717 = t99716 ^ t99716;
    wire t99718 = t99717 ^ t99717;
    wire t99719 = t99718 ^ t99718;
    wire t99720 = t99719 ^ t99719;
    wire t99721 = t99720 ^ t99720;
    wire t99722 = t99721 ^ t99721;
    wire t99723 = t99722 ^ t99722;
    wire t99724 = t99723 ^ t99723;
    wire t99725 = t99724 ^ t99724;
    wire t99726 = t99725 ^ t99725;
    wire t99727 = t99726 ^ t99726;
    wire t99728 = t99727 ^ t99727;
    wire t99729 = t99728 ^ t99728;
    wire t99730 = t99729 ^ t99729;
    wire t99731 = t99730 ^ t99730;
    wire t99732 = t99731 ^ t99731;
    wire t99733 = t99732 ^ t99732;
    wire t99734 = t99733 ^ t99733;
    wire t99735 = t99734 ^ t99734;
    wire t99736 = t99735 ^ t99735;
    wire t99737 = t99736 ^ t99736;
    wire t99738 = t99737 ^ t99737;
    wire t99739 = t99738 ^ t99738;
    wire t99740 = t99739 ^ t99739;
    wire t99741 = t99740 ^ t99740;
    wire t99742 = t99741 ^ t99741;
    wire t99743 = t99742 ^ t99742;
    wire t99744 = t99743 ^ t99743;
    wire t99745 = t99744 ^ t99744;
    wire t99746 = t99745 ^ t99745;
    wire t99747 = t99746 ^ t99746;
    wire t99748 = t99747 ^ t99747;
    wire t99749 = t99748 ^ t99748;
    wire t99750 = t99749 ^ t99749;
    wire t99751 = t99750 ^ t99750;
    wire t99752 = t99751 ^ t99751;
    wire t99753 = t99752 ^ t99752;
    wire t99754 = t99753 ^ t99753;
    wire t99755 = t99754 ^ t99754;
    wire t99756 = t99755 ^ t99755;
    wire t99757 = t99756 ^ t99756;
    wire t99758 = t99757 ^ t99757;
    wire t99759 = t99758 ^ t99758;
    wire t99760 = t99759 ^ t99759;
    wire t99761 = t99760 ^ t99760;
    wire t99762 = t99761 ^ t99761;
    wire t99763 = t99762 ^ t99762;
    wire t99764 = t99763 ^ t99763;
    wire t99765 = t99764 ^ t99764;
    wire t99766 = t99765 ^ t99765;
    wire t99767 = t99766 ^ t99766;
    wire t99768 = t99767 ^ t99767;
    wire t99769 = t99768 ^ t99768;
    wire t99770 = t99769 ^ t99769;
    wire t99771 = t99770 ^ t99770;
    wire t99772 = t99771 ^ t99771;
    wire t99773 = t99772 ^ t99772;
    wire t99774 = t99773 ^ t99773;
    wire t99775 = t99774 ^ t99774;
    wire t99776 = t99775 ^ t99775;
    wire t99777 = t99776 ^ t99776;
    wire t99778 = t99777 ^ t99777;
    wire t99779 = t99778 ^ t99778;
    wire t99780 = t99779 ^ t99779;
    wire t99781 = t99780 ^ t99780;
    wire t99782 = t99781 ^ t99781;
    wire t99783 = t99782 ^ t99782;
    wire t99784 = t99783 ^ t99783;
    wire t99785 = t99784 ^ t99784;
    wire t99786 = t99785 ^ t99785;
    wire t99787 = t99786 ^ t99786;
    wire t99788 = t99787 ^ t99787;
    wire t99789 = t99788 ^ t99788;
    wire t99790 = t99789 ^ t99789;
    wire t99791 = t99790 ^ t99790;
    wire t99792 = t99791 ^ t99791;
    wire t99793 = t99792 ^ t99792;
    wire t99794 = t99793 ^ t99793;
    wire t99795 = t99794 ^ t99794;
    wire t99796 = t99795 ^ t99795;
    wire t99797 = t99796 ^ t99796;
    wire t99798 = t99797 ^ t99797;
    wire t99799 = t99798 ^ t99798;
    wire t99800 = t99799 ^ t99799;
    wire t99801 = t99800 ^ t99800;
    wire t99802 = t99801 ^ t99801;
    wire t99803 = t99802 ^ t99802;
    wire t99804 = t99803 ^ t99803;
    wire t99805 = t99804 ^ t99804;
    wire t99806 = t99805 ^ t99805;
    wire t99807 = t99806 ^ t99806;
    wire t99808 = t99807 ^ t99807;
    wire t99809 = t99808 ^ t99808;
    wire t99810 = t99809 ^ t99809;
    wire t99811 = t99810 ^ t99810;
    wire t99812 = t99811 ^ t99811;
    wire t99813 = t99812 ^ t99812;
    wire t99814 = t99813 ^ t99813;
    wire t99815 = t99814 ^ t99814;
    wire t99816 = t99815 ^ t99815;
    wire t99817 = t99816 ^ t99816;
    wire t99818 = t99817 ^ t99817;
    wire t99819 = t99818 ^ t99818;
    wire t99820 = t99819 ^ t99819;
    wire t99821 = t99820 ^ t99820;
    wire t99822 = t99821 ^ t99821;
    wire t99823 = t99822 ^ t99822;
    wire t99824 = t99823 ^ t99823;
    wire t99825 = t99824 ^ t99824;
    wire t99826 = t99825 ^ t99825;
    wire t99827 = t99826 ^ t99826;
    wire t99828 = t99827 ^ t99827;
    wire t99829 = t99828 ^ t99828;
    wire t99830 = t99829 ^ t99829;
    wire t99831 = t99830 ^ t99830;
    wire t99832 = t99831 ^ t99831;
    wire t99833 = t99832 ^ t99832;
    wire t99834 = t99833 ^ t99833;
    wire t99835 = t99834 ^ t99834;
    wire t99836 = t99835 ^ t99835;
    wire t99837 = t99836 ^ t99836;
    wire t99838 = t99837 ^ t99837;
    wire t99839 = t99838 ^ t99838;
    wire t99840 = t99839 ^ t99839;
    wire t99841 = t99840 ^ t99840;
    wire t99842 = t99841 ^ t99841;
    wire t99843 = t99842 ^ t99842;
    wire t99844 = t99843 ^ t99843;
    wire t99845 = t99844 ^ t99844;
    wire t99846 = t99845 ^ t99845;
    wire t99847 = t99846 ^ t99846;
    wire t99848 = t99847 ^ t99847;
    wire t99849 = t99848 ^ t99848;
    wire t99850 = t99849 ^ t99849;
    wire t99851 = t99850 ^ t99850;
    wire t99852 = t99851 ^ t99851;
    wire t99853 = t99852 ^ t99852;
    wire t99854 = t99853 ^ t99853;
    wire t99855 = t99854 ^ t99854;
    wire t99856 = t99855 ^ t99855;
    wire t99857 = t99856 ^ t99856;
    wire t99858 = t99857 ^ t99857;
    wire t99859 = t99858 ^ t99858;
    wire t99860 = t99859 ^ t99859;
    wire t99861 = t99860 ^ t99860;
    wire t99862 = t99861 ^ t99861;
    wire t99863 = t99862 ^ t99862;
    wire t99864 = t99863 ^ t99863;
    wire t99865 = t99864 ^ t99864;
    wire t99866 = t99865 ^ t99865;
    wire t99867 = t99866 ^ t99866;
    wire t99868 = t99867 ^ t99867;
    wire t99869 = t99868 ^ t99868;
    wire t99870 = t99869 ^ t99869;
    wire t99871 = t99870 ^ t99870;
    wire t99872 = t99871 ^ t99871;
    wire t99873 = t99872 ^ t99872;
    wire t99874 = t99873 ^ t99873;
    wire t99875 = t99874 ^ t99874;
    wire t99876 = t99875 ^ t99875;
    wire t99877 = t99876 ^ t99876;
    wire t99878 = t99877 ^ t99877;
    wire t99879 = t99878 ^ t99878;
    wire t99880 = t99879 ^ t99879;
    wire t99881 = t99880 ^ t99880;
    wire t99882 = t99881 ^ t99881;
    wire t99883 = t99882 ^ t99882;
    wire t99884 = t99883 ^ t99883;
    wire t99885 = t99884 ^ t99884;
    wire t99886 = t99885 ^ t99885;
    wire t99887 = t99886 ^ t99886;
    wire t99888 = t99887 ^ t99887;
    wire t99889 = t99888 ^ t99888;
    wire t99890 = t99889 ^ t99889;
    wire t99891 = t99890 ^ t99890;
    wire t99892 = t99891 ^ t99891;
    wire t99893 = t99892 ^ t99892;
    wire t99894 = t99893 ^ t99893;
    wire t99895 = t99894 ^ t99894;
    wire t99896 = t99895 ^ t99895;
    wire t99897 = t99896 ^ t99896;
    wire t99898 = t99897 ^ t99897;
    wire t99899 = t99898 ^ t99898;
    wire t99900 = t99899 ^ t99899;
    wire t99901 = t99900 ^ t99900;
    wire t99902 = t99901 ^ t99901;
    wire t99903 = t99902 ^ t99902;
    wire t99904 = t99903 ^ t99903;
    wire t99905 = t99904 ^ t99904;
    wire t99906 = t99905 ^ t99905;
    wire t99907 = t99906 ^ t99906;
    wire t99908 = t99907 ^ t99907;
    wire t99909 = t99908 ^ t99908;
    wire t99910 = t99909 ^ t99909;
    wire t99911 = t99910 ^ t99910;
    wire t99912 = t99911 ^ t99911;
    wire t99913 = t99912 ^ t99912;
    wire t99914 = t99913 ^ t99913;
    wire t99915 = t99914 ^ t99914;
    wire t99916 = t99915 ^ t99915;
    wire t99917 = t99916 ^ t99916;
    wire t99918 = t99917 ^ t99917;
    wire t99919 = t99918 ^ t99918;
    wire t99920 = t99919 ^ t99919;
    wire t99921 = t99920 ^ t99920;
    wire t99922 = t99921 ^ t99921;
    wire t99923 = t99922 ^ t99922;
    wire t99924 = t99923 ^ t99923;
    wire t99925 = t99924 ^ t99924;
    wire t99926 = t99925 ^ t99925;
    wire t99927 = t99926 ^ t99926;
    wire t99928 = t99927 ^ t99927;
    wire t99929 = t99928 ^ t99928;
    wire t99930 = t99929 ^ t99929;
    wire t99931 = t99930 ^ t99930;
    wire t99932 = t99931 ^ t99931;
    wire t99933 = t99932 ^ t99932;
    wire t99934 = t99933 ^ t99933;
    wire t99935 = t99934 ^ t99934;
    wire t99936 = t99935 ^ t99935;
    wire t99937 = t99936 ^ t99936;
    wire t99938 = t99937 ^ t99937;
    wire t99939 = t99938 ^ t99938;
    wire t99940 = t99939 ^ t99939;
    wire t99941 = t99940 ^ t99940;
    wire t99942 = t99941 ^ t99941;
    wire t99943 = t99942 ^ t99942;
    wire t99944 = t99943 ^ t99943;
    wire t99945 = t99944 ^ t99944;
    wire t99946 = t99945 ^ t99945;
    wire t99947 = t99946 ^ t99946;
    wire t99948 = t99947 ^ t99947;
    wire t99949 = t99948 ^ t99948;
    wire t99950 = t99949 ^ t99949;
    wire t99951 = t99950 ^ t99950;
    wire t99952 = t99951 ^ t99951;
    wire t99953 = t99952 ^ t99952;
    wire t99954 = t99953 ^ t99953;
    wire t99955 = t99954 ^ t99954;
    wire t99956 = t99955 ^ t99955;
    wire t99957 = t99956 ^ t99956;
    wire t99958 = t99957 ^ t99957;
    wire t99959 = t99958 ^ t99958;
    wire t99960 = t99959 ^ t99959;
    wire t99961 = t99960 ^ t99960;
    wire t99962 = t99961 ^ t99961;
    wire t99963 = t99962 ^ t99962;
    wire t99964 = t99963 ^ t99963;
    wire t99965 = t99964 ^ t99964;
    wire t99966 = t99965 ^ t99965;
    wire t99967 = t99966 ^ t99966;
    wire t99968 = t99967 ^ t99967;
    wire t99969 = t99968 ^ t99968;
    wire t99970 = t99969 ^ t99969;
    wire t99971 = t99970 ^ t99970;
    wire t99972 = t99971 ^ t99971;
    wire t99973 = t99972 ^ t99972;
    wire t99974 = t99973 ^ t99973;
    wire t99975 = t99974 ^ t99974;
    wire t99976 = t99975 ^ t99975;
    wire t99977 = t99976 ^ t99976;
    wire t99978 = t99977 ^ t99977;
    wire t99979 = t99978 ^ t99978;
    wire t99980 = t99979 ^ t99979;
    wire t99981 = t99980 ^ t99980;
    wire t99982 = t99981 ^ t99981;
    wire t99983 = t99982 ^ t99982;
    wire t99984 = t99983 ^ t99983;
    wire t99985 = t99984 ^ t99984;
    wire t99986 = t99985 ^ t99985;
    wire t99987 = t99986 ^ t99986;
    wire t99988 = t99987 ^ t99987;
    wire t99989 = t99988 ^ t99988;
    wire t99990 = t99989 ^ t99989;
    wire t99991 = t99990 ^ t99990;
    wire t99992 = t99991 ^ t99991;
    wire t99993 = t99992 ^ t99992;
    wire t99994 = t99993 ^ t99993;
    wire t99995 = t99994 ^ t99994;
    wire t99996 = t99995 ^ t99995;
    wire t99997 = t99996 ^ t99996;
    wire t99998 = t99997 ^ t99997;
    wire z = t99998 ^ t99998;


endmodule