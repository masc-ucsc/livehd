module pick( input [2:0] a, output [2:0] x);
assign x = a[2:1];
endmodule

