/* verilator lint_off WIDTH */
module pyrm_write_back_block(
	pc_pyri,
	pc_valid_pyri,
	pc_retry_pyro,
	branch_pc_pyri,
	branch_pc_valid_pyri,
	branch_pc_retry_pyro,
	raddr_pyri,
	raddr_valid_pyri,
	raddr_retry_pyro,
	rdata_pyri,
	rdata_valid_pyri,
	rdata_retry_pyro,
	inst_pyri,
	inst_valid_pyri,
	inst_retry_pyro,
	reset_pyri,
	pc_pyro,
	pc_valid_pyro,
	pc_retry_pyri,
	branch_pc_pyro,
	branch_pc_valid_pyro,
	branch_pc_retry_pyri,
	decode_reg_addr_pyro,
	decode_reg_addr_valid_pyro,
	decode_reg_addr_retry_pyri,
	debug_reg_addr_pyro,
	debug_reg_addr_valid_pyro,
	debug_reg_addr_retry_pyri,
	decode_reg_data_pyro,
	decode_reg_data_valid_pyro,
	decode_reg_data_retry_pyri,
	debug_reg_data_pyro,
	debug_reg_data_valid_pyro,
	debug_reg_data_retry_pyri,
	clk
);


  

  

  

  

  

  


input [64-1:0] pc_pyri;
input pc_valid_pyri;
output pc_retry_pyro;
input [64-1:0] branch_pc_pyri;
input branch_pc_valid_pyri;
output branch_pc_retry_pyro;
input [64-1:0] raddr_pyri;
input raddr_valid_pyri;
output raddr_retry_pyro;
input [64-1:0] rdata_pyri;
input rdata_valid_pyri;
output rdata_retry_pyro;
input [32-1:0] inst_pyri;
input inst_valid_pyri;
output inst_retry_pyro;
input  reset_pyri;
output[64-1:0] pc_pyro;
output pc_valid_pyro;
input pc_retry_pyri;
output[64-1:0] branch_pc_pyro;
output branch_pc_valid_pyro;
input branch_pc_retry_pyri;
output[64-1:0] decode_reg_addr_pyro;
output decode_reg_addr_valid_pyro;
input decode_reg_addr_retry_pyri;
output[64-1:0] debug_reg_addr_pyro;
output debug_reg_addr_valid_pyro;
input debug_reg_addr_retry_pyri;
output[64-1:0] decode_reg_data_pyro;
output decode_reg_data_valid_pyro;
input decode_reg_data_retry_pyri;
output[64-1:0] debug_reg_data_pyro;
output debug_reg_data_valid_pyro;
input debug_reg_data_retry_pyri;
input clk;
logic [64-1:0] __tid17237;
logic [64-1:0] __tid17239;
logic dcache__write__11813;
logic debug_reg_data__write__11814;
logic debug_reg_addr__write__11815;
logic decode_reg_data__write__11816;
logic decode_reg_addr__write__11817;
logic rdata__read__11821;
logic raddr__read__11822;
logic __tid333__11897;
logic __tid341__11911;
logic __tid349__11925;
logic __tid391__11946;
logic __tid399__11960;
logic __tid407__11974;
logic __tid9539__12042;
logic branch_pc__write__12067;
logic branch_pc__read__12068;
logic decode_reg_addr__write__12073;
logic decode_reg_data__write__12077;
logic debug_reg_addr__write__12081;
logic raddr__read__12082;
logic debug_reg_data__write__12085;
logic rdata__read__12086;
logic branch_pc__write__12096;
logic branch_pc__read__12098;
logic [64-1:0] __tid9641__12109;
logic rdata__read__12110;
logic [64-1:0] dcaddr__12112;
logic [64-1:0] __tid450__12126;
logic [64-1:0] fpx10559__index__12128;
logic [64-1:0] __tid464__12131;
logic [64-1:0] __tid473__12136;
logic [64-1:0] fpx10559__first_read_remainder__12138;
logic [64-1:0] __tid481__12139;
logic __tid487__12141;
logic __tid489__12142;
logic [64-1:0] fpx10790__data__12195;
logic [64-1:0] fpx10790__data__12196;
logic [6-1:0] __tid692__12197;
logic __tid694__12198;
logic __tid696__12199;
logic __tid702__12201;
logic __tid704__12202;
logic [64-1:0] fpx10790__data__12206;
logic [64-1:0] fpx10790__data__12207;
logic [64-1:0] fpx10790__data__12210;
logic [64-1:0] fpx10790__data__12213;
logic [64-1:0] fpx10790__data__12214;
logic [6-1:0] __tid726__12215;
logic __tid728__12216;
logic __tid730__12217;
logic __tid736__12219;
logic __tid738__12220;
logic [64-1:0] fpx10790__data__12224;
logic [64-1:0] fpx10790__data__12225;
logic [64-1:0] fpx10790__data__12228;
logic [64-1:0] fpx10790__data__12231;
logic [64-1:0] fpx10790__data__12232;
logic [64-1:0] fpx10790__data__12235;
logic [64-1:0] fpx10790__data__12236;
logic [64-1:0] fpx10790__data__12239;
logic [64-1:0] fpx10790__data__12240;
logic [6-1:0] __tid772__12241;
logic __tid774__12242;
logic __tid776__12243;
logic __tid782__12245;
logic __tid784__12246;
logic [64-1:0] fpx10790__data__12250;
logic [64-1:0] fpx10790__data__12251;
logic [64-1:0] fpx10790__data__12254;
logic [64-1:0] fpx10790__data__12257;
logic [64-1:0] fpx10790__data__12258;
logic [64-1:0] __tid507__12343;
logic [64-1:0] __tid509__12345;
logic [6-1:0] __tid513__12347;
logic [64-1:0] fpx10559__result__12348;
logic [64-1:0] __tid833__12357;
logic [64-1:0] fpx10807__remainder__12359;
logic [8-1:0] fpx11255__rtrn__12365;
logic __tid1730__12384;
logic __tid1762__12406;
logic __tid1794__12428;
logic [8-1:0] fpx11255__rtrn__12437;
logic [8-1:0] fpx11255__rtrn__12440;
logic [8-1:0] fpx11255__rtrn__12443;
logic [64-1:0] __tid852__12452;
logic [64-1:0] fpx10807__bytes_after_remainder__12453;
logic [64-1:0] __tid861__12455;
logic [64-1:0] __tid535__12460;
logic [64-1:0] __tid541__12462;
logic [64-1:0] __tid543__12464;
logic [64-1:0] __tid883__12477;
logic [64-1:0] fpx10891__remainder__12479;
logic [8-1:0] __tid899__12483;
logic [8-1:0] __tid910__12488;
logic [8-1:0] fpx10891__bytes_already_read__12489;
logic __tid936__12509;
logic __tid968__12531;
logic [8-1:0] __tid1007__12548;
logic [8-1:0] fpx10891__bytes_to_read__12549;
logic [8-1:0] __tid1017__12554;
logic [8-1:0] fpx10891__bytes_to_read__12555;
logic [8-1:0] __tid1027__12560;
logic [8-1:0] fpx10891__bytes_to_read__12561;
logic [8-1:0] fpx10891__bytes_to_read__12566;
logic [64-1:0] __tid1065__12595;
logic [64-1:0] fpx10559__result__12601;
logic [6-1:0] __tid692__12783;
logic [6-1:0] __tid726__12801;
logic [6-1:0] __tid772__12827;
logic raddr__read__13187;
logic [64-1:0] __tid9682__13195;
logic [64-1:0] dcaddr__13198;
logic [64-1:0] __tid1141__13237;
logic [64-1:0] fpx10696__remainder__13239;
logic [64-1:0] __tid1152__13242;
logic [64-1:0] fpx10696__index__13244;
logic [64-1:0] fpx10696__write_overflow_val__13246;
logic fpx10696__has_overflow__13247;
logic [64-1:0] __tid1169__13248;
logic __tid1175__13250;
logic __tid1177__13251;
logic [64-1:0] fpx10696__index__13264;
logic [64-1:0] __tid1203__13265;
logic [64-1:0] fpx10696__current__13287;
logic [64-1:0] fpx10696__current__13288;
logic [64-1:0] fpx10696__current__13293;
logic [64-1:0] fpx10696__current__13294;
logic [64-1:0] fpx10696__current__13297;
logic [64-1:0] fpx10696__current__13298;
logic [64-1:0] fpx11078__data__13360;
logic [64-1:0] fpx11078__data__13361;
logic [6-1:0] __tid692__13362;
logic __tid694__13363;
logic __tid696__13364;
logic __tid702__13366;
logic __tid704__13367;
logic [64-1:0] fpx11078__data__13371;
logic [64-1:0] fpx11078__data__13372;
logic [64-1:0] fpx11078__data__13375;
logic [64-1:0] fpx11078__data__13378;
logic [64-1:0] fpx11078__data__13379;
logic [6-1:0] __tid726__13380;
logic __tid728__13381;
logic __tid730__13382;
logic __tid736__13384;
logic __tid738__13385;
logic [64-1:0] fpx11078__data__13389;
logic [64-1:0] fpx11078__data__13390;
logic [64-1:0] fpx11078__data__13393;
logic [64-1:0] fpx11078__data__13396;
logic [64-1:0] fpx11078__data__13397;
logic [64-1:0] fpx11078__data__13400;
logic [64-1:0] fpx11078__data__13401;
logic [64-1:0] fpx11078__data__13404;
logic [64-1:0] fpx11078__data__13405;
logic [6-1:0] __tid772__13406;
logic __tid774__13407;
logic __tid776__13408;
logic __tid782__13410;
logic __tid784__13411;
logic [64-1:0] fpx11078__data__13415;
logic [64-1:0] fpx11078__data__13416;
logic [64-1:0] fpx11078__data__13419;
logic [64-1:0] fpx11078__data__13422;
logic [64-1:0] fpx11078__data__13423;
logic [64-1:0] fpx11347__data__13714;
logic [64-1:0] fpx11347__data__13715;
logic [6-1:0] __tid692__13716;
logic __tid694__13717;
logic __tid696__13718;
logic __tid702__13720;
logic __tid704__13721;
logic [64-1:0] fpx11347__data__13725;
logic [64-1:0] fpx11347__data__13726;
logic [64-1:0] fpx11347__data__13729;
logic [64-1:0] fpx11347__data__13732;
logic [64-1:0] fpx11347__data__13733;
logic [6-1:0] __tid726__13734;
logic __tid728__13735;
logic __tid730__13736;
logic __tid736__13738;
logic __tid738__13739;
logic [64-1:0] fpx11347__data__13743;
logic [64-1:0] fpx11347__data__13744;
logic [64-1:0] fpx11347__data__13747;
logic [64-1:0] fpx11347__data__13750;
logic [64-1:0] fpx11347__data__13751;
logic [64-1:0] fpx11347__data__13754;
logic [64-1:0] fpx11347__data__13755;
logic [64-1:0] fpx11347__data__13758;
logic [64-1:0] fpx11347__data__13759;
logic [6-1:0] __tid772__13760;
logic __tid774__13761;
logic __tid776__13762;
logic __tid782__13764;
logic __tid784__13765;
logic [64-1:0] fpx11347__data__13769;
logic [64-1:0] fpx11347__data__13770;
logic [64-1:0] fpx11347__data__13773;
logic [64-1:0] fpx11347__data__13776;
logic [64-1:0] fpx11347__data__13777;
logic [8-1:0] fpx11703__rtrn__13870;
logic __tid1730__13889;
logic __tid1762__13911;
logic __tid1794__13933;
logic [8-1:0] fpx11703__rtrn__13942;
logic [8-1:0] fpx11703__rtrn__13945;
logic [8-1:0] fpx11703__rtrn__13948;
logic [64-1:0] __tid1944__13956;
logic [64-1:0] fpx11377__remainder__13958;
logic [64-1:0] __tid1953__13959;
logic [64-1:0] fpx11377__rtrn__13962;
logic [8-1:0] fpx11437__rtrn__14004;
logic [8-1:0] fpx11437__rtrn__14076;
logic [8-1:0] fpx11437__rtrn__14079;
logic [8-1:0] fpx11437__rtrn__14082;
logic [64-1:0] __tid1307__14180;
logic [6-1:0] fpx10696__low_bit_count__14182;
logic [64-1:0] fpx10696__index__14185;
logic [64-1:0] __tid1323__14186;
logic [64-1:0] __tid1334__14192;
logic [64-1:0] fpx10696__to_shift_out__14193;
logic [64-1:0] __tid1342__14194;
logic [6-1:0] __tid1344__14195;
logic [64-1:0] __tid1346__14196;
logic [6-1:0] __tid1348__14197;
logic [64-1:0] fpx10696__low_bits__14198;
logic [64-1:0] __tid1357__14200;
logic [64-1:0] __tid1857__14211;
logic [64-1:0] fpx11145__remainder__14213;
logic [8-1:0] fpx11496__rtrn__14217;
logic [8-1:0] fpx11496__rtrn__14274;
logic [8-1:0] fpx11496__rtrn__14277;
logic [8-1:0] fpx11496__rtrn__14280;
logic [64-1:0] __tid1872__14286;
logic [64-1:0] fpx11145__rtrn__14289;
logic [8-1:0] fpx11555__rtrn__14331;
logic [8-1:0] fpx11555__rtrn__14403;
logic [8-1:0] fpx11555__rtrn__14406;
logic [8-1:0] fpx11555__rtrn__14409;
logic [64-1:0] __tid1944__14417;
logic [64-1:0] fpx11175__remainder__14419;
logic [64-1:0] __tid1953__14420;
logic [64-1:0] fpx11175__rtrn__14423;
logic [64-1:0] fpx11194__rtrn__14466;
logic [8-1:0] fpx11614__rtrn__14472;
logic [8-1:0] fpx11614__rtrn__14544;
logic [8-1:0] fpx11614__rtrn__14547;
logic [8-1:0] fpx11614__rtrn__14550;
logic [8-1:0] fpx11762__rtrn__14572;
logic [8-1:0] fpx11762__rtrn__14635;
logic [8-1:0] fpx11762__rtrn__14638;
logic [8-1:0] fpx11762__rtrn__14641;
logic [64-1:0] __tid1944__14649;
logic [64-1:0] fpx11643__remainder__14651;
logic [64-1:0] __tid1953__14652;
logic [64-1:0] fpx11643__rtrn__14655;
logic [64-1:0] __tid1416__14687;
logic [64-1:0] __tid1422__14689;
logic [64-1:0] __tid1424__14691;
logic [64-1:0] __tid1432__14694;
logic [64-1:0] fpx10696__write_overflow_val__14833;
logic fpx10696__has_overflow__14835;
logic [64-1:0] __tid1475__14844;
logic [64-1:0] __tid1512__15420;
logic [64-1:0] __tid1518__15422;
logic dcache__write__15790;
logic __tid14922__17256;
logic __tid14938__17264;
logic __tid14942__17266;
logic __tid14944__17267;
logic __tid14948__17269;
logic __tid14954__17272;
logic __tid14960__17275;
logic __tid14966__17278;
logic __tid14972__17281;
logic [64-1:0] __tid17011__17374;
logic __tid17013__17375;
logic [64-1:0] __tid17017__17377;
logic [64-1:0] __tid17021__17379;
logic [64-1:0] __tid17027__17382;
logic [64-1:0] __tid17031__17384;
logic [64-1:0] __tid17037__17387;
logic [64-1:0] __tid17041__17389;
logic [64-1:0] __tid17047__17392;
logic [64-1:0] __tid17051__17394;
logic [64-1:0] __tid17055__17396;
logic [64-1:0] __tid17059__17398;
logic [7-1:0] __tid9503__11853;
logic [7-1:0] __tid9516__11862;
logic __tid9522__11864;
logic __tid9524__11865;
logic [7-1:0] __tid9533__11868;
logic __tid9537__11870;
logic __tid9543__11871;
logic [7-1:0] __tid323__11883;
logic __tid327__11885;
logic __tid353__11886;
logic [7-1:0] __tid329__11889;
logic __tid333__11892;
logic __tid333__11898;
logic __tid335__11899;
logic __tid359__11900;
logic [7-1:0] __tid337__11903;
logic __tid341__11906;
logic __tid341__11912;
logic __tid343__11913;
logic __tid365__11914;
logic [7-1:0] __tid345__11917;
logic __tid349__11920;
logic __tid349__11926;
logic fpx10518__rtrn__11927;
logic __tid385__11934;
logic __tid411__11935;
logic [7-1:0] __tid387__11938;
logic __tid391__11941;
logic __tid391__11947;
logic __tid393__11948;
logic __tid417__11949;
logic [7-1:0] __tid395__11952;
logic __tid399__11955;
logic __tid399__11961;
logic __tid401__11962;
logic __tid423__11963;
logic [7-1:0] __tid403__11966;
logic __tid407__11969;
logic __tid407__11975;
logic fpx10518__rtrn__11976;
logic __tid9539__12043;
logic __tid9549__12044;
logic __tid9551__12045;
logic [7-1:0] __tid9557__12048;
logic __tid9563__12050;
logic __tid9565__12051;
logic [7-1:0] __tid9571__12054;
logic __tid9577__12056;
logic __tid9579__12057;
logic __tid9581__12058;
logic __tid9583__12059;
logic __tid9585__12060;
logic __tid9587__12061;
logic __tid9589__12062;
logic __tid9591__12063;
logic __tid9583__12069;
logic __tid9587__12100;
logic [3-1:0] __tid9657__12116;
logic [3-1:0] __tid585__12150;
logic __tid591__12152;
logic __tid593__12153;
logic [3-1:0] __tid599__12156;
logic __tid605__12158;
logic __tid607__12159;
logic [3-1:0] __tid613__12162;
logic __tid619__12164;
logic __tid621__12165;
logic [3-1:0] __tid627__12168;
logic __tid633__12170;
logic __tid635__12171;
logic [3-1:0] __tid641__12174;
logic __tid647__12176;
logic __tid649__12177;
logic [3-1:0] __tid655__12180;
logic __tid661__12182;
logic __tid663__12183;
logic __tid665__12184;
logic __tid667__12185;
logic __tid669__12186;
logic __tid671__12187;
logic __tid673__12188;
logic __tid675__12189;
logic __tid677__12190;
logic __tid679__12191;
logic __tid681__12192;
logic __tid683__12193;
logic __tid667__12211;
logic __tid671__12229;
logic __tid675__12233;
logic __tid679__12237;
logic __tid683__12255;
logic [64-1:0] fpx10790__data__12259;
logic [64-1:0] fpx10790__data__12260;
logic [64-1:0] fpx10790__data__12274;
logic [64-1:0] fpx10790__data__12282;
logic [64-1:0] fpx10790__data__12290;
logic [64-1:0] fpx10790__data__12311;
logic [3-1:0] __tid1720__12370;
logic __tid1724__12372;
logic __tid1734__12373;
logic [3-1:0] __tid1726__12376;
logic __tid1730__12379;
logic __tid1730__12385;
logic __tid1740__12386;
logic __tid1742__12387;
logic [3-1:0] __tid1752__12392;
logic __tid1756__12394;
logic __tid1766__12395;
logic [3-1:0] __tid1758__12398;
logic __tid1762__12401;
logic __tid1762__12407;
logic __tid1772__12408;
logic __tid1774__12409;
logic [3-1:0] __tid1784__12414;
logic __tid1788__12416;
logic __tid1798__12417;
logic [3-1:0] __tid1790__12420;
logic __tid1794__12423;
logic __tid1794__12429;
logic __tid1804__12430;
logic __tid1806__12431;
logic __tid1808__12432;
logic __tid1810__12433;
logic __tid1812__12434;
logic __tid1814__12435;
logic __tid1810__12438;
logic __tid1814__12441;
logic [8-1:0] fpx11255__rtrn__12445;
logic [8-1:0] fpx11255__rtrn__12446;
logic [8-1:0] fpx11255__rtrn__12447;
logic [8-1:0] __tid859__12454;
logic __tid526__12456;
logic __tid528__12457;
logic [3-1:0] __tid926__12495;
logic __tid930__12497;
logic __tid940__12498;
logic [3-1:0] __tid932__12501;
logic __tid936__12504;
logic __tid936__12510;
logic __tid946__12511;
logic __tid948__12512;
logic [3-1:0] __tid958__12517;
logic __tid962__12519;
logic __tid972__12520;
logic [3-1:0] __tid964__12523;
logic __tid968__12526;
logic __tid968__12532;
logic __tid978__12533;
logic __tid980__12534;
logic [3-1:0] __tid986__12537;
logic __tid992__12539;
logic __tid994__12540;
logic __tid996__12541;
logic __tid998__12542;
logic __tid1000__12543;
logic __tid1002__12544;
logic __tid998__12550;
logic __tid1002__12556;
logic [8-1:0] fpx10891__bytes_to_read__12567;
logic [8-1:0] fpx10891__bytes_to_read__12572;
logic [8-1:0] fpx10891__bytes_to_read__12579;
logic [8-1:0] __tid1046__12588;
logic [8-1:0] fpx10891__bytes_to_shift_out__12589;
logic [8-1:0] __tid1055__12592;
logic [8-1:0] fpx10891__bits_to_shift_out__12594;
logic [8-1:0] __tid1067__12596;
logic [64-1:0] __tid1069__12597;
logic [8-1:0] __tid1071__12598;
logic [64-1:0] fpx10891__data__12599;
logic [64-1:0] fpx10559__second_read__12600;
logic [64-1:0] fpx10559__result__12602;
logic [64-1:0] fpx10559__result__12735;
logic [3-1:0] __tid585__12740;
logic __tid591__12742;
logic __tid593__12743;
logic [3-1:0] __tid599__12745;
logic __tid605__12747;
logic __tid607__12748;
logic [3-1:0] __tid613__12751;
logic __tid619__12753;
logic __tid621__12754;
logic [3-1:0] __tid627__12756;
logic __tid633__12758;
logic __tid635__12759;
logic [3-1:0] __tid641__12761;
logic __tid647__12763;
logic __tid649__12764;
logic [3-1:0] __tid655__12766;
logic __tid661__12768;
logic __tid663__12769;
logic __tid665__12770;
logic __tid667__12771;
logic __tid669__12772;
logic __tid671__12773;
logic __tid673__12774;
logic __tid675__12775;
logic __tid677__12776;
logic __tid679__12777;
logic __tid681__12778;
logic __tid683__12779;
logic [64-1:0] fpx10985__data__12781;
logic [64-1:0] fpx10985__data__12782;
logic __tid694__12784;
logic __tid696__12785;
logic __tid702__12787;
logic __tid704__12788;
logic [64-1:0] fpx10985__data__12792;
logic [64-1:0] fpx10985__data__12793;
logic [64-1:0] fpx10985__data__12796;
logic __tid667__12797;
logic [64-1:0] fpx10985__data__12799;
logic [64-1:0] fpx10985__data__12800;
logic __tid728__12802;
logic __tid730__12803;
logic __tid736__12805;
logic __tid738__12806;
logic [64-1:0] fpx10985__data__12810;
logic [64-1:0] fpx10985__data__12811;
logic [64-1:0] fpx10985__data__12814;
logic __tid671__12815;
logic [64-1:0] fpx10985__data__12817;
logic [64-1:0] fpx10985__data__12818;
logic __tid675__12819;
logic [64-1:0] fpx10985__data__12821;
logic [64-1:0] fpx10985__data__12822;
logic __tid679__12823;
logic [64-1:0] fpx10985__data__12825;
logic [64-1:0] fpx10985__data__12826;
logic __tid774__12828;
logic __tid776__12829;
logic __tid782__12831;
logic __tid784__12832;
logic [64-1:0] fpx10985__data__12836;
logic [64-1:0] fpx10985__data__12837;
logic [64-1:0] fpx10985__data__12840;
logic __tid683__12841;
logic [64-1:0] fpx10985__data__12843;
logic [64-1:0] fpx10985__data__12844;
logic [64-1:0] fpx10985__data__12845;
logic [64-1:0] fpx10985__data__12846;
logic [64-1:0] fpx10985__data__12860;
logic [64-1:0] fpx10985__data__12868;
logic [64-1:0] fpx10985__data__12876;
logic [64-1:0] fpx10985__data__12897;
logic [64-1:0] fpx10559__result__12991;
logic __tid9591__13190;
logic [32-1:0] inst__13201;
logic [3-1:0] __tid9701__13202;
logic [3-1:0] __tid1183__13256;
logic __tid1189__13258;
logic __tid1191__13259;
logic [3-1:0] __tid1212__13271;
logic __tid1218__13273;
logic __tid1220__13274;
logic [3-1:0] __tid1226__13278;
logic __tid1232__13280;
logic __tid1234__13281;
logic __tid1236__13282;
logic __tid1238__13283;
logic __tid1238__13289;
logic [64-1:0] fpx10696__current__13301;
logic [64-1:0] fpx10696__current__13306;
logic [3-1:0] __tid585__13315;
logic __tid591__13317;
logic __tid593__13318;
logic [3-1:0] __tid599__13321;
logic __tid605__13323;
logic __tid607__13324;
logic [3-1:0] __tid613__13327;
logic __tid619__13329;
logic __tid621__13330;
logic [3-1:0] __tid627__13333;
logic __tid633__13335;
logic __tid635__13336;
logic [3-1:0] __tid641__13339;
logic __tid647__13341;
logic __tid649__13342;
logic [3-1:0] __tid655__13345;
logic __tid661__13347;
logic __tid663__13348;
logic __tid665__13349;
logic __tid667__13350;
logic __tid669__13351;
logic __tid671__13352;
logic __tid673__13353;
logic __tid675__13354;
logic __tid677__13355;
logic __tid679__13356;
logic __tid681__13357;
logic __tid683__13358;
logic __tid667__13376;
logic __tid671__13394;
logic __tid675__13398;
logic __tid679__13402;
logic __tid683__13420;
logic [64-1:0] fpx11078__data__13424;
logic [64-1:0] fpx11078__data__13425;
logic [64-1:0] fpx11078__data__13439;
logic [64-1:0] fpx11078__data__13447;
logic [64-1:0] fpx11078__data__13455;
logic [64-1:0] fpx11078__data__13476;
logic [64-1:0] __tid1280__13505;
logic [64-1:0] __tid1282__13506;
logic [64-1:0] fpx10696__write_val__13507;
logic [64-1:0] fpx10696__write_val__13508;
logic [3-1:0] __tid585__13669;
logic __tid591__13671;
logic __tid593__13672;
logic [3-1:0] __tid599__13675;
logic __tid605__13677;
logic __tid607__13678;
logic [3-1:0] __tid613__13681;
logic __tid619__13683;
logic __tid621__13684;
logic [3-1:0] __tid627__13687;
logic __tid633__13689;
logic __tid635__13690;
logic [3-1:0] __tid641__13693;
logic __tid647__13695;
logic __tid649__13696;
logic [3-1:0] __tid655__13699;
logic __tid661__13701;
logic __tid663__13702;
logic __tid665__13703;
logic __tid667__13704;
logic __tid669__13705;
logic __tid671__13706;
logic __tid673__13707;
logic __tid675__13708;
logic __tid677__13709;
logic __tid679__13710;
logic __tid681__13711;
logic __tid683__13712;
logic __tid667__13730;
logic __tid671__13748;
logic __tid675__13752;
logic __tid679__13756;
logic __tid683__13774;
logic [64-1:0] fpx11347__data__13778;
logic [64-1:0] fpx11347__data__13779;
logic [64-1:0] fpx11347__data__13793;
logic [64-1:0] fpx11347__data__13801;
logic [64-1:0] fpx11347__data__13809;
logic [64-1:0] fpx11347__data__13830;
logic [3-1:0] __tid1720__13875;
logic __tid1724__13877;
logic __tid1734__13878;
logic [3-1:0] __tid1726__13881;
logic __tid1730__13884;
logic __tid1730__13890;
logic __tid1740__13891;
logic __tid1742__13892;
logic [3-1:0] __tid1752__13897;
logic __tid1756__13899;
logic __tid1766__13900;
logic [3-1:0] __tid1758__13903;
logic __tid1762__13906;
logic __tid1762__13912;
logic __tid1772__13913;
logic __tid1774__13914;
logic [3-1:0] __tid1784__13919;
logic __tid1788__13921;
logic __tid1798__13922;
logic [3-1:0] __tid1790__13925;
logic __tid1794__13928;
logic __tid1794__13934;
logic __tid1804__13935;
logic __tid1806__13936;
logic __tid1808__13937;
logic __tid1810__13938;
logic __tid1812__13939;
logic __tid1814__13940;
logic __tid1810__13943;
logic __tid1814__13946;
logic [8-1:0] fpx11703__rtrn__13950;
logic [8-1:0] fpx11703__rtrn__13951;
logic [8-1:0] fpx11703__rtrn__13952;
logic [8-1:0] __tid1955__13960;
logic [64-1:0] fpx11377__needed__13961;
logic [64-1:0] __tid1967__13965;
logic __tid1973__13967;
logic __tid1975__13968;
logic [64-1:0] __tid1981__13973;
logic [64-1:0] fpx11377__rtrn__13975;
logic [64-1:0] fpx11377__rtrn__13982;
logic [64-1:0] __tid1996__13985;
logic [64-1:0] fpx11114__overflow_bit_count__13987;
logic [8-1:0] __tid1567__13991;
logic [64-1:0] __tid1573__13993;
logic __tid1579__13995;
logic __tid1581__13996;
logic [3-1:0] __tid1720__14009;
logic __tid1724__14011;
logic __tid1734__14012;
logic [3-1:0] __tid1726__14015;
logic __tid1730__14018;
logic __tid1730__14024;
logic __tid1740__14025;
logic __tid1742__14026;
logic [3-1:0] __tid1752__14031;
logic __tid1756__14033;
logic __tid1766__14034;
logic [3-1:0] __tid1758__14037;
logic __tid1762__14040;
logic __tid1762__14046;
logic __tid1772__14047;
logic __tid1774__14048;
logic [3-1:0] __tid1784__14053;
logic __tid1788__14055;
logic __tid1798__14056;
logic [3-1:0] __tid1790__14059;
logic __tid1794__14062;
logic __tid1794__14068;
logic __tid1804__14069;
logic __tid1806__14070;
logic __tid1808__14071;
logic __tid1810__14072;
logic __tid1812__14073;
logic __tid1814__14074;
logic __tid1810__14077;
logic __tid1814__14080;
logic [8-1:0] fpx11437__rtrn__14084;
logic [8-1:0] fpx11437__rtrn__14085;
logic [8-1:0] fpx11437__rtrn__14086;
logic [8-1:0] __tid1599__14093;
logic [8-1:0] __tid1601__14094;
logic [8-1:0] __tid1605__14096;
logic [8-1:0] __tid1607__14098;
logic [8-1:0] fpx11114__to_shift_off__14099;
logic [64-1:0] __tid1615__14101;
logic [8-1:0] __tid1617__14102;
logic [64-1:0] __tid1619__14103;
logic [8-1:0] __tid1621__14104;
logic [64-1:0] fpx11114__rtrn__14105;
logic __tid1730__14119;
logic __tid1762__14130;
logic __tid1794__14141;
logic [64-1:0] fpx11114__rtrn__14176;
logic [64-1:0] fpx10696__data_low__14177;
logic [64-1:0] fpx10696__data_low__14183;
logic [64-1:0] __tid1355__14199;
logic [64-1:0] fpx10696__write_val__14201;
logic [3-1:0] __tid1720__14220;
logic __tid1724__14222;
logic __tid1734__14223;
logic [3-1:0] __tid1726__14226;
logic __tid1730__14229;
logic __tid1730__14232;
logic __tid1740__14233;
logic __tid1742__14234;
logic [3-1:0] __tid1752__14237;
logic __tid1756__14239;
logic __tid1766__14240;
logic [3-1:0] __tid1758__14243;
logic __tid1762__14246;
logic __tid1762__14249;
logic __tid1772__14250;
logic __tid1774__14251;
logic [3-1:0] __tid1784__14254;
logic __tid1788__14256;
logic __tid1798__14257;
logic [3-1:0] __tid1790__14260;
logic __tid1794__14263;
logic __tid1794__14266;
logic __tid1804__14267;
logic __tid1806__14268;
logic __tid1808__14269;
logic __tid1810__14270;
logic __tid1812__14271;
logic __tid1814__14272;
logic __tid1810__14275;
logic __tid1814__14278;
logic [8-1:0] fpx11496__rtrn__14282;
logic [8-1:0] fpx11496__rtrn__14283;
logic [8-1:0] fpx11496__rtrn__14284;
logic [8-1:0] __tid1874__14287;
logic [64-1:0] fpx11145__needed__14288;
logic [64-1:0] __tid1886__14291;
logic __tid1892__14293;
logic __tid1894__14294;
logic [64-1:0] __tid1902__14300;
logic [64-1:0] fpx11145__rtrn__14301;
logic [64-1:0] fpx11145__rtrn__14308;
logic [64-1:0] __tid1915__14310;
logic [64-1:0] fpx10696__high_bit_count__14312;
logic [64-1:0] __tid1372__14313;
logic __tid1378__14315;
logic __tid1380__14316;
logic [3-1:0] __tid1720__14336;
logic __tid1724__14338;
logic __tid1734__14339;
logic [3-1:0] __tid1726__14342;
logic __tid1730__14345;
logic __tid1730__14351;
logic __tid1740__14352;
logic __tid1742__14353;
logic [3-1:0] __tid1752__14358;
logic __tid1756__14360;
logic __tid1766__14361;
logic [3-1:0] __tid1758__14364;
logic __tid1762__14367;
logic __tid1762__14373;
logic __tid1772__14374;
logic __tid1774__14375;
logic [3-1:0] __tid1784__14380;
logic __tid1788__14382;
logic __tid1798__14383;
logic [3-1:0] __tid1790__14386;
logic __tid1794__14389;
logic __tid1794__14395;
logic __tid1804__14396;
logic __tid1806__14397;
logic __tid1808__14398;
logic __tid1810__14399;
logic __tid1812__14400;
logic __tid1814__14401;
logic __tid1810__14404;
logic __tid1814__14407;
logic [8-1:0] fpx11555__rtrn__14411;
logic [8-1:0] fpx11555__rtrn__14412;
logic [8-1:0] fpx11555__rtrn__14413;
logic [8-1:0] __tid1955__14421;
logic [64-1:0] fpx11175__needed__14422;
logic [64-1:0] __tid1967__14426;
logic __tid1973__14428;
logic __tid1975__14429;
logic [64-1:0] __tid1981__14434;
logic [64-1:0] fpx11175__rtrn__14436;
logic [64-1:0] fpx11175__rtrn__14443;
logic [64-1:0] __tid1996__14446;
logic [64-1:0] fpx10696__overflow_bit_count__14448;
logic [64-1:0] __tid1392__14449;
logic __tid1398__14451;
logic __tid1400__14452;
logic [3-1:0] __tid1720__14477;
logic __tid1724__14479;
logic __tid1734__14480;
logic [3-1:0] __tid1726__14483;
logic __tid1730__14486;
logic __tid1730__14492;
logic __tid1740__14493;
logic __tid1742__14494;
logic [3-1:0] __tid1752__14499;
logic __tid1756__14501;
logic __tid1766__14502;
logic [3-1:0] __tid1758__14505;
logic __tid1762__14508;
logic __tid1762__14514;
logic __tid1772__14515;
logic __tid1774__14516;
logic [3-1:0] __tid1784__14521;
logic __tid1788__14523;
logic __tid1798__14524;
logic [3-1:0] __tid1790__14527;
logic __tid1794__14530;
logic __tid1794__14536;
logic __tid1804__14537;
logic __tid1806__14538;
logic __tid1808__14539;
logic __tid1810__14540;
logic __tid1812__14541;
logic __tid1814__14542;
logic __tid1810__14545;
logic __tid1814__14548;
logic [8-1:0] fpx11614__rtrn__14552;
logic [8-1:0] fpx11614__rtrn__14553;
logic [8-1:0] fpx11614__rtrn__14554;
logic [8-1:0] __tid1665__14558;
logic [8-1:0] fpx11194__access_width_bits__14560;
logic [3-1:0] __tid1720__14577;
logic __tid1724__14579;
logic __tid1734__14580;
logic [3-1:0] __tid1726__14583;
logic __tid1730__14586;
logic __tid1730__14589;
logic __tid1740__14590;
logic __tid1742__14591;
logic [3-1:0] __tid1752__14596;
logic __tid1756__14598;
logic __tid1766__14599;
logic [3-1:0] __tid1758__14602;
logic __tid1762__14605;
logic __tid1762__14608;
logic __tid1772__14609;
logic __tid1774__14610;
logic [3-1:0] __tid1784__14615;
logic __tid1788__14617;
logic __tid1798__14618;
logic [3-1:0] __tid1790__14621;
logic __tid1794__14624;
logic __tid1794__14627;
logic __tid1804__14628;
logic __tid1806__14629;
logic __tid1808__14630;
logic __tid1810__14631;
logic __tid1812__14632;
logic __tid1814__14633;
logic __tid1810__14636;
logic __tid1814__14639;
logic [8-1:0] fpx11762__rtrn__14643;
logic [8-1:0] fpx11762__rtrn__14644;
logic [8-1:0] fpx11762__rtrn__14645;
logic [8-1:0] __tid1955__14653;
logic [64-1:0] fpx11643__needed__14654;
logic [64-1:0] __tid1967__14658;
logic __tid1973__14660;
logic __tid1975__14661;
logic [64-1:0] __tid1981__14666;
logic [64-1:0] fpx11643__rtrn__14668;
logic [64-1:0] fpx11643__rtrn__14675;
logic [64-1:0] __tid1996__14678;
logic [64-1:0] fpx11194__overflow_bits__14680;
logic [8-1:0] __tid1683__14681;
logic [64-1:0] __tid1685__14682;
logic [6-1:0] fpx11194__to_shift_off__14683;
logic [64-1:0] fpx11194__rtrn__14684;
logic [6-1:0] __tid1434__14696;
logic [64-1:0] __tid1436__14697;
logic [6-1:0] __tid1438__14699;
logic [64-1:0] fpx10696__high_bits__14700;
logic [64-1:0] __tid1445__14701;
logic [64-1:0] __tid1447__14702;
logic [64-1:0] fpx10696__write_overflow_val__14703;
logic [64-1:0] fpx10696__write_overflow_val__14834;
logic [64-1:0] __tid1467__14841;
logic [64-1:0] fpx10696__to_shift_out__14842;
logic [6-1:0] __tid1477__14845;
logic [64-1:0] __tid1479__14846;
logic [6-1:0] __tid1481__14847;
logic [64-1:0] fpx10696__high_bits__14848;
logic [64-1:0] fpx10696__write_val__14849;
logic [64-1:0] fpx10696__write_val__14850;
logic [64-1:0] fpx10696__write_overflow_val__14978;
logic fpx10696__has_overflow__14979;
logic [64-1:0] fpx10696__write_val__14995;
logic [64-1:0] fpx10696__write_val__15006;
logic [64-1:0] fpx10696__write_overflow_val__15405;
logic fpx10696__has_overflow__15406;
logic __tid1505__15417;
logic raddr__read__15801;
logic rdata__read__15806;
logic dcache__write__16282;
logic decode_reg_addr__write__16288;
logic raddr__read__16289;
logic [64-1:0] decode_reg_data__16290;
logic decode_reg_data__write__16291;
logic rdata__read__16292;
logic debug_reg_addr__write__16294;
logic [64-1:0] debug_reg_data__16295;
logic debug_reg_data__write__16296;
logic branch_pc__write__16302;
logic branch_pc__read__16303;
logic dcache__write__16750;
logic branch_pc__write__16756;
logic branch_pc__read__16757;
logic decode_reg_addr__write__16759;
logic raddr__read__16760;
logic decode_reg_data__write__16762;
logic rdata__read__16763;
logic debug_reg_addr__write__16766;
logic debug_reg_data__write__16769;
logic dcache__write__17216;
logic dcache__write__17228;
logic debug_reg_data__write__17229;
logic debug_reg_addr__write__17230;
logic decode_reg_data__write__17231;
logic decode_reg_addr__write__17232;
logic branch_pc__write__17233;
logic rdata__read__17236;
logic raddr__read__17237;
logic branch_pc__read__17238;
logic __tid14924__17257;
logic __tid14926__17258;
logic __tid14928__17259;
logic __tid14930__17260;
logic __tid14932__17261;
logic __tid14934__17262;
logic __tid14946__17268;
logic __tid14950__17270;
logic __tid14952__17271;
logic __tid14956__17273;
logic __tid14958__17274;
logic __tid14962__17276;
logic __tid14964__17277;
logic __tid14968__17279;
logic __tid14970__17280;
logic __tid14974__17282;
logic __tid14983__17286;
logic __tid14985__17287;
logic __tid14987__17288;
logic __tid14989__17289;
logic __tid14991__17290;
logic __tid14993__17291;
logic __tid14995__17292;
logic __tid14997__17293;
logic __tid14999__17294;
logic __tid15001__17295;
logic __block_valid__17297;
logic __tid15012__17310;
logic __tid15026__17317;
logic __tid15031__17320;
logic __tid15035__17322;
logic __tid15039__17324;
logic __tid15043__17326;
logic __tid15047__17328;
logic [64-1:0] __tid17015__17376;
logic [64-1:0] __tid17019__17378;
logic __tid17025__17381;
logic [64-1:0] __tid17029__17383;
logic __tid17035__17386;
logic [64-1:0] __tid17039__17388;
logic __tid17045__17391;
logic [64-1:0] __tid17049__17393;
logic [64-1:0] __tid17057__17397;
logic [64-1:0] __tid15978__17354;
logic [64-1:0] __tid17023__17380;
logic [64-1:0] __tid17033__17385;
logic [64-1:0] __tid17043__17390;
logic [64-1:0] __tid17053__17395;
logic [64-1:0] __tid17061__17399;
logic [64-1:0] pc_pyri;
logic pc_retry_pyro;
logic pc_valid_pyri;
logic [64-1:0] branch_pc_pyri;
logic branch_pc_retry_pyro;
logic branch_pc_valid_pyri;
logic [64-1:0] raddr_pyri;
logic raddr_retry_pyro;
logic raddr_valid_pyri;
logic [64-1:0] rdata_pyri;
logic rdata_retry_pyro;
logic rdata_valid_pyri;
logic [32-1:0] inst_pyri;
logic inst_retry_pyro;
logic inst_valid_pyri;
logic reset_pyri;
logic reset_retry_pyro;
logic reset_valid_pyri;
logic [64-1:0] dcache_pyri;
logic [64-1:0] pc_pyro;
logic pc_valid_pyro;
logic pc_retry_pyri;
logic [64-1:0] branch_pc_pyro;
logic branch_pc_valid_pyro;
logic branch_pc_retry_pyri;
logic [64-1:0] decode_reg_addr_pyro;
logic decode_reg_addr_valid_pyro;
logic decode_reg_addr_retry_pyri;
logic [64-1:0] debug_reg_addr_pyro;
logic debug_reg_addr_valid_pyro;
logic debug_reg_addr_retry_pyri;
logic [64-1:0] decode_reg_data_pyro;
logic decode_reg_data_valid_pyro;
logic decode_reg_data_retry_pyri;
logic [64-1:0] debug_reg_data_pyro;
logic debug_reg_data_valid_pyro;
logic debug_reg_data_retry_pyri;
logic [64-1:0] dcache_pyro;
logic dcache_valid_pyro;



  
    logic[63:0] dcache[2048-1:0];
  



assign dcache__write__11813 = 0; // asn dcache__write__11813, false

assign debug_reg_data__write__11814 = 0; // asn debug_reg_data__write__11814, false

assign debug_reg_addr__write__11815 = 0; // asn debug_reg_addr__write__11815, false

assign decode_reg_data__write__11816 = 0; // asn decode_reg_data__write__11816, false

assign decode_reg_addr__write__11817 = 0; // asn decode_reg_addr__write__11817, false

assign rdata__read__11821 = 0; // asn rdata__read__11821, false

assign raddr__read__11822 = 0; // asn raddr__read__11822, false

assign pc_pyro = pc_pyri; // asn pc_pyro, pc_pyri

assign __tid333__11897 = 0; // asn __tid333__11897, false

assign __tid341__11911 = 0; // asn __tid341__11911, false

assign __tid349__11925 = 0; // asn __tid349__11925, false

assign __tid391__11946 = 0; // asn __tid391__11946, false

assign __tid399__11960 = 0; // asn __tid399__11960, false

assign __tid407__11974 = 0; // asn __tid407__11974, false

assign __tid9539__12042 = 0; // asn __tid9539__12042, false

assign branch_pc__write__12067 = 1; // asn branch_pc__write__12067, true

assign branch_pc__read__12068 = 1; // asn branch_pc__read__12068, true

assign decode_reg_addr__write__12073 = 1; // asn decode_reg_addr__write__12073, true

assign decode_reg_data__write__12077 = 1; // asn decode_reg_data__write__12077, true

assign debug_reg_addr__write__12081 = 1; // asn debug_reg_addr__write__12081, true

assign raddr__read__12082 = 1; // asn raddr__read__12082, true

assign debug_reg_data__write__12085 = 1; // asn debug_reg_data__write__12085, true

assign rdata__read__12086 = 1; // asn rdata__read__12086, true

assign branch_pc__write__12096 = 0; // asn branch_pc__write__12096, false

assign branch_pc__read__12098 = 0; // asn branch_pc__read__12098, false

assign __tid9641__12109 = rdata_pyri; // asn __tid9641__12109, rdata_pyri

assign rdata__read__12110 = 1; // asn rdata__read__12110, true

assign dcaddr__12112 = __tid9641__12109 & 64'd65535; // asn dcaddr__12112, %numeric_and(__tid9641__12109, 65535<uint<64>>)

assign __tid450__12126 = dcaddr__12112; // asn __tid450__12126, dcaddr__12112

assign fpx10559__index__12128 = __tid450__12126 >> 64'd3; // asn fpx10559__index__12128, %right_shift(__tid450__12126, 3<uint<64>>)

assign __tid473__12136 = dcaddr__12112; // asn __tid473__12136, dcaddr__12112

assign fpx10559__first_read_remainder__12138 = __tid473__12136 & 64'd7; // asn fpx10559__first_read_remainder__12138, %numeric_and(__tid473__12136, 7<uint<64>>)

assign __tid481__12139 = fpx10559__first_read_remainder__12138; // asn __tid481__12139, fpx10559__first_read_remainder__12138

assign __tid487__12141 = __tid481__12139 == 64'd0; // asn __tid487__12141, %is_equal(__tid481__12139, 0<uint<64>>)

assign __tid489__12142 = __tid487__12141; // asn __tid489__12142, __tid487__12141

assign fpx10790__data__12195 = __tid464__12131; // asn fpx10790__data__12195, __tid464__12131

assign fpx10790__data__12196 = fpx10790__data__12195 & 64'd255; // asn fpx10790__data__12196, %numeric_and(fpx10790__data__12195, 255<uint<64>>)

assign __tid692__12197 = 6'd7; // asn __tid692__12197, 7<uint<6>>

assign __tid694__12198 = fpx10790__data__12196[__tid692__12197]; // asn __tid694__12198, %bit_read(fpx10790__data__12196, __tid692__12197)

assign __tid696__12199 = __tid694__12198; // asn __tid696__12199, __tid694__12198

assign __tid702__12201 = __tid696__12199 == 1'd1; // asn __tid702__12201, %is_equal(__tid696__12199, 1<uint<1>>)

assign __tid704__12202 = __tid702__12201; // asn __tid704__12202, __tid702__12201

assign fpx10790__data__12206 = fpx10790__data__12196; // asn fpx10790__data__12206, fpx10790__data__12196

assign fpx10790__data__12207 = fpx10790__data__12206 | 64'd18446744073709551360; // asn fpx10790__data__12207, %numeric_or(fpx10790__data__12206, 18446744073709551360<uint<64>>)

assign fpx10790__data__12210 = (__tid704__12202) ? fpx10790__data__12207 : fpx10790__data__12196;

assign fpx10790__data__12213 = __tid464__12131; // asn fpx10790__data__12213, __tid464__12131

assign fpx10790__data__12214 = fpx10790__data__12213 & 64'd65535; // asn fpx10790__data__12214, %numeric_and(fpx10790__data__12213, 65535<uint<64>>)

assign __tid726__12215 = 6'd15; // asn __tid726__12215, 15<uint<6>>

assign __tid728__12216 = fpx10790__data__12214[__tid726__12215]; // asn __tid728__12216, %bit_read(fpx10790__data__12214, __tid726__12215)

assign __tid730__12217 = __tid728__12216; // asn __tid730__12217, __tid728__12216

assign __tid736__12219 = __tid730__12217 == 1'd1; // asn __tid736__12219, %is_equal(__tid730__12217, 1<uint<1>>)

assign __tid738__12220 = __tid736__12219; // asn __tid738__12220, __tid736__12219

assign fpx10790__data__12224 = fpx10790__data__12214; // asn fpx10790__data__12224, fpx10790__data__12214

assign fpx10790__data__12225 = fpx10790__data__12224 | 64'd18446744073709486080; // asn fpx10790__data__12225, %numeric_or(fpx10790__data__12224, 18446744073709486080<uint<64>>)

assign fpx10790__data__12228 = (__tid738__12220) ? fpx10790__data__12225 : fpx10790__data__12214;

assign fpx10790__data__12231 = __tid464__12131; // asn fpx10790__data__12231, __tid464__12131

assign fpx10790__data__12232 = fpx10790__data__12231 & 64'd255; // asn fpx10790__data__12232, %numeric_and(fpx10790__data__12231, 255<uint<64>>)

assign fpx10790__data__12235 = __tid464__12131; // asn fpx10790__data__12235, __tid464__12131

assign fpx10790__data__12236 = fpx10790__data__12235 & 64'd65535; // asn fpx10790__data__12236, %numeric_and(fpx10790__data__12235, 65535<uint<64>>)

assign fpx10790__data__12239 = __tid464__12131; // asn fpx10790__data__12239, __tid464__12131

assign fpx10790__data__12240 = fpx10790__data__12239 & 64'd4294967295; // asn fpx10790__data__12240, %numeric_and(fpx10790__data__12239, 4294967295<uint<64>>)

assign __tid772__12241 = 6'd31; // asn __tid772__12241, 31<uint<6>>

assign __tid774__12242 = fpx10790__data__12240[__tid772__12241]; // asn __tid774__12242, %bit_read(fpx10790__data__12240, __tid772__12241)

assign __tid776__12243 = __tid774__12242; // asn __tid776__12243, __tid774__12242

assign __tid782__12245 = __tid776__12243 == 1'd1; // asn __tid782__12245, %is_equal(__tid776__12243, 1<uint<1>>)

assign __tid784__12246 = __tid782__12245; // asn __tid784__12246, __tid782__12245

assign fpx10790__data__12250 = fpx10790__data__12240; // asn fpx10790__data__12250, fpx10790__data__12240

assign fpx10790__data__12251 = fpx10790__data__12250 | 64'd18446744069414584320; // asn fpx10790__data__12251, %numeric_or(fpx10790__data__12250, 18446744069414584320<uint<64>>)

assign fpx10790__data__12254 = (__tid784__12246) ? fpx10790__data__12251 : fpx10790__data__12240;

assign fpx10790__data__12257 = __tid464__12131; // asn fpx10790__data__12257, __tid464__12131

assign fpx10790__data__12258 = fpx10790__data__12257 & 64'd4294967295; // asn fpx10790__data__12258, %numeric_and(fpx10790__data__12257, 4294967295<uint<64>>)

assign __tid507__12343 = __tid464__12131; // asn __tid507__12343, __tid464__12131

assign __tid509__12345 = fpx10559__first_read_remainder__12138; // asn __tid509__12345, fpx10559__first_read_remainder__12138

assign __tid513__12347 = __tid509__12345 << 64'd3; // asn __tid513__12347, %left_shift(__tid509__12345, 3<uint<64>>)

assign fpx10559__result__12348 = __tid507__12343 >> __tid513__12347; // asn fpx10559__result__12348, %right_shift(__tid507__12343, __tid513__12347)

assign __tid833__12357 = dcaddr__12112; // asn __tid833__12357, dcaddr__12112

assign fpx10807__remainder__12359 = __tid833__12357 & 64'd7; // asn fpx10807__remainder__12359, %numeric_and(__tid833__12357, 7<uint<64>>)

assign fpx11255__rtrn__12365 = 8'd8; // asn fpx11255__rtrn__12365, 8<uint<4>>

assign __tid1730__12384 = 0; // asn __tid1730__12384, false

assign __tid1762__12406 = 0; // asn __tid1762__12406, false

assign __tid1794__12428 = 0; // asn __tid1794__12428, false

assign fpx11255__rtrn__12437 = 8'd1; // asn fpx11255__rtrn__12437, 1<uint<8>>

assign fpx11255__rtrn__12440 = 8'd2; // asn fpx11255__rtrn__12440, 2<uint<8>>

assign fpx11255__rtrn__12443 = 8'd4; // asn fpx11255__rtrn__12443, 4<uint<8>>

assign __tid852__12452 = fpx10807__remainder__12359; // asn __tid852__12452, fpx10807__remainder__12359

assign fpx10807__bytes_after_remainder__12453 = 64'd8 - __tid852__12452; // asn fpx10807__bytes_after_remainder__12453, %subtraction(8<uint<64>>, __tid852__12452)

assign __tid861__12455 = fpx10807__bytes_after_remainder__12453; // asn __tid861__12455, fpx10807__bytes_after_remainder__12453

assign __tid535__12460 = fpx10559__index__12128; // asn __tid535__12460, fpx10559__index__12128

assign __tid541__12462 = __tid535__12460 + 64'd1; // asn __tid541__12462, %addition(__tid535__12460, 1<uint<64>>)

assign __tid883__12477 = dcaddr__12112; // asn __tid883__12477, dcaddr__12112

assign fpx10891__remainder__12479 = __tid883__12477 & 64'd7; // asn fpx10891__remainder__12479, %numeric_and(__tid883__12477, 7<uint<64>>)

assign __tid899__12483 = fpx10891__remainder__12479[7:0]; // asn __tid899__12483, %bit_read(fpx10891__remainder__12479, 7<uint<4>>, 0<uint<1>>)

assign __tid910__12488 = __tid899__12483; // asn __tid910__12488, __tid899__12483

assign fpx10891__bytes_already_read__12489 = 8'd8 - __tid910__12488; // asn fpx10891__bytes_already_read__12489, %subtraction(8<uint<8>>, __tid910__12488)

assign __tid936__12509 = 0; // asn __tid936__12509, false

assign __tid968__12531 = 0; // asn __tid968__12531, false

assign __tid1007__12548 = fpx10891__bytes_already_read__12489; // asn __tid1007__12548, fpx10891__bytes_already_read__12489

assign fpx10891__bytes_to_read__12549 = 8'd2 - __tid1007__12548; // asn fpx10891__bytes_to_read__12549, %subtraction(2<uint<8>>, __tid1007__12548)

assign __tid1017__12554 = fpx10891__bytes_already_read__12489; // asn __tid1017__12554, fpx10891__bytes_already_read__12489

assign fpx10891__bytes_to_read__12555 = 8'd4 - __tid1017__12554; // asn fpx10891__bytes_to_read__12555, %subtraction(4<uint<8>>, __tid1017__12554)

assign __tid1027__12560 = fpx10891__bytes_already_read__12489; // asn __tid1027__12560, fpx10891__bytes_already_read__12489

assign fpx10891__bytes_to_read__12561 = 8'd8 - __tid1027__12560; // asn fpx10891__bytes_to_read__12561, %subtraction(8<uint<8>>, __tid1027__12560)

assign fpx10891__bytes_to_read__12566 = 8'd0; // asn fpx10891__bytes_to_read__12566, 0<uint<8>>

assign __tid1065__12595 = __tid543__12464; // asn __tid1065__12595, __tid543__12464

assign fpx10559__result__12601 = fpx10559__result__12348; // asn fpx10559__result__12601, fpx10559__result__12348

assign __tid692__12783 = 6'd7; // asn __tid692__12783, 7<uint<6>>

assign __tid726__12801 = 6'd15; // asn __tid726__12801, 15<uint<6>>

assign __tid772__12827 = 6'd31; // asn __tid772__12827, 31<uint<6>>

assign raddr__read__13187 = 1; // asn raddr__read__13187, true

assign __tid9682__13195 = raddr_pyri; // asn __tid9682__13195, raddr_pyri

assign dcaddr__13198 = __tid9682__13195 & 64'd65535; // asn dcaddr__13198, %numeric_and(__tid9682__13195, 65535<uint<64>>)

assign __tid1141__13237 = dcaddr__13198; // asn __tid1141__13237, dcaddr__13198

assign fpx10696__remainder__13239 = __tid1141__13237 & 64'd7; // asn fpx10696__remainder__13239, %numeric_and(__tid1141__13237, 7<uint<64>>)

assign __tid1152__13242 = dcaddr__13198; // asn __tid1152__13242, dcaddr__13198

assign fpx10696__index__13244 = __tid1152__13242 >> 64'd3; // asn fpx10696__index__13244, %right_shift(__tid1152__13242, 3<uint<64>>)

assign fpx10696__write_overflow_val__13246 = 64'd0; // asn fpx10696__write_overflow_val__13246, 0<uint<1>>

assign fpx10696__has_overflow__13247 = 0; // asn fpx10696__has_overflow__13247, false

assign __tid1169__13248 = fpx10696__remainder__13239; // asn __tid1169__13248, fpx10696__remainder__13239

assign __tid1175__13250 = __tid1169__13248 == 64'd0; // asn __tid1175__13250, %is_equal(__tid1169__13248, 0<uint<64>>)

assign __tid1177__13251 = __tid1175__13250; // asn __tid1177__13251, __tid1175__13250

assign fpx10696__index__13264 = fpx10696__index__13244; // asn fpx10696__index__13264, fpx10696__index__13244

assign fpx10696__current__13287 = __tid1203__13265; // asn fpx10696__current__13287, __tid1203__13265

assign fpx10696__current__13288 = fpx10696__current__13287 & 64'd18446744069414584320; // asn fpx10696__current__13288, %numeric_and(fpx10696__current__13287, 18446744069414584320<uint<64>>)

assign fpx10696__current__13293 = __tid1203__13265; // asn fpx10696__current__13293, __tid1203__13265

assign fpx10696__current__13294 = fpx10696__current__13293 & 64'd18446744073709486080; // asn fpx10696__current__13294, %numeric_and(fpx10696__current__13293, 18446744073709486080<uint<64>>)

assign fpx10696__current__13297 = __tid1203__13265; // asn fpx10696__current__13297, __tid1203__13265

assign fpx10696__current__13298 = fpx10696__current__13297 & 64'd18446744073709551360; // asn fpx10696__current__13298, %numeric_and(fpx10696__current__13297, 18446744073709551360<uint<64>>)

assign fpx11078__data__13360 = rdata_pyri; // asn fpx11078__data__13360, rdata_pyri

assign fpx11078__data__13361 = fpx11078__data__13360 & 64'd255; // asn fpx11078__data__13361, %numeric_and(fpx11078__data__13360, 255<uint<64>>)

assign __tid692__13362 = 6'd7; // asn __tid692__13362, 7<uint<6>>

assign __tid694__13363 = fpx11078__data__13361[__tid692__13362]; // asn __tid694__13363, %bit_read(fpx11078__data__13361, __tid692__13362)

assign __tid696__13364 = __tid694__13363; // asn __tid696__13364, __tid694__13363

assign __tid702__13366 = __tid696__13364 == 1'd1; // asn __tid702__13366, %is_equal(__tid696__13364, 1<uint<1>>)

assign __tid704__13367 = __tid702__13366; // asn __tid704__13367, __tid702__13366

assign fpx11078__data__13371 = fpx11078__data__13361; // asn fpx11078__data__13371, fpx11078__data__13361

assign fpx11078__data__13372 = fpx11078__data__13371 | 64'd18446744073709551360; // asn fpx11078__data__13372, %numeric_or(fpx11078__data__13371, 18446744073709551360<uint<64>>)

assign fpx11078__data__13375 = (__tid704__13367) ? fpx11078__data__13372 : fpx11078__data__13361;

assign fpx11078__data__13378 = rdata_pyri; // asn fpx11078__data__13378, rdata_pyri

assign fpx11078__data__13379 = fpx11078__data__13378 & 64'd65535; // asn fpx11078__data__13379, %numeric_and(fpx11078__data__13378, 65535<uint<64>>)

assign __tid726__13380 = 6'd15; // asn __tid726__13380, 15<uint<6>>

assign __tid728__13381 = fpx11078__data__13379[__tid726__13380]; // asn __tid728__13381, %bit_read(fpx11078__data__13379, __tid726__13380)

assign __tid730__13382 = __tid728__13381; // asn __tid730__13382, __tid728__13381

assign __tid736__13384 = __tid730__13382 == 1'd1; // asn __tid736__13384, %is_equal(__tid730__13382, 1<uint<1>>)

assign __tid738__13385 = __tid736__13384; // asn __tid738__13385, __tid736__13384

assign fpx11078__data__13389 = fpx11078__data__13379; // asn fpx11078__data__13389, fpx11078__data__13379

assign fpx11078__data__13390 = fpx11078__data__13389 | 64'd18446744073709486080; // asn fpx11078__data__13390, %numeric_or(fpx11078__data__13389, 18446744073709486080<uint<64>>)

assign fpx11078__data__13393 = (__tid738__13385) ? fpx11078__data__13390 : fpx11078__data__13379;

assign fpx11078__data__13396 = rdata_pyri; // asn fpx11078__data__13396, rdata_pyri

assign fpx11078__data__13397 = fpx11078__data__13396 & 64'd255; // asn fpx11078__data__13397, %numeric_and(fpx11078__data__13396, 255<uint<64>>)

assign fpx11078__data__13400 = rdata_pyri; // asn fpx11078__data__13400, rdata_pyri

assign fpx11078__data__13401 = fpx11078__data__13400 & 64'd65535; // asn fpx11078__data__13401, %numeric_and(fpx11078__data__13400, 65535<uint<64>>)

assign fpx11078__data__13404 = rdata_pyri; // asn fpx11078__data__13404, rdata_pyri

assign fpx11078__data__13405 = fpx11078__data__13404 & 64'd4294967295; // asn fpx11078__data__13405, %numeric_and(fpx11078__data__13404, 4294967295<uint<64>>)

assign __tid772__13406 = 6'd31; // asn __tid772__13406, 31<uint<6>>

assign __tid774__13407 = fpx11078__data__13405[__tid772__13406]; // asn __tid774__13407, %bit_read(fpx11078__data__13405, __tid772__13406)

assign __tid776__13408 = __tid774__13407; // asn __tid776__13408, __tid774__13407

assign __tid782__13410 = __tid776__13408 == 1'd1; // asn __tid782__13410, %is_equal(__tid776__13408, 1<uint<1>>)

assign __tid784__13411 = __tid782__13410; // asn __tid784__13411, __tid782__13410

assign fpx11078__data__13415 = fpx11078__data__13405; // asn fpx11078__data__13415, fpx11078__data__13405

assign fpx11078__data__13416 = fpx11078__data__13415 | 64'd18446744069414584320; // asn fpx11078__data__13416, %numeric_or(fpx11078__data__13415, 18446744069414584320<uint<64>>)

assign fpx11078__data__13419 = (__tid784__13411) ? fpx11078__data__13416 : fpx11078__data__13405;

assign fpx11078__data__13422 = rdata_pyri; // asn fpx11078__data__13422, rdata_pyri

assign fpx11078__data__13423 = fpx11078__data__13422 & 64'd4294967295; // asn fpx11078__data__13423, %numeric_and(fpx11078__data__13422, 4294967295<uint<64>>)

assign fpx11347__data__13714 = rdata_pyri; // asn fpx11347__data__13714, rdata_pyri

assign fpx11347__data__13715 = fpx11347__data__13714 & 64'd255; // asn fpx11347__data__13715, %numeric_and(fpx11347__data__13714, 255<uint<64>>)

assign __tid692__13716 = 6'd7; // asn __tid692__13716, 7<uint<6>>

assign __tid694__13717 = fpx11347__data__13715[__tid692__13716]; // asn __tid694__13717, %bit_read(fpx11347__data__13715, __tid692__13716)

assign __tid696__13718 = __tid694__13717; // asn __tid696__13718, __tid694__13717

assign __tid702__13720 = __tid696__13718 == 1'd1; // asn __tid702__13720, %is_equal(__tid696__13718, 1<uint<1>>)

assign __tid704__13721 = __tid702__13720; // asn __tid704__13721, __tid702__13720

assign fpx11347__data__13725 = fpx11347__data__13715; // asn fpx11347__data__13725, fpx11347__data__13715

assign fpx11347__data__13726 = fpx11347__data__13725 | 64'd18446744073709551360; // asn fpx11347__data__13726, %numeric_or(fpx11347__data__13725, 18446744073709551360<uint<64>>)

assign fpx11347__data__13729 = (__tid704__13721) ? fpx11347__data__13726 : fpx11347__data__13715;

assign fpx11347__data__13732 = rdata_pyri; // asn fpx11347__data__13732, rdata_pyri

assign fpx11347__data__13733 = fpx11347__data__13732 & 64'd65535; // asn fpx11347__data__13733, %numeric_and(fpx11347__data__13732, 65535<uint<64>>)

assign __tid726__13734 = 6'd15; // asn __tid726__13734, 15<uint<6>>

assign __tid728__13735 = fpx11347__data__13733[__tid726__13734]; // asn __tid728__13735, %bit_read(fpx11347__data__13733, __tid726__13734)

assign __tid730__13736 = __tid728__13735; // asn __tid730__13736, __tid728__13735

assign __tid736__13738 = __tid730__13736 == 1'd1; // asn __tid736__13738, %is_equal(__tid730__13736, 1<uint<1>>)

assign __tid738__13739 = __tid736__13738; // asn __tid738__13739, __tid736__13738

assign fpx11347__data__13743 = fpx11347__data__13733; // asn fpx11347__data__13743, fpx11347__data__13733

assign fpx11347__data__13744 = fpx11347__data__13743 | 64'd18446744073709486080; // asn fpx11347__data__13744, %numeric_or(fpx11347__data__13743, 18446744073709486080<uint<64>>)

assign fpx11347__data__13747 = (__tid738__13739) ? fpx11347__data__13744 : fpx11347__data__13733;

assign fpx11347__data__13750 = rdata_pyri; // asn fpx11347__data__13750, rdata_pyri

assign fpx11347__data__13751 = fpx11347__data__13750 & 64'd255; // asn fpx11347__data__13751, %numeric_and(fpx11347__data__13750, 255<uint<64>>)

assign fpx11347__data__13754 = rdata_pyri; // asn fpx11347__data__13754, rdata_pyri

assign fpx11347__data__13755 = fpx11347__data__13754 & 64'd65535; // asn fpx11347__data__13755, %numeric_and(fpx11347__data__13754, 65535<uint<64>>)

assign fpx11347__data__13758 = rdata_pyri; // asn fpx11347__data__13758, rdata_pyri

assign fpx11347__data__13759 = fpx11347__data__13758 & 64'd4294967295; // asn fpx11347__data__13759, %numeric_and(fpx11347__data__13758, 4294967295<uint<64>>)

assign __tid772__13760 = 6'd31; // asn __tid772__13760, 31<uint<6>>

assign __tid774__13761 = fpx11347__data__13759[__tid772__13760]; // asn __tid774__13761, %bit_read(fpx11347__data__13759, __tid772__13760)

assign __tid776__13762 = __tid774__13761; // asn __tid776__13762, __tid774__13761

assign __tid782__13764 = __tid776__13762 == 1'd1; // asn __tid782__13764, %is_equal(__tid776__13762, 1<uint<1>>)

assign __tid784__13765 = __tid782__13764; // asn __tid784__13765, __tid782__13764

assign fpx11347__data__13769 = fpx11347__data__13759; // asn fpx11347__data__13769, fpx11347__data__13759

assign fpx11347__data__13770 = fpx11347__data__13769 | 64'd18446744069414584320; // asn fpx11347__data__13770, %numeric_or(fpx11347__data__13769, 18446744069414584320<uint<64>>)

assign fpx11347__data__13773 = (__tid784__13765) ? fpx11347__data__13770 : fpx11347__data__13759;

assign fpx11347__data__13776 = rdata_pyri; // asn fpx11347__data__13776, rdata_pyri

assign fpx11347__data__13777 = fpx11347__data__13776 & 64'd4294967295; // asn fpx11347__data__13777, %numeric_and(fpx11347__data__13776, 4294967295<uint<64>>)

assign fpx11703__rtrn__13870 = 8'd8; // asn fpx11703__rtrn__13870, 8<uint<4>>

assign __tid1730__13889 = 0; // asn __tid1730__13889, false

assign __tid1762__13911 = 0; // asn __tid1762__13911, false

assign __tid1794__13933 = 0; // asn __tid1794__13933, false

assign fpx11703__rtrn__13942 = 8'd1; // asn fpx11703__rtrn__13942, 1<uint<8>>

assign fpx11703__rtrn__13945 = 8'd2; // asn fpx11703__rtrn__13945, 2<uint<8>>

assign fpx11703__rtrn__13948 = 8'd4; // asn fpx11703__rtrn__13948, 4<uint<8>>

assign __tid1944__13956 = dcaddr__13198; // asn __tid1944__13956, dcaddr__13198

assign fpx11377__remainder__13958 = __tid1944__13956 & 64'd7; // asn fpx11377__remainder__13958, %numeric_and(__tid1944__13956, 7<uint<64>>)

assign __tid1953__13959 = fpx11377__remainder__13958; // asn __tid1953__13959, fpx11377__remainder__13958

assign fpx11377__rtrn__13962 = 64'd0; // asn fpx11377__rtrn__13962, 0<uint<1>>

assign fpx11437__rtrn__14004 = 8'd8; // asn fpx11437__rtrn__14004, 8<uint<4>>

assign fpx11437__rtrn__14076 = 8'd1; // asn fpx11437__rtrn__14076, 1<uint<8>>

assign fpx11437__rtrn__14079 = 8'd2; // asn fpx11437__rtrn__14079, 2<uint<8>>

assign fpx11437__rtrn__14082 = 8'd4; // asn fpx11437__rtrn__14082, 4<uint<8>>

assign __tid1307__14180 = fpx10696__remainder__13239; // asn __tid1307__14180, fpx10696__remainder__13239

assign fpx10696__low_bit_count__14182 = __tid1307__14180 << 64'd3; // asn fpx10696__low_bit_count__14182, %left_shift(__tid1307__14180, 3<uint<64>>)

assign fpx10696__index__14185 = fpx10696__index__13244; // asn fpx10696__index__14185, fpx10696__index__13244

assign __tid1334__14192 = fpx10696__low_bit_count__14182; // asn __tid1334__14192, fpx10696__low_bit_count__14182

assign fpx10696__to_shift_out__14193 = 64'd64 - __tid1334__14192; // asn fpx10696__to_shift_out__14193, %subtraction(64<uint<64>>, __tid1334__14192)

assign __tid1342__14194 = __tid1323__14186; // asn __tid1342__14194, __tid1323__14186

assign __tid1344__14195 = fpx10696__to_shift_out__14193; // asn __tid1344__14195, fpx10696__to_shift_out__14193

assign __tid1346__14196 = __tid1342__14194 << __tid1344__14195; // asn __tid1346__14196, %left_shift(__tid1342__14194, __tid1344__14195)

assign __tid1348__14197 = fpx10696__to_shift_out__14193; // asn __tid1348__14197, fpx10696__to_shift_out__14193

assign fpx10696__low_bits__14198 = __tid1346__14196 >> __tid1348__14197; // asn fpx10696__low_bits__14198, %right_shift(__tid1346__14196, __tid1348__14197)

assign __tid1357__14200 = fpx10696__low_bits__14198; // asn __tid1357__14200, fpx10696__low_bits__14198

assign __tid1857__14211 = dcaddr__13198; // asn __tid1857__14211, dcaddr__13198

assign fpx11145__remainder__14213 = __tid1857__14211 & 64'd7; // asn fpx11145__remainder__14213, %numeric_and(__tid1857__14211, 7<uint<64>>)

assign fpx11496__rtrn__14217 = 8'd8; // asn fpx11496__rtrn__14217, 8<uint<4>>

assign fpx11496__rtrn__14274 = 8'd1; // asn fpx11496__rtrn__14274, 1<uint<8>>

assign fpx11496__rtrn__14277 = 8'd2; // asn fpx11496__rtrn__14277, 2<uint<8>>

assign fpx11496__rtrn__14280 = 8'd4; // asn fpx11496__rtrn__14280, 4<uint<8>>

assign __tid1872__14286 = fpx11145__remainder__14213; // asn __tid1872__14286, fpx11145__remainder__14213

assign fpx11145__rtrn__14289 = 64'd0; // asn fpx11145__rtrn__14289, 0<uint<1>>

assign fpx11555__rtrn__14331 = 8'd8; // asn fpx11555__rtrn__14331, 8<uint<4>>

assign fpx11555__rtrn__14403 = 8'd1; // asn fpx11555__rtrn__14403, 1<uint<8>>

assign fpx11555__rtrn__14406 = 8'd2; // asn fpx11555__rtrn__14406, 2<uint<8>>

assign fpx11555__rtrn__14409 = 8'd4; // asn fpx11555__rtrn__14409, 4<uint<8>>

assign __tid1944__14417 = dcaddr__13198; // asn __tid1944__14417, dcaddr__13198

assign fpx11175__remainder__14419 = __tid1944__14417 & 64'd7; // asn fpx11175__remainder__14419, %numeric_and(__tid1944__14417, 7<uint<64>>)

assign __tid1953__14420 = fpx11175__remainder__14419; // asn __tid1953__14420, fpx11175__remainder__14419

assign fpx11175__rtrn__14423 = 64'd0; // asn fpx11175__rtrn__14423, 0<uint<1>>

assign fpx11194__rtrn__14466 = rdata_pyri; // asn fpx11194__rtrn__14466, rdata_pyri

assign fpx11614__rtrn__14472 = 8'd8; // asn fpx11614__rtrn__14472, 8<uint<4>>

assign fpx11614__rtrn__14544 = 8'd1; // asn fpx11614__rtrn__14544, 1<uint<8>>

assign fpx11614__rtrn__14547 = 8'd2; // asn fpx11614__rtrn__14547, 2<uint<8>>

assign fpx11614__rtrn__14550 = 8'd4; // asn fpx11614__rtrn__14550, 4<uint<8>>

assign fpx11762__rtrn__14572 = 8'd8; // asn fpx11762__rtrn__14572, 8<uint<4>>

assign fpx11762__rtrn__14635 = 8'd1; // asn fpx11762__rtrn__14635, 1<uint<8>>

assign fpx11762__rtrn__14638 = 8'd2; // asn fpx11762__rtrn__14638, 2<uint<8>>

assign fpx11762__rtrn__14641 = 8'd4; // asn fpx11762__rtrn__14641, 4<uint<8>>

assign __tid1944__14649 = dcaddr__13198; // asn __tid1944__14649, dcaddr__13198

assign fpx11643__remainder__14651 = __tid1944__14649 & 64'd7; // asn fpx11643__remainder__14651, %numeric_and(__tid1944__14649, 7<uint<64>>)

assign __tid1953__14652 = fpx11643__remainder__14651; // asn __tid1953__14652, fpx11643__remainder__14651

assign fpx11643__rtrn__14655 = 64'd0; // asn fpx11643__rtrn__14655, 0<uint<1>>

assign __tid1416__14687 = fpx10696__index__13244; // asn __tid1416__14687, fpx10696__index__13244

assign __tid1422__14689 = __tid1416__14687 + 64'd1; // asn __tid1422__14689, %addition(__tid1416__14687, 1<uint<64>>)

assign __tid1432__14694 = __tid1424__14691; // asn __tid1432__14694, __tid1424__14691

assign fpx10696__write_overflow_val__14833 = 64'd0; // asn fpx10696__write_overflow_val__14833, 0<uint<1>>

assign fpx10696__has_overflow__14835 = 0; // asn fpx10696__has_overflow__14835, false

assign __tid1475__14844 = __tid1323__14186; // asn __tid1475__14844, __tid1323__14186

assign __tid1512__15420 = fpx10696__index__13244; // asn __tid1512__15420, fpx10696__index__13244

assign __tid1518__15422 = __tid1512__15420 + 64'd1; // asn __tid1518__15422, %addition(__tid1512__15420, 1<uint<64>>)

assign dcache__write__15790 = 0; // asn dcache__write__15790, false

assign branch_pc_pyro = branch_pc_pyri; // asn branch_pc_pyro, branch_pc_pyri

assign decode_reg_addr_pyro = raddr_pyri; // asn decode_reg_addr_pyro, raddr_pyri

assign debug_reg_addr_pyro = raddr_pyri; // asn debug_reg_addr_pyro, raddr_pyri

assign __tid14922__17256 = pc_valid_pyri; // asn __tid14922__17256, pc_valid_pyri

assign __tid14938__17264 = inst_valid_pyri; // asn __tid14938__17264, inst_valid_pyri

assign __tid14942__17266 = ! pc_retry_pyri; // asn __tid14942__17266, %logical_not(pc_retry_pyri)

assign __tid14944__17267 = __tid14942__17266; // asn __tid14944__17267, __tid14942__17266

assign __tid14948__17269 = ! branch_pc_retry_pyri; // asn __tid14948__17269, %logical_not(branch_pc_retry_pyri)

assign __tid14954__17272 = ! decode_reg_addr_retry_pyri; // asn __tid14954__17272, %logical_not(decode_reg_addr_retry_pyri)

assign __tid14960__17275 = ! decode_reg_data_retry_pyri; // asn __tid14960__17275, %logical_not(decode_reg_data_retry_pyri)

assign __tid14966__17278 = ! debug_reg_addr_retry_pyri; // asn __tid14966__17278, %logical_not(debug_reg_addr_retry_pyri)

assign __tid14972__17281 = ! debug_reg_data_retry_pyri; // asn __tid14972__17281, %logical_not(debug_reg_data_retry_pyri)

assign dcache_valid_pyro = 1; // asn dcache_valid_pyro, true

assign __tid17013__17375 = __tid1518__15422 == fpx10696__index__13244; // asn __tid17013__17375, %is_equal(__tid1518__15422, fpx10696__index__13244)

assign __tid9503__11853 = inst_pyri[6:0]; // asn __tid9503__11853, %bit_read(inst_pyri, 6<uint<4>>, 0<uint<1>>)

assign __tid9516__11862 = __tid9503__11853; // asn __tid9516__11862, __tid9503__11853

assign __tid9522__11864 = __tid9516__11862 == 7'd99; // asn __tid9522__11864, %is_equal(__tid9516__11862, 99<uint<7>>)

assign __tid9524__11865 = __tid9522__11864; // asn __tid9524__11865, __tid9522__11864

assign __tid9533__11868 = __tid9503__11853; // asn __tid9533__11868, __tid9503__11853

assign __tid9537__11870 = __tid9533__11868 == 7'd103; // asn __tid9537__11870, %is_equal(__tid9533__11868, 103<uint<7>>)

assign __tid9543__11871 = ! __tid9537__11870; // asn __tid9543__11871, %logical_not(__tid9537__11870)

assign __tid323__11883 = __tid9503__11853; // asn __tid323__11883, __tid9503__11853

assign __tid327__11885 = __tid323__11883 == 7'd51; // asn __tid327__11885, %is_equal(__tid323__11883, 51<uint<7>>)

assign __tid353__11886 = ! __tid327__11885; // asn __tid353__11886, %logical_not(__tid327__11885)

assign __tid329__11889 = __tid9503__11853; // asn __tid329__11889, __tid9503__11853

assign __tid333__11892 = __tid329__11889 == 7'd19; // asn __tid333__11892, %is_equal(__tid329__11889, 19<uint<7>>)

assign __tid333__11898 = (__tid353__11886) ? __tid333__11892 : __tid333__11897;

assign __tid335__11899 = __tid327__11885 | __tid333__11898; // asn __tid335__11899, %logical_or(__tid327__11885, __tid333__11898)

assign __tid359__11900 = ! __tid335__11899; // asn __tid359__11900, %logical_not(__tid335__11899)

assign __tid337__11903 = __tid9503__11853; // asn __tid337__11903, __tid9503__11853

assign __tid341__11906 = __tid337__11903 == 7'd59; // asn __tid341__11906, %is_equal(__tid337__11903, 59<uint<7>>)

assign __tid341__11912 = (__tid359__11900) ? __tid341__11906 : __tid341__11911;

assign __tid343__11913 = __tid335__11899 | __tid341__11912; // asn __tid343__11913, %logical_or(__tid335__11899, __tid341__11912)

assign __tid365__11914 = ! __tid343__11913; // asn __tid365__11914, %logical_not(__tid343__11913)

assign __tid345__11917 = __tid9503__11853; // asn __tid345__11917, __tid9503__11853

assign __tid349__11920 = __tid345__11917 == 7'd27; // asn __tid349__11920, %is_equal(__tid345__11917, 27<uint<7>>)

assign __tid349__11926 = (__tid365__11914) ? __tid349__11920 : __tid349__11925;

assign fpx10518__rtrn__11927 = __tid343__11913 | __tid349__11926; // asn fpx10518__rtrn__11927, %logical_or(__tid343__11913, __tid349__11926)

assign __tid385__11934 = fpx10518__rtrn__11927; // asn __tid385__11934, fpx10518__rtrn__11927

assign __tid411__11935 = ! __tid385__11934; // asn __tid411__11935, %logical_not(__tid385__11934)

assign __tid387__11938 = __tid9503__11853; // asn __tid387__11938, __tid9503__11853

assign __tid391__11941 = __tid387__11938 == 7'd55; // asn __tid391__11941, %is_equal(__tid387__11938, 55<uint<7>>)

assign __tid391__11947 = (__tid411__11935) ? __tid391__11941 : __tid391__11946;

assign __tid393__11948 = __tid385__11934 | __tid391__11947; // asn __tid393__11948, %logical_or(__tid385__11934, __tid391__11947)

assign __tid417__11949 = ! __tid393__11948; // asn __tid417__11949, %logical_not(__tid393__11948)

assign __tid395__11952 = __tid9503__11853; // asn __tid395__11952, __tid9503__11853

assign __tid399__11955 = __tid395__11952 == 7'd23; // asn __tid399__11955, %is_equal(__tid395__11952, 23<uint<7>>)

assign __tid399__11961 = (__tid417__11949) ? __tid399__11955 : __tid399__11960;

assign __tid401__11962 = __tid393__11948 | __tid399__11961; // asn __tid401__11962, %logical_or(__tid393__11948, __tid399__11961)

assign __tid423__11963 = ! __tid401__11962; // asn __tid423__11963, %logical_not(__tid401__11962)

assign __tid403__11966 = __tid9503__11853; // asn __tid403__11966, __tid9503__11853

assign __tid407__11969 = __tid403__11966 == 7'd111; // asn __tid407__11969, %is_equal(__tid403__11966, 111<uint<7>>)

assign __tid407__11975 = (__tid423__11963) ? __tid407__11969 : __tid407__11974;

assign fpx10518__rtrn__11976 = __tid401__11962 | __tid407__11975; // asn fpx10518__rtrn__11976, %logical_or(__tid401__11962, __tid407__11975)

assign __tid9539__12043 = (__tid9543__11871) ? fpx10518__rtrn__11976 : __tid9539__12042;

assign __tid9549__12044 = __tid9537__11870 | __tid9539__12043; // asn __tid9549__12044, %logical_or(__tid9537__11870, __tid9539__12043)

assign __tid9551__12045 = __tid9549__12044; // asn __tid9551__12045, __tid9549__12044

assign __tid9557__12048 = __tid9503__11853; // asn __tid9557__12048, __tid9503__11853

assign __tid9563__12050 = __tid9557__12048 == 7'd3; // asn __tid9563__12050, %is_equal(__tid9557__12048, 3<uint<7>>)

assign __tid9565__12051 = __tid9563__12050; // asn __tid9565__12051, __tid9563__12050

assign __tid9571__12054 = __tid9503__11853; // asn __tid9571__12054, __tid9503__11853

assign __tid9577__12056 = __tid9571__12054 == 7'd35; // asn __tid9577__12056, %is_equal(__tid9571__12054, 35<uint<7>>)

assign __tid9579__12057 = __tid9577__12056; // asn __tid9579__12057, __tid9577__12056

assign __tid9581__12058 = ! __tid9524__11865; // asn __tid9581__12058, %logical_not(__tid9524__11865)

assign __tid9583__12059 = __tid9581__12058 & __tid9551__12045; // asn __tid9583__12059, %logical_and(__tid9581__12058, __tid9551__12045)

assign __tid9585__12060 = ! __tid9583__12059; // asn __tid9585__12060, %logical_not(__tid9583__12059)

assign __tid9587__12061 = __tid9585__12060 & __tid9565__12051; // asn __tid9587__12061, %logical_and(__tid9585__12060, __tid9565__12051)

assign __tid9589__12062 = ! __tid9587__12061; // asn __tid9589__12062, %logical_not(__tid9587__12061)

assign __tid9591__12063 = __tid9589__12062 & __tid9579__12057; // asn __tid9591__12063, %logical_and(__tid9589__12062, __tid9579__12057)

assign __tid9583__12069 = __tid9583__12059; // asn __tid9583__12069, __tid9583__12059

assign __tid9587__12100 = __tid9587__12061; // asn __tid9587__12100, __tid9587__12061

assign __tid9657__12116 = inst_pyri[14:12]; // asn __tid9657__12116, %bit_read(inst_pyri, 14<uint<5>>, 12<uint<5>>)

assign __tid585__12150 = __tid9657__12116; // asn __tid585__12150, __tid9657__12116

assign __tid591__12152 = __tid585__12150 == 3'd0; // asn __tid591__12152, %is_equal(__tid585__12150, 0<uint<3>>)

assign __tid593__12153 = __tid591__12152; // asn __tid593__12153, __tid591__12152

assign __tid599__12156 = __tid9657__12116; // asn __tid599__12156, __tid9657__12116

assign __tid605__12158 = __tid599__12156 == 3'd1; // asn __tid605__12158, %is_equal(__tid599__12156, 1<uint<3>>)

assign __tid607__12159 = __tid605__12158; // asn __tid607__12159, __tid605__12158

assign __tid613__12162 = __tid9657__12116; // asn __tid613__12162, __tid9657__12116

assign __tid619__12164 = __tid613__12162 == 3'd4; // asn __tid619__12164, %is_equal(__tid613__12162, 4<uint<3>>)

assign __tid621__12165 = __tid619__12164; // asn __tid621__12165, __tid619__12164

assign __tid627__12168 = __tid9657__12116; // asn __tid627__12168, __tid9657__12116

assign __tid633__12170 = { 1'd0, __tid627__12168 } == 4'd5; // asn __tid633__12170, %is_equal(__tid627__12168, 5<uint<4>>)

assign __tid635__12171 = __tid633__12170; // asn __tid635__12171, __tid633__12170

assign __tid641__12174 = __tid9657__12116; // asn __tid641__12174, __tid9657__12116

assign __tid647__12176 = __tid641__12174 == 3'd2; // asn __tid647__12176, %is_equal(__tid641__12174, 2<uint<3>>)

assign __tid649__12177 = __tid647__12176; // asn __tid649__12177, __tid647__12176

assign __tid655__12180 = __tid9657__12116; // asn __tid655__12180, __tid9657__12116

assign __tid661__12182 = { 1'd0, __tid655__12180 } == 4'd6; // asn __tid661__12182, %is_equal(__tid655__12180, 6<uint<4>>)

assign __tid663__12183 = __tid661__12182; // asn __tid663__12183, __tid661__12182

assign __tid665__12184 = ! __tid593__12153; // asn __tid665__12184, %logical_not(__tid593__12153)

assign __tid667__12185 = __tid665__12184 & __tid607__12159; // asn __tid667__12185, %logical_and(__tid665__12184, __tid607__12159)

assign __tid669__12186 = ! __tid667__12185; // asn __tid669__12186, %logical_not(__tid667__12185)

assign __tid671__12187 = __tid669__12186 & __tid621__12165; // asn __tid671__12187, %logical_and(__tid669__12186, __tid621__12165)

assign __tid673__12188 = ! __tid671__12187; // asn __tid673__12188, %logical_not(__tid671__12187)

assign __tid675__12189 = __tid673__12188 & __tid635__12171; // asn __tid675__12189, %logical_and(__tid673__12188, __tid635__12171)

assign __tid677__12190 = ! __tid675__12189; // asn __tid677__12190, %logical_not(__tid675__12189)

assign __tid679__12191 = __tid677__12190 & __tid649__12177; // asn __tid679__12191, %logical_and(__tid677__12190, __tid649__12177)

assign __tid681__12192 = ! __tid679__12191; // asn __tid681__12192, %logical_not(__tid679__12191)

assign __tid683__12193 = __tid681__12192 & __tid663__12183; // asn __tid683__12193, %logical_and(__tid681__12192, __tid663__12183)

assign __tid667__12211 = __tid667__12185; // asn __tid667__12211, __tid667__12185

assign __tid671__12229 = __tid671__12187; // asn __tid671__12229, __tid671__12187

assign __tid675__12233 = __tid675__12189; // asn __tid675__12233, __tid675__12189

assign __tid679__12237 = __tid679__12191; // asn __tid679__12237, __tid679__12191

assign __tid683__12255 = __tid683__12193; // asn __tid683__12255, __tid683__12193

assign fpx10790__data__12259 = (__tid683__12255) ? fpx10790__data__12258 : __tid464__12131;

assign fpx10790__data__12260 = (__tid679__12237) ? fpx10790__data__12254 : fpx10790__data__12259;

assign fpx10790__data__12274 = (__tid675__12233) ? fpx10790__data__12236 : fpx10790__data__12260;

assign fpx10790__data__12282 = (__tid671__12229) ? fpx10790__data__12232 : fpx10790__data__12274;

assign fpx10790__data__12290 = (__tid667__12211) ? fpx10790__data__12228 : fpx10790__data__12282;

assign fpx10790__data__12311 = (__tid593__12153) ? fpx10790__data__12210 : fpx10790__data__12290;

assign __tid1720__12370 = __tid9657__12116; // asn __tid1720__12370, __tid9657__12116

assign __tid1724__12372 = __tid1720__12370 == 3'd0; // asn __tid1724__12372, %is_equal(__tid1720__12370, 0<uint<3>>)

assign __tid1734__12373 = ! __tid1724__12372; // asn __tid1734__12373, %logical_not(__tid1724__12372)

assign __tid1726__12376 = __tid9657__12116; // asn __tid1726__12376, __tid9657__12116

assign __tid1730__12379 = __tid1726__12376 == 3'd4; // asn __tid1730__12379, %is_equal(__tid1726__12376, 4<uint<3>>)

assign __tid1730__12385 = (__tid1734__12373) ? __tid1730__12379 : __tid1730__12384;

assign __tid1740__12386 = __tid1724__12372 | __tid1730__12385; // asn __tid1740__12386, %logical_or(__tid1724__12372, __tid1730__12385)

assign __tid1742__12387 = __tid1740__12386; // asn __tid1742__12387, __tid1740__12386

assign __tid1752__12392 = __tid9657__12116; // asn __tid1752__12392, __tid9657__12116

assign __tid1756__12394 = __tid1752__12392 == 3'd1; // asn __tid1756__12394, %is_equal(__tid1752__12392, 1<uint<3>>)

assign __tid1766__12395 = ! __tid1756__12394; // asn __tid1766__12395, %logical_not(__tid1756__12394)

assign __tid1758__12398 = __tid9657__12116; // asn __tid1758__12398, __tid9657__12116

assign __tid1762__12401 = { 1'd0, __tid1758__12398 } == 4'd5; // asn __tid1762__12401, %is_equal(__tid1758__12398, 5<uint<4>>)

assign __tid1762__12407 = (__tid1766__12395) ? __tid1762__12401 : __tid1762__12406;

assign __tid1772__12408 = __tid1756__12394 | __tid1762__12407; // asn __tid1772__12408, %logical_or(__tid1756__12394, __tid1762__12407)

assign __tid1774__12409 = __tid1772__12408; // asn __tid1774__12409, __tid1772__12408

assign __tid1784__12414 = __tid9657__12116; // asn __tid1784__12414, __tid9657__12116

assign __tid1788__12416 = __tid1784__12414 == 3'd2; // asn __tid1788__12416, %is_equal(__tid1784__12414, 2<uint<3>>)

assign __tid1798__12417 = ! __tid1788__12416; // asn __tid1798__12417, %logical_not(__tid1788__12416)

assign __tid1790__12420 = __tid9657__12116; // asn __tid1790__12420, __tid9657__12116

assign __tid1794__12423 = { 1'd0, __tid1790__12420 } == 4'd6; // asn __tid1794__12423, %is_equal(__tid1790__12420, 6<uint<4>>)

assign __tid1794__12429 = (__tid1798__12417) ? __tid1794__12423 : __tid1794__12428;

assign __tid1804__12430 = __tid1788__12416 | __tid1794__12429; // asn __tid1804__12430, %logical_or(__tid1788__12416, __tid1794__12429)

assign __tid1806__12431 = __tid1804__12430; // asn __tid1806__12431, __tid1804__12430

assign __tid1808__12432 = ! __tid1742__12387; // asn __tid1808__12432, %logical_not(__tid1742__12387)

assign __tid1810__12433 = __tid1808__12432 & __tid1774__12409; // asn __tid1810__12433, %logical_and(__tid1808__12432, __tid1774__12409)

assign __tid1812__12434 = ! __tid1810__12433; // asn __tid1812__12434, %logical_not(__tid1810__12433)

assign __tid1814__12435 = __tid1812__12434 & __tid1806__12431; // asn __tid1814__12435, %logical_and(__tid1812__12434, __tid1806__12431)

assign __tid1810__12438 = __tid1810__12433; // asn __tid1810__12438, __tid1810__12433

assign __tid1814__12441 = __tid1814__12435; // asn __tid1814__12441, __tid1814__12435

assign fpx11255__rtrn__12445 = (__tid1814__12441) ? fpx11255__rtrn__12443 : fpx11255__rtrn__12365;

assign fpx11255__rtrn__12446 = (__tid1810__12438) ? fpx11255__rtrn__12440 : fpx11255__rtrn__12445;

assign fpx11255__rtrn__12447 = (__tid1742__12387) ? fpx11255__rtrn__12437 : fpx11255__rtrn__12446;

assign __tid859__12454 = fpx11255__rtrn__12447; // asn __tid859__12454, fpx11255__rtrn__12447

assign __tid526__12456 = { 56'd0, __tid859__12454 } > __tid861__12455; // asn __tid526__12456, %greater_than(__tid859__12454, __tid861__12455)

assign __tid528__12457 = __tid526__12456; // asn __tid528__12457, __tid526__12456

assign __tid926__12495 = __tid9657__12116; // asn __tid926__12495, __tid9657__12116

assign __tid930__12497 = __tid926__12495 == 3'd1; // asn __tid930__12497, %is_equal(__tid926__12495, 1<uint<3>>)

assign __tid940__12498 = ! __tid930__12497; // asn __tid940__12498, %logical_not(__tid930__12497)

assign __tid932__12501 = __tid9657__12116; // asn __tid932__12501, __tid9657__12116

assign __tid936__12504 = { 1'd0, __tid932__12501 } == 4'd5; // asn __tid936__12504, %is_equal(__tid932__12501, 5<uint<4>>)

assign __tid936__12510 = (__tid940__12498) ? __tid936__12504 : __tid936__12509;

assign __tid946__12511 = __tid930__12497 | __tid936__12510; // asn __tid946__12511, %logical_or(__tid930__12497, __tid936__12510)

assign __tid948__12512 = __tid946__12511; // asn __tid948__12512, __tid946__12511

assign __tid958__12517 = __tid9657__12116; // asn __tid958__12517, __tid9657__12116

assign __tid962__12519 = __tid958__12517 == 3'd2; // asn __tid962__12519, %is_equal(__tid958__12517, 2<uint<3>>)

assign __tid972__12520 = ! __tid962__12519; // asn __tid972__12520, %logical_not(__tid962__12519)

assign __tid964__12523 = __tid9657__12116; // asn __tid964__12523, __tid9657__12116

assign __tid968__12526 = { 1'd0, __tid964__12523 } == 4'd6; // asn __tid968__12526, %is_equal(__tid964__12523, 6<uint<4>>)

assign __tid968__12532 = (__tid972__12520) ? __tid968__12526 : __tid968__12531;

assign __tid978__12533 = __tid962__12519 | __tid968__12532; // asn __tid978__12533, %logical_or(__tid962__12519, __tid968__12532)

assign __tid980__12534 = __tid978__12533; // asn __tid980__12534, __tid978__12533

assign __tid986__12537 = __tid9657__12116; // asn __tid986__12537, __tid9657__12116

assign __tid992__12539 = __tid986__12537 == 3'd3; // asn __tid992__12539, %is_equal(__tid986__12537, 3<uint<3>>)

assign __tid994__12540 = __tid992__12539; // asn __tid994__12540, __tid992__12539

assign __tid996__12541 = ! __tid948__12512; // asn __tid996__12541, %logical_not(__tid948__12512)

assign __tid998__12542 = __tid996__12541 & __tid980__12534; // asn __tid998__12542, %logical_and(__tid996__12541, __tid980__12534)

assign __tid1000__12543 = ! __tid998__12542; // asn __tid1000__12543, %logical_not(__tid998__12542)

assign __tid1002__12544 = __tid1000__12543 & __tid994__12540; // asn __tid1002__12544, %logical_and(__tid1000__12543, __tid994__12540)

assign __tid998__12550 = __tid998__12542; // asn __tid998__12550, __tid998__12542

assign __tid1002__12556 = __tid1002__12544; // asn __tid1002__12556, __tid1002__12544

assign fpx10891__bytes_to_read__12567 = (__tid1002__12556) ? fpx10891__bytes_to_read__12561 : fpx10891__bytes_to_read__12566;

assign fpx10891__bytes_to_read__12572 = (__tid998__12550) ? fpx10891__bytes_to_read__12555 : fpx10891__bytes_to_read__12567;

assign fpx10891__bytes_to_read__12579 = (__tid948__12512) ? fpx10891__bytes_to_read__12549 : fpx10891__bytes_to_read__12572;

assign __tid1046__12588 = fpx10891__bytes_to_read__12579; // asn __tid1046__12588, fpx10891__bytes_to_read__12579

assign fpx10891__bytes_to_shift_out__12589 = 8'd8 - __tid1046__12588; // asn fpx10891__bytes_to_shift_out__12589, %subtraction(8<uint<8>>, __tid1046__12588)

assign __tid1055__12592 = fpx10891__bytes_to_shift_out__12589; // asn __tid1055__12592, fpx10891__bytes_to_shift_out__12589

assign fpx10891__bits_to_shift_out__12594 = __tid1055__12592 << 8'd3; // asn fpx10891__bits_to_shift_out__12594, %left_shift(__tid1055__12592, 3<uint<8>>)

assign __tid1067__12596 = fpx10891__bits_to_shift_out__12594; // asn __tid1067__12596, fpx10891__bits_to_shift_out__12594

assign __tid1069__12597 = __tid1065__12595 << __tid1067__12596; // asn __tid1069__12597, %left_shift(__tid1065__12595, __tid1067__12596)

assign __tid1071__12598 = fpx10891__bits_to_shift_out__12594; // asn __tid1071__12598, fpx10891__bits_to_shift_out__12594

assign fpx10891__data__12599 = __tid1069__12597 >> __tid1071__12598; // asn fpx10891__data__12599, %right_shift(__tid1069__12597, __tid1071__12598)

assign fpx10559__second_read__12600 = fpx10891__data__12599; // asn fpx10559__second_read__12600, fpx10891__data__12599

assign fpx10559__result__12602 = fpx10559__result__12601 | fpx10559__second_read__12600; // asn fpx10559__result__12602, %numeric_or(fpx10559__result__12601, fpx10559__second_read__12600)

assign fpx10559__result__12735 = (__tid528__12457) ? fpx10559__result__12602 : fpx10559__result__12348;

assign __tid585__12740 = __tid9657__12116; // asn __tid585__12740, __tid9657__12116

assign __tid591__12742 = __tid585__12740 == 3'd0; // asn __tid591__12742, %is_equal(__tid585__12740, 0<uint<3>>)

assign __tid593__12743 = __tid591__12742; // asn __tid593__12743, __tid591__12742

assign __tid599__12745 = __tid9657__12116; // asn __tid599__12745, __tid9657__12116

assign __tid605__12747 = __tid599__12745 == 3'd1; // asn __tid605__12747, %is_equal(__tid599__12745, 1<uint<3>>)

assign __tid607__12748 = __tid605__12747; // asn __tid607__12748, __tid605__12747

assign __tid613__12751 = __tid9657__12116; // asn __tid613__12751, __tid9657__12116

assign __tid619__12753 = __tid613__12751 == 3'd4; // asn __tid619__12753, %is_equal(__tid613__12751, 4<uint<3>>)

assign __tid621__12754 = __tid619__12753; // asn __tid621__12754, __tid619__12753

assign __tid627__12756 = __tid9657__12116; // asn __tid627__12756, __tid9657__12116

assign __tid633__12758 = { 1'd0, __tid627__12756 } == 4'd5; // asn __tid633__12758, %is_equal(__tid627__12756, 5<uint<4>>)

assign __tid635__12759 = __tid633__12758; // asn __tid635__12759, __tid633__12758

assign __tid641__12761 = __tid9657__12116; // asn __tid641__12761, __tid9657__12116

assign __tid647__12763 = __tid641__12761 == 3'd2; // asn __tid647__12763, %is_equal(__tid641__12761, 2<uint<3>>)

assign __tid649__12764 = __tid647__12763; // asn __tid649__12764, __tid647__12763

assign __tid655__12766 = __tid9657__12116; // asn __tid655__12766, __tid9657__12116

assign __tid661__12768 = { 1'd0, __tid655__12766 } == 4'd6; // asn __tid661__12768, %is_equal(__tid655__12766, 6<uint<4>>)

assign __tid663__12769 = __tid661__12768; // asn __tid663__12769, __tid661__12768

assign __tid665__12770 = ! __tid593__12743; // asn __tid665__12770, %logical_not(__tid593__12743)

assign __tid667__12771 = __tid665__12770 & __tid607__12748; // asn __tid667__12771, %logical_and(__tid665__12770, __tid607__12748)

assign __tid669__12772 = ! __tid667__12771; // asn __tid669__12772, %logical_not(__tid667__12771)

assign __tid671__12773 = __tid669__12772 & __tid621__12754; // asn __tid671__12773, %logical_and(__tid669__12772, __tid621__12754)

assign __tid673__12774 = ! __tid671__12773; // asn __tid673__12774, %logical_not(__tid671__12773)

assign __tid675__12775 = __tid673__12774 & __tid635__12759; // asn __tid675__12775, %logical_and(__tid673__12774, __tid635__12759)

assign __tid677__12776 = ! __tid675__12775; // asn __tid677__12776, %logical_not(__tid675__12775)

assign __tid679__12777 = __tid677__12776 & __tid649__12764; // asn __tid679__12777, %logical_and(__tid677__12776, __tid649__12764)

assign __tid681__12778 = ! __tid679__12777; // asn __tid681__12778, %logical_not(__tid679__12777)

assign __tid683__12779 = __tid681__12778 & __tid663__12769; // asn __tid683__12779, %logical_and(__tid681__12778, __tid663__12769)

assign fpx10985__data__12781 = fpx10559__result__12735; // asn fpx10985__data__12781, fpx10559__result__12735

assign fpx10985__data__12782 = fpx10985__data__12781 & 64'd255; // asn fpx10985__data__12782, %numeric_and(fpx10985__data__12781, 255<uint<64>>)

assign __tid694__12784 = fpx10985__data__12782[__tid692__12783]; // asn __tid694__12784, %bit_read(fpx10985__data__12782, __tid692__12783)

assign __tid696__12785 = __tid694__12784; // asn __tid696__12785, __tid694__12784

assign __tid702__12787 = __tid696__12785 == 1'd1; // asn __tid702__12787, %is_equal(__tid696__12785, 1<uint<1>>)

assign __tid704__12788 = __tid702__12787; // asn __tid704__12788, __tid702__12787

assign fpx10985__data__12792 = fpx10985__data__12782; // asn fpx10985__data__12792, fpx10985__data__12782

assign fpx10985__data__12793 = fpx10985__data__12792 | 64'd18446744073709551360; // asn fpx10985__data__12793, %numeric_or(fpx10985__data__12792, 18446744073709551360<uint<64>>)

assign fpx10985__data__12796 = (__tid704__12788) ? fpx10985__data__12793 : fpx10985__data__12782;

assign __tid667__12797 = __tid667__12771; // asn __tid667__12797, __tid667__12771

assign fpx10985__data__12799 = fpx10559__result__12735; // asn fpx10985__data__12799, fpx10559__result__12735

assign fpx10985__data__12800 = fpx10985__data__12799 & 64'd65535; // asn fpx10985__data__12800, %numeric_and(fpx10985__data__12799, 65535<uint<64>>)

assign __tid728__12802 = fpx10985__data__12800[__tid726__12801]; // asn __tid728__12802, %bit_read(fpx10985__data__12800, __tid726__12801)

assign __tid730__12803 = __tid728__12802; // asn __tid730__12803, __tid728__12802

assign __tid736__12805 = __tid730__12803 == 1'd1; // asn __tid736__12805, %is_equal(__tid730__12803, 1<uint<1>>)

assign __tid738__12806 = __tid736__12805; // asn __tid738__12806, __tid736__12805

assign fpx10985__data__12810 = fpx10985__data__12800; // asn fpx10985__data__12810, fpx10985__data__12800

assign fpx10985__data__12811 = fpx10985__data__12810 | 64'd18446744073709486080; // asn fpx10985__data__12811, %numeric_or(fpx10985__data__12810, 18446744073709486080<uint<64>>)

assign fpx10985__data__12814 = (__tid738__12806) ? fpx10985__data__12811 : fpx10985__data__12800;

assign __tid671__12815 = __tid671__12773; // asn __tid671__12815, __tid671__12773

assign fpx10985__data__12817 = fpx10559__result__12735; // asn fpx10985__data__12817, fpx10559__result__12735

assign fpx10985__data__12818 = fpx10985__data__12817 & 64'd255; // asn fpx10985__data__12818, %numeric_and(fpx10985__data__12817, 255<uint<64>>)

assign __tid675__12819 = __tid675__12775; // asn __tid675__12819, __tid675__12775

assign fpx10985__data__12821 = fpx10559__result__12735; // asn fpx10985__data__12821, fpx10559__result__12735

assign fpx10985__data__12822 = fpx10985__data__12821 & 64'd65535; // asn fpx10985__data__12822, %numeric_and(fpx10985__data__12821, 65535<uint<64>>)

assign __tid679__12823 = __tid679__12777; // asn __tid679__12823, __tid679__12777

assign fpx10985__data__12825 = fpx10559__result__12735; // asn fpx10985__data__12825, fpx10559__result__12735

assign fpx10985__data__12826 = fpx10985__data__12825 & 64'd4294967295; // asn fpx10985__data__12826, %numeric_and(fpx10985__data__12825, 4294967295<uint<64>>)

assign __tid774__12828 = fpx10985__data__12826[__tid772__12827]; // asn __tid774__12828, %bit_read(fpx10985__data__12826, __tid772__12827)

assign __tid776__12829 = __tid774__12828; // asn __tid776__12829, __tid774__12828

assign __tid782__12831 = __tid776__12829 == 1'd1; // asn __tid782__12831, %is_equal(__tid776__12829, 1<uint<1>>)

assign __tid784__12832 = __tid782__12831; // asn __tid784__12832, __tid782__12831

assign fpx10985__data__12836 = fpx10985__data__12826; // asn fpx10985__data__12836, fpx10985__data__12826

assign fpx10985__data__12837 = fpx10985__data__12836 | 64'd18446744069414584320; // asn fpx10985__data__12837, %numeric_or(fpx10985__data__12836, 18446744069414584320<uint<64>>)

assign fpx10985__data__12840 = (__tid784__12832) ? fpx10985__data__12837 : fpx10985__data__12826;

assign __tid683__12841 = __tid683__12779; // asn __tid683__12841, __tid683__12779

assign fpx10985__data__12843 = fpx10559__result__12735; // asn fpx10985__data__12843, fpx10559__result__12735

assign fpx10985__data__12844 = fpx10985__data__12843 & 64'd4294967295; // asn fpx10985__data__12844, %numeric_and(fpx10985__data__12843, 4294967295<uint<64>>)

assign fpx10985__data__12845 = (__tid683__12841) ? fpx10985__data__12844 : fpx10559__result__12735;

assign fpx10985__data__12846 = (__tid679__12823) ? fpx10985__data__12840 : fpx10985__data__12845;

assign fpx10985__data__12860 = (__tid675__12819) ? fpx10985__data__12822 : fpx10985__data__12846;

assign fpx10985__data__12868 = (__tid671__12815) ? fpx10985__data__12818 : fpx10985__data__12860;

assign fpx10985__data__12876 = (__tid667__12797) ? fpx10985__data__12814 : fpx10985__data__12868;

assign fpx10985__data__12897 = (__tid593__12743) ? fpx10985__data__12796 : fpx10985__data__12876;

assign fpx10559__result__12991 = (__tid489__12142) ? fpx10790__data__12311 : fpx10985__data__12897;

assign __tid9591__13190 = __tid9591__12063; // asn __tid9591__13190, __tid9591__12063

assign inst__13201 = inst_pyri; // asn inst__13201, inst_pyri

assign __tid9701__13202 = inst__13201[14:12]; // asn __tid9701__13202, %bit_read(inst__13201, 14<uint<5>>, 12<uint<5>>)

assign __tid1183__13256 = __tid9701__13202; // asn __tid1183__13256, __tid9701__13202

assign __tid1189__13258 = __tid1183__13256 == 3'd3; // asn __tid1189__13258, %is_equal(__tid1183__13256, 3<uint<3>>)

assign __tid1191__13259 = __tid1189__13258; // asn __tid1191__13259, __tid1189__13258

assign __tid1212__13271 = __tid9701__13202; // asn __tid1212__13271, __tid9701__13202

assign __tid1218__13273 = __tid1212__13271 == 3'd2; // asn __tid1218__13273, %is_equal(__tid1212__13271, 2<uint<3>>)

assign __tid1220__13274 = __tid1218__13273; // asn __tid1220__13274, __tid1218__13273

assign __tid1226__13278 = __tid9701__13202; // asn __tid1226__13278, __tid9701__13202

assign __tid1232__13280 = __tid1226__13278 == 3'd1; // asn __tid1232__13280, %is_equal(__tid1226__13278, 1<uint<3>>)

assign __tid1234__13281 = __tid1232__13280; // asn __tid1234__13281, __tid1232__13280

assign __tid1236__13282 = ! __tid1220__13274; // asn __tid1236__13282, %logical_not(__tid1220__13274)

assign __tid1238__13283 = __tid1236__13282 & __tid1234__13281; // asn __tid1238__13283, %logical_and(__tid1236__13282, __tid1234__13281)

assign __tid1238__13289 = __tid1238__13283; // asn __tid1238__13289, __tid1238__13283

assign fpx10696__current__13301 = (__tid1238__13289) ? fpx10696__current__13294 : fpx10696__current__13298;

assign fpx10696__current__13306 = (__tid1220__13274) ? fpx10696__current__13288 : fpx10696__current__13301;

assign __tid585__13315 = __tid9701__13202; // asn __tid585__13315, __tid9701__13202

assign __tid591__13317 = __tid585__13315 == 3'd0; // asn __tid591__13317, %is_equal(__tid585__13315, 0<uint<3>>)

assign __tid593__13318 = __tid591__13317; // asn __tid593__13318, __tid591__13317

assign __tid599__13321 = __tid9701__13202; // asn __tid599__13321, __tid9701__13202

assign __tid605__13323 = __tid599__13321 == 3'd1; // asn __tid605__13323, %is_equal(__tid599__13321, 1<uint<3>>)

assign __tid607__13324 = __tid605__13323; // asn __tid607__13324, __tid605__13323

assign __tid613__13327 = __tid9701__13202; // asn __tid613__13327, __tid9701__13202

assign __tid619__13329 = __tid613__13327 == 3'd4; // asn __tid619__13329, %is_equal(__tid613__13327, 4<uint<3>>)

assign __tid621__13330 = __tid619__13329; // asn __tid621__13330, __tid619__13329

assign __tid627__13333 = __tid9701__13202; // asn __tid627__13333, __tid9701__13202

assign __tid633__13335 = { 1'd0, __tid627__13333 } == 4'd5; // asn __tid633__13335, %is_equal(__tid627__13333, 5<uint<4>>)

assign __tid635__13336 = __tid633__13335; // asn __tid635__13336, __tid633__13335

assign __tid641__13339 = __tid9701__13202; // asn __tid641__13339, __tid9701__13202

assign __tid647__13341 = __tid641__13339 == 3'd2; // asn __tid647__13341, %is_equal(__tid641__13339, 2<uint<3>>)

assign __tid649__13342 = __tid647__13341; // asn __tid649__13342, __tid647__13341

assign __tid655__13345 = __tid9701__13202; // asn __tid655__13345, __tid9701__13202

assign __tid661__13347 = { 1'd0, __tid655__13345 } == 4'd6; // asn __tid661__13347, %is_equal(__tid655__13345, 6<uint<4>>)

assign __tid663__13348 = __tid661__13347; // asn __tid663__13348, __tid661__13347

assign __tid665__13349 = ! __tid593__13318; // asn __tid665__13349, %logical_not(__tid593__13318)

assign __tid667__13350 = __tid665__13349 & __tid607__13324; // asn __tid667__13350, %logical_and(__tid665__13349, __tid607__13324)

assign __tid669__13351 = ! __tid667__13350; // asn __tid669__13351, %logical_not(__tid667__13350)

assign __tid671__13352 = __tid669__13351 & __tid621__13330; // asn __tid671__13352, %logical_and(__tid669__13351, __tid621__13330)

assign __tid673__13353 = ! __tid671__13352; // asn __tid673__13353, %logical_not(__tid671__13352)

assign __tid675__13354 = __tid673__13353 & __tid635__13336; // asn __tid675__13354, %logical_and(__tid673__13353, __tid635__13336)

assign __tid677__13355 = ! __tid675__13354; // asn __tid677__13355, %logical_not(__tid675__13354)

assign __tid679__13356 = __tid677__13355 & __tid649__13342; // asn __tid679__13356, %logical_and(__tid677__13355, __tid649__13342)

assign __tid681__13357 = ! __tid679__13356; // asn __tid681__13357, %logical_not(__tid679__13356)

assign __tid683__13358 = __tid681__13357 & __tid663__13348; // asn __tid683__13358, %logical_and(__tid681__13357, __tid663__13348)

assign __tid667__13376 = __tid667__13350; // asn __tid667__13376, __tid667__13350

assign __tid671__13394 = __tid671__13352; // asn __tid671__13394, __tid671__13352

assign __tid675__13398 = __tid675__13354; // asn __tid675__13398, __tid675__13354

assign __tid679__13402 = __tid679__13356; // asn __tid679__13402, __tid679__13356

assign __tid683__13420 = __tid683__13358; // asn __tid683__13420, __tid683__13358

assign fpx11078__data__13424 = (__tid683__13420) ? fpx11078__data__13423 : rdata_pyri;

assign fpx11078__data__13425 = (__tid679__13402) ? fpx11078__data__13419 : fpx11078__data__13424;

assign fpx11078__data__13439 = (__tid675__13398) ? fpx11078__data__13401 : fpx11078__data__13425;

assign fpx11078__data__13447 = (__tid671__13394) ? fpx11078__data__13397 : fpx11078__data__13439;

assign fpx11078__data__13455 = (__tid667__13376) ? fpx11078__data__13393 : fpx11078__data__13447;

assign fpx11078__data__13476 = (__tid593__13318) ? fpx11078__data__13375 : fpx11078__data__13455;

assign __tid1280__13505 = fpx10696__current__13306; // asn __tid1280__13505, fpx10696__current__13306

assign __tid1282__13506 = fpx11078__data__13476; // asn __tid1282__13506, fpx11078__data__13476

assign fpx10696__write_val__13507 = __tid1280__13505 | __tid1282__13506; // asn fpx10696__write_val__13507, %numeric_or(__tid1280__13505, __tid1282__13506)

assign fpx10696__write_val__13508 = (__tid1191__13259) ? rdata_pyri : fpx10696__write_val__13507;

assign __tid585__13669 = __tid9701__13202; // asn __tid585__13669, __tid9701__13202

assign __tid591__13671 = __tid585__13669 == 3'd0; // asn __tid591__13671, %is_equal(__tid585__13669, 0<uint<3>>)

assign __tid593__13672 = __tid591__13671; // asn __tid593__13672, __tid591__13671

assign __tid599__13675 = __tid9701__13202; // asn __tid599__13675, __tid9701__13202

assign __tid605__13677 = __tid599__13675 == 3'd1; // asn __tid605__13677, %is_equal(__tid599__13675, 1<uint<3>>)

assign __tid607__13678 = __tid605__13677; // asn __tid607__13678, __tid605__13677

assign __tid613__13681 = __tid9701__13202; // asn __tid613__13681, __tid9701__13202

assign __tid619__13683 = __tid613__13681 == 3'd4; // asn __tid619__13683, %is_equal(__tid613__13681, 4<uint<3>>)

assign __tid621__13684 = __tid619__13683; // asn __tid621__13684, __tid619__13683

assign __tid627__13687 = __tid9701__13202; // asn __tid627__13687, __tid9701__13202

assign __tid633__13689 = { 1'd0, __tid627__13687 } == 4'd5; // asn __tid633__13689, %is_equal(__tid627__13687, 5<uint<4>>)

assign __tid635__13690 = __tid633__13689; // asn __tid635__13690, __tid633__13689

assign __tid641__13693 = __tid9701__13202; // asn __tid641__13693, __tid9701__13202

assign __tid647__13695 = __tid641__13693 == 3'd2; // asn __tid647__13695, %is_equal(__tid641__13693, 2<uint<3>>)

assign __tid649__13696 = __tid647__13695; // asn __tid649__13696, __tid647__13695

assign __tid655__13699 = __tid9701__13202; // asn __tid655__13699, __tid9701__13202

assign __tid661__13701 = { 1'd0, __tid655__13699 } == 4'd6; // asn __tid661__13701, %is_equal(__tid655__13699, 6<uint<4>>)

assign __tid663__13702 = __tid661__13701; // asn __tid663__13702, __tid661__13701

assign __tid665__13703 = ! __tid593__13672; // asn __tid665__13703, %logical_not(__tid593__13672)

assign __tid667__13704 = __tid665__13703 & __tid607__13678; // asn __tid667__13704, %logical_and(__tid665__13703, __tid607__13678)

assign __tid669__13705 = ! __tid667__13704; // asn __tid669__13705, %logical_not(__tid667__13704)

assign __tid671__13706 = __tid669__13705 & __tid621__13684; // asn __tid671__13706, %logical_and(__tid669__13705, __tid621__13684)

assign __tid673__13707 = ! __tid671__13706; // asn __tid673__13707, %logical_not(__tid671__13706)

assign __tid675__13708 = __tid673__13707 & __tid635__13690; // asn __tid675__13708, %logical_and(__tid673__13707, __tid635__13690)

assign __tid677__13709 = ! __tid675__13708; // asn __tid677__13709, %logical_not(__tid675__13708)

assign __tid679__13710 = __tid677__13709 & __tid649__13696; // asn __tid679__13710, %logical_and(__tid677__13709, __tid649__13696)

assign __tid681__13711 = ! __tid679__13710; // asn __tid681__13711, %logical_not(__tid679__13710)

assign __tid683__13712 = __tid681__13711 & __tid663__13702; // asn __tid683__13712, %logical_and(__tid681__13711, __tid663__13702)

assign __tid667__13730 = __tid667__13704; // asn __tid667__13730, __tid667__13704

assign __tid671__13748 = __tid671__13706; // asn __tid671__13748, __tid671__13706

assign __tid675__13752 = __tid675__13708; // asn __tid675__13752, __tid675__13708

assign __tid679__13756 = __tid679__13710; // asn __tid679__13756, __tid679__13710

assign __tid683__13774 = __tid683__13712; // asn __tid683__13774, __tid683__13712

assign fpx11347__data__13778 = (__tid683__13774) ? fpx11347__data__13777 : rdata_pyri;

assign fpx11347__data__13779 = (__tid679__13756) ? fpx11347__data__13773 : fpx11347__data__13778;

assign fpx11347__data__13793 = (__tid675__13752) ? fpx11347__data__13755 : fpx11347__data__13779;

assign fpx11347__data__13801 = (__tid671__13748) ? fpx11347__data__13751 : fpx11347__data__13793;

assign fpx11347__data__13809 = (__tid667__13730) ? fpx11347__data__13747 : fpx11347__data__13801;

assign fpx11347__data__13830 = (__tid593__13672) ? fpx11347__data__13729 : fpx11347__data__13809;

assign __tid1720__13875 = __tid9701__13202; // asn __tid1720__13875, __tid9701__13202

assign __tid1724__13877 = __tid1720__13875 == 3'd0; // asn __tid1724__13877, %is_equal(__tid1720__13875, 0<uint<3>>)

assign __tid1734__13878 = ! __tid1724__13877; // asn __tid1734__13878, %logical_not(__tid1724__13877)

assign __tid1726__13881 = __tid9701__13202; // asn __tid1726__13881, __tid9701__13202

assign __tid1730__13884 = __tid1726__13881 == 3'd4; // asn __tid1730__13884, %is_equal(__tid1726__13881, 4<uint<3>>)

assign __tid1730__13890 = (__tid1734__13878) ? __tid1730__13884 : __tid1730__13889;

assign __tid1740__13891 = __tid1724__13877 | __tid1730__13890; // asn __tid1740__13891, %logical_or(__tid1724__13877, __tid1730__13890)

assign __tid1742__13892 = __tid1740__13891; // asn __tid1742__13892, __tid1740__13891

assign __tid1752__13897 = __tid9701__13202; // asn __tid1752__13897, __tid9701__13202

assign __tid1756__13899 = __tid1752__13897 == 3'd1; // asn __tid1756__13899, %is_equal(__tid1752__13897, 1<uint<3>>)

assign __tid1766__13900 = ! __tid1756__13899; // asn __tid1766__13900, %logical_not(__tid1756__13899)

assign __tid1758__13903 = __tid9701__13202; // asn __tid1758__13903, __tid9701__13202

assign __tid1762__13906 = { 1'd0, __tid1758__13903 } == 4'd5; // asn __tid1762__13906, %is_equal(__tid1758__13903, 5<uint<4>>)

assign __tid1762__13912 = (__tid1766__13900) ? __tid1762__13906 : __tid1762__13911;

assign __tid1772__13913 = __tid1756__13899 | __tid1762__13912; // asn __tid1772__13913, %logical_or(__tid1756__13899, __tid1762__13912)

assign __tid1774__13914 = __tid1772__13913; // asn __tid1774__13914, __tid1772__13913

assign __tid1784__13919 = __tid9701__13202; // asn __tid1784__13919, __tid9701__13202

assign __tid1788__13921 = __tid1784__13919 == 3'd2; // asn __tid1788__13921, %is_equal(__tid1784__13919, 2<uint<3>>)

assign __tid1798__13922 = ! __tid1788__13921; // asn __tid1798__13922, %logical_not(__tid1788__13921)

assign __tid1790__13925 = __tid9701__13202; // asn __tid1790__13925, __tid9701__13202

assign __tid1794__13928 = { 1'd0, __tid1790__13925 } == 4'd6; // asn __tid1794__13928, %is_equal(__tid1790__13925, 6<uint<4>>)

assign __tid1794__13934 = (__tid1798__13922) ? __tid1794__13928 : __tid1794__13933;

assign __tid1804__13935 = __tid1788__13921 | __tid1794__13934; // asn __tid1804__13935, %logical_or(__tid1788__13921, __tid1794__13934)

assign __tid1806__13936 = __tid1804__13935; // asn __tid1806__13936, __tid1804__13935

assign __tid1808__13937 = ! __tid1742__13892; // asn __tid1808__13937, %logical_not(__tid1742__13892)

assign __tid1810__13938 = __tid1808__13937 & __tid1774__13914; // asn __tid1810__13938, %logical_and(__tid1808__13937, __tid1774__13914)

assign __tid1812__13939 = ! __tid1810__13938; // asn __tid1812__13939, %logical_not(__tid1810__13938)

assign __tid1814__13940 = __tid1812__13939 & __tid1806__13936; // asn __tid1814__13940, %logical_and(__tid1812__13939, __tid1806__13936)

assign __tid1810__13943 = __tid1810__13938; // asn __tid1810__13943, __tid1810__13938

assign __tid1814__13946 = __tid1814__13940; // asn __tid1814__13946, __tid1814__13940

assign fpx11703__rtrn__13950 = (__tid1814__13946) ? fpx11703__rtrn__13948 : fpx11703__rtrn__13870;

assign fpx11703__rtrn__13951 = (__tid1810__13943) ? fpx11703__rtrn__13945 : fpx11703__rtrn__13950;

assign fpx11703__rtrn__13952 = (__tid1742__13892) ? fpx11703__rtrn__13942 : fpx11703__rtrn__13951;

assign __tid1955__13960 = fpx11703__rtrn__13952; // asn __tid1955__13960, fpx11703__rtrn__13952

assign fpx11377__needed__13961 = __tid1953__13959 + { 56'd0, __tid1955__13960 }; // asn fpx11377__needed__13961, %addition(__tid1953__13959, __tid1955__13960)

assign __tid1967__13965 = fpx11377__needed__13961; // asn __tid1967__13965, fpx11377__needed__13961

assign __tid1973__13967 = __tid1967__13965 > 64'd8; // asn __tid1973__13967, %greater_than(__tid1967__13965, 8<uint<64>>)

assign __tid1975__13968 = __tid1973__13967; // asn __tid1975__13968, __tid1973__13967

assign __tid1981__13973 = fpx11377__needed__13961; // asn __tid1981__13973, fpx11377__needed__13961

assign fpx11377__rtrn__13975 = __tid1981__13973 - 64'd8; // asn fpx11377__rtrn__13975, %subtraction(__tid1981__13973, 8<uint<64>>)

assign fpx11377__rtrn__13982 = (__tid1975__13968) ? fpx11377__rtrn__13975 : fpx11377__rtrn__13962;

assign __tid1996__13985 = fpx11377__rtrn__13982; // asn __tid1996__13985, fpx11377__rtrn__13982

assign fpx11114__overflow_bit_count__13987 = __tid1996__13985 << 64'd3; // asn fpx11114__overflow_bit_count__13987, %left_shift(__tid1996__13985, 3<uint<64>>)

assign __tid1567__13991 = fpx11114__overflow_bit_count__13987[7:0]; // asn __tid1567__13991, %bit_read(fpx11114__overflow_bit_count__13987, 7<uint<4>>, 0<uint<1>>)

assign __tid1573__13993 = fpx11114__overflow_bit_count__13987; // asn __tid1573__13993, fpx11114__overflow_bit_count__13987

assign __tid1579__13995 = __tid1573__13993 > 64'd0; // asn __tid1579__13995, %greater_than(__tid1573__13993, 0<uint<64>>)

assign __tid1581__13996 = __tid1579__13995; // asn __tid1581__13996, __tid1579__13995

assign __tid1720__14009 = __tid9701__13202; // asn __tid1720__14009, __tid9701__13202

assign __tid1724__14011 = __tid1720__14009 == 3'd0; // asn __tid1724__14011, %is_equal(__tid1720__14009, 0<uint<3>>)

assign __tid1734__14012 = ! __tid1724__14011; // asn __tid1734__14012, %logical_not(__tid1724__14011)

assign __tid1726__14015 = __tid9701__13202; // asn __tid1726__14015, __tid9701__13202

assign __tid1730__14018 = __tid1726__14015 == 3'd4; // asn __tid1730__14018, %is_equal(__tid1726__14015, 4<uint<3>>)

assign __tid1730__14024 = (__tid1734__14012) ? __tid1730__14018 : __tid1730__13890;

assign __tid1740__14025 = __tid1724__14011 | __tid1730__14024; // asn __tid1740__14025, %logical_or(__tid1724__14011, __tid1730__14024)

assign __tid1742__14026 = __tid1740__14025; // asn __tid1742__14026, __tid1740__14025

assign __tid1752__14031 = __tid9701__13202; // asn __tid1752__14031, __tid9701__13202

assign __tid1756__14033 = __tid1752__14031 == 3'd1; // asn __tid1756__14033, %is_equal(__tid1752__14031, 1<uint<3>>)

assign __tid1766__14034 = ! __tid1756__14033; // asn __tid1766__14034, %logical_not(__tid1756__14033)

assign __tid1758__14037 = __tid9701__13202; // asn __tid1758__14037, __tid9701__13202

assign __tid1762__14040 = { 1'd0, __tid1758__14037 } == 4'd5; // asn __tid1762__14040, %is_equal(__tid1758__14037, 5<uint<4>>)

assign __tid1762__14046 = (__tid1766__14034) ? __tid1762__14040 : __tid1762__13912;

assign __tid1772__14047 = __tid1756__14033 | __tid1762__14046; // asn __tid1772__14047, %logical_or(__tid1756__14033, __tid1762__14046)

assign __tid1774__14048 = __tid1772__14047; // asn __tid1774__14048, __tid1772__14047

assign __tid1784__14053 = __tid9701__13202; // asn __tid1784__14053, __tid9701__13202

assign __tid1788__14055 = __tid1784__14053 == 3'd2; // asn __tid1788__14055, %is_equal(__tid1784__14053, 2<uint<3>>)

assign __tid1798__14056 = ! __tid1788__14055; // asn __tid1798__14056, %logical_not(__tid1788__14055)

assign __tid1790__14059 = __tid9701__13202; // asn __tid1790__14059, __tid9701__13202

assign __tid1794__14062 = { 1'd0, __tid1790__14059 } == 4'd6; // asn __tid1794__14062, %is_equal(__tid1790__14059, 6<uint<4>>)

assign __tid1794__14068 = (__tid1798__14056) ? __tid1794__14062 : __tid1794__13934;

assign __tid1804__14069 = __tid1788__14055 | __tid1794__14068; // asn __tid1804__14069, %logical_or(__tid1788__14055, __tid1794__14068)

assign __tid1806__14070 = __tid1804__14069; // asn __tid1806__14070, __tid1804__14069

assign __tid1808__14071 = ! __tid1742__14026; // asn __tid1808__14071, %logical_not(__tid1742__14026)

assign __tid1810__14072 = __tid1808__14071 & __tid1774__14048; // asn __tid1810__14072, %logical_and(__tid1808__14071, __tid1774__14048)

assign __tid1812__14073 = ! __tid1810__14072; // asn __tid1812__14073, %logical_not(__tid1810__14072)

assign __tid1814__14074 = __tid1812__14073 & __tid1806__14070; // asn __tid1814__14074, %logical_and(__tid1812__14073, __tid1806__14070)

assign __tid1810__14077 = __tid1810__14072; // asn __tid1810__14077, __tid1810__14072

assign __tid1814__14080 = __tid1814__14074; // asn __tid1814__14080, __tid1814__14074

assign fpx11437__rtrn__14084 = (__tid1814__14080) ? fpx11437__rtrn__14082 : fpx11437__rtrn__14004;

assign fpx11437__rtrn__14085 = (__tid1810__14077) ? fpx11437__rtrn__14079 : fpx11437__rtrn__14084;

assign fpx11437__rtrn__14086 = (__tid1742__14026) ? fpx11437__rtrn__14076 : fpx11437__rtrn__14085;

assign __tid1599__14093 = fpx11437__rtrn__14086; // asn __tid1599__14093, fpx11437__rtrn__14086

assign __tid1601__14094 = 8'd8 - __tid1599__14093; // asn __tid1601__14094, %subtraction(8<uint<8>>, __tid1599__14093)

assign __tid1605__14096 = __tid1601__14094 << 8'd3; // asn __tid1605__14096, %left_shift(__tid1601__14094, 3<uint<8>>)

assign __tid1607__14098 = __tid1567__13991; // asn __tid1607__14098, __tid1567__13991

assign fpx11114__to_shift_off__14099 = __tid1605__14096 + __tid1607__14098; // asn fpx11114__to_shift_off__14099, %addition(__tid1605__14096, __tid1607__14098)

assign __tid1615__14101 = fpx11347__data__13830; // asn __tid1615__14101, fpx11347__data__13830

assign __tid1617__14102 = fpx11114__to_shift_off__14099; // asn __tid1617__14102, fpx11114__to_shift_off__14099

assign __tid1619__14103 = __tid1615__14101 << __tid1617__14102; // asn __tid1619__14103, %left_shift(__tid1615__14101, __tid1617__14102)

assign __tid1621__14104 = fpx11114__to_shift_off__14099; // asn __tid1621__14104, fpx11114__to_shift_off__14099

assign fpx11114__rtrn__14105 = __tid1619__14103 >> __tid1621__14104; // asn fpx11114__rtrn__14105, %right_shift(__tid1619__14103, __tid1621__14104)

assign __tid1730__14119 = (__tid1581__13996) ? __tid1730__14024 : __tid1730__13890;

assign __tid1762__14130 = (__tid1581__13996) ? __tid1762__14046 : __tid1762__13912;

assign __tid1794__14141 = (__tid1581__13996) ? __tid1794__14068 : __tid1794__13934;

assign fpx11114__rtrn__14176 = (__tid1581__13996) ? fpx11114__rtrn__14105 : fpx11347__data__13830;

assign fpx10696__data_low__14177 = fpx11114__rtrn__14176; // asn fpx10696__data_low__14177, fpx11114__rtrn__14176

assign fpx10696__data_low__14183 = fpx10696__data_low__14177 << fpx10696__low_bit_count__14182; // asn fpx10696__data_low__14183, %left_shift(fpx10696__data_low__14177, fpx10696__low_bit_count__14182)

assign __tid1355__14199 = fpx10696__data_low__14183; // asn __tid1355__14199, fpx10696__data_low__14183

assign fpx10696__write_val__14201 = __tid1355__14199 | __tid1357__14200; // asn fpx10696__write_val__14201, %numeric_or(__tid1355__14199, __tid1357__14200)

assign __tid1720__14220 = __tid9701__13202; // asn __tid1720__14220, __tid9701__13202

assign __tid1724__14222 = __tid1720__14220 == 3'd0; // asn __tid1724__14222, %is_equal(__tid1720__14220, 0<uint<3>>)

assign __tid1734__14223 = ! __tid1724__14222; // asn __tid1734__14223, %logical_not(__tid1724__14222)

assign __tid1726__14226 = __tid9701__13202; // asn __tid1726__14226, __tid9701__13202

assign __tid1730__14229 = __tid1726__14226 == 3'd4; // asn __tid1730__14229, %is_equal(__tid1726__14226, 4<uint<3>>)

assign __tid1730__14232 = (__tid1734__14223) ? __tid1730__14229 : __tid1730__14119;

assign __tid1740__14233 = __tid1724__14222 | __tid1730__14232; // asn __tid1740__14233, %logical_or(__tid1724__14222, __tid1730__14232)

assign __tid1742__14234 = __tid1740__14233; // asn __tid1742__14234, __tid1740__14233

assign __tid1752__14237 = __tid9701__13202; // asn __tid1752__14237, __tid9701__13202

assign __tid1756__14239 = __tid1752__14237 == 3'd1; // asn __tid1756__14239, %is_equal(__tid1752__14237, 1<uint<3>>)

assign __tid1766__14240 = ! __tid1756__14239; // asn __tid1766__14240, %logical_not(__tid1756__14239)

assign __tid1758__14243 = __tid9701__13202; // asn __tid1758__14243, __tid9701__13202

assign __tid1762__14246 = { 1'd0, __tid1758__14243 } == 4'd5; // asn __tid1762__14246, %is_equal(__tid1758__14243, 5<uint<4>>)

assign __tid1762__14249 = (__tid1766__14240) ? __tid1762__14246 : __tid1762__14130;

assign __tid1772__14250 = __tid1756__14239 | __tid1762__14249; // asn __tid1772__14250, %logical_or(__tid1756__14239, __tid1762__14249)

assign __tid1774__14251 = __tid1772__14250; // asn __tid1774__14251, __tid1772__14250

assign __tid1784__14254 = __tid9701__13202; // asn __tid1784__14254, __tid9701__13202

assign __tid1788__14256 = __tid1784__14254 == 3'd2; // asn __tid1788__14256, %is_equal(__tid1784__14254, 2<uint<3>>)

assign __tid1798__14257 = ! __tid1788__14256; // asn __tid1798__14257, %logical_not(__tid1788__14256)

assign __tid1790__14260 = __tid9701__13202; // asn __tid1790__14260, __tid9701__13202

assign __tid1794__14263 = { 1'd0, __tid1790__14260 } == 4'd6; // asn __tid1794__14263, %is_equal(__tid1790__14260, 6<uint<4>>)

assign __tid1794__14266 = (__tid1798__14257) ? __tid1794__14263 : __tid1794__14141;

assign __tid1804__14267 = __tid1788__14256 | __tid1794__14266; // asn __tid1804__14267, %logical_or(__tid1788__14256, __tid1794__14266)

assign __tid1806__14268 = __tid1804__14267; // asn __tid1806__14268, __tid1804__14267

assign __tid1808__14269 = ! __tid1742__14234; // asn __tid1808__14269, %logical_not(__tid1742__14234)

assign __tid1810__14270 = __tid1808__14269 & __tid1774__14251; // asn __tid1810__14270, %logical_and(__tid1808__14269, __tid1774__14251)

assign __tid1812__14271 = ! __tid1810__14270; // asn __tid1812__14271, %logical_not(__tid1810__14270)

assign __tid1814__14272 = __tid1812__14271 & __tid1806__14268; // asn __tid1814__14272, %logical_and(__tid1812__14271, __tid1806__14268)

assign __tid1810__14275 = __tid1810__14270; // asn __tid1810__14275, __tid1810__14270

assign __tid1814__14278 = __tid1814__14272; // asn __tid1814__14278, __tid1814__14272

assign fpx11496__rtrn__14282 = (__tid1814__14278) ? fpx11496__rtrn__14280 : fpx11496__rtrn__14217;

assign fpx11496__rtrn__14283 = (__tid1810__14275) ? fpx11496__rtrn__14277 : fpx11496__rtrn__14282;

assign fpx11496__rtrn__14284 = (__tid1742__14234) ? fpx11496__rtrn__14274 : fpx11496__rtrn__14283;

assign __tid1874__14287 = fpx11496__rtrn__14284; // asn __tid1874__14287, fpx11496__rtrn__14284

assign fpx11145__needed__14288 = __tid1872__14286 + { 56'd0, __tid1874__14287 }; // asn fpx11145__needed__14288, %addition(__tid1872__14286, __tid1874__14287)

assign __tid1886__14291 = fpx11145__needed__14288; // asn __tid1886__14291, fpx11145__needed__14288

assign __tid1892__14293 = __tid1886__14291 < 64'd8; // asn __tid1892__14293, %less_than(__tid1886__14291, 8<uint<64>>)

assign __tid1894__14294 = __tid1892__14293; // asn __tid1894__14294, __tid1892__14293

assign __tid1902__14300 = fpx11145__needed__14288; // asn __tid1902__14300, fpx11145__needed__14288

assign fpx11145__rtrn__14301 = 64'd8 - __tid1902__14300; // asn fpx11145__rtrn__14301, %subtraction(8<uint<64>>, __tid1902__14300)

assign fpx11145__rtrn__14308 = (__tid1894__14294) ? fpx11145__rtrn__14301 : fpx11145__rtrn__14289;

assign __tid1915__14310 = fpx11145__rtrn__14308; // asn __tid1915__14310, fpx11145__rtrn__14308

assign fpx10696__high_bit_count__14312 = __tid1915__14310 << 64'd3; // asn fpx10696__high_bit_count__14312, %left_shift(__tid1915__14310, 3<uint<64>>)

assign __tid1372__14313 = fpx10696__high_bit_count__14312; // asn __tid1372__14313, fpx10696__high_bit_count__14312

assign __tid1378__14315 = __tid1372__14313 == 64'd0; // asn __tid1378__14315, %is_equal(__tid1372__14313, 0<uint<64>>)

assign __tid1380__14316 = __tid1378__14315; // asn __tid1380__14316, __tid1378__14315

assign __tid1720__14336 = __tid9701__13202; // asn __tid1720__14336, __tid9701__13202

assign __tid1724__14338 = __tid1720__14336 == 3'd0; // asn __tid1724__14338, %is_equal(__tid1720__14336, 0<uint<3>>)

assign __tid1734__14339 = ! __tid1724__14338; // asn __tid1734__14339, %logical_not(__tid1724__14338)

assign __tid1726__14342 = __tid9701__13202; // asn __tid1726__14342, __tid9701__13202

assign __tid1730__14345 = __tid1726__14342 == 3'd4; // asn __tid1730__14345, %is_equal(__tid1726__14342, 4<uint<3>>)

assign __tid1730__14351 = (__tid1734__14339) ? __tid1730__14345 : __tid1730__14232;

assign __tid1740__14352 = __tid1724__14338 | __tid1730__14351; // asn __tid1740__14352, %logical_or(__tid1724__14338, __tid1730__14351)

assign __tid1742__14353 = __tid1740__14352; // asn __tid1742__14353, __tid1740__14352

assign __tid1752__14358 = __tid9701__13202; // asn __tid1752__14358, __tid9701__13202

assign __tid1756__14360 = __tid1752__14358 == 3'd1; // asn __tid1756__14360, %is_equal(__tid1752__14358, 1<uint<3>>)

assign __tid1766__14361 = ! __tid1756__14360; // asn __tid1766__14361, %logical_not(__tid1756__14360)

assign __tid1758__14364 = __tid9701__13202; // asn __tid1758__14364, __tid9701__13202

assign __tid1762__14367 = { 1'd0, __tid1758__14364 } == 4'd5; // asn __tid1762__14367, %is_equal(__tid1758__14364, 5<uint<4>>)

assign __tid1762__14373 = (__tid1766__14361) ? __tid1762__14367 : __tid1762__14249;

assign __tid1772__14374 = __tid1756__14360 | __tid1762__14373; // asn __tid1772__14374, %logical_or(__tid1756__14360, __tid1762__14373)

assign __tid1774__14375 = __tid1772__14374; // asn __tid1774__14375, __tid1772__14374

assign __tid1784__14380 = __tid9701__13202; // asn __tid1784__14380, __tid9701__13202

assign __tid1788__14382 = __tid1784__14380 == 3'd2; // asn __tid1788__14382, %is_equal(__tid1784__14380, 2<uint<3>>)

assign __tid1798__14383 = ! __tid1788__14382; // asn __tid1798__14383, %logical_not(__tid1788__14382)

assign __tid1790__14386 = __tid9701__13202; // asn __tid1790__14386, __tid9701__13202

assign __tid1794__14389 = { 1'd0, __tid1790__14386 } == 4'd6; // asn __tid1794__14389, %is_equal(__tid1790__14386, 6<uint<4>>)

assign __tid1794__14395 = (__tid1798__14383) ? __tid1794__14389 : __tid1794__14266;

assign __tid1804__14396 = __tid1788__14382 | __tid1794__14395; // asn __tid1804__14396, %logical_or(__tid1788__14382, __tid1794__14395)

assign __tid1806__14397 = __tid1804__14396; // asn __tid1806__14397, __tid1804__14396

assign __tid1808__14398 = ! __tid1742__14353; // asn __tid1808__14398, %logical_not(__tid1742__14353)

assign __tid1810__14399 = __tid1808__14398 & __tid1774__14375; // asn __tid1810__14399, %logical_and(__tid1808__14398, __tid1774__14375)

assign __tid1812__14400 = ! __tid1810__14399; // asn __tid1812__14400, %logical_not(__tid1810__14399)

assign __tid1814__14401 = __tid1812__14400 & __tid1806__14397; // asn __tid1814__14401, %logical_and(__tid1812__14400, __tid1806__14397)

assign __tid1810__14404 = __tid1810__14399; // asn __tid1810__14404, __tid1810__14399

assign __tid1814__14407 = __tid1814__14401; // asn __tid1814__14407, __tid1814__14401

assign fpx11555__rtrn__14411 = (__tid1814__14407) ? fpx11555__rtrn__14409 : fpx11555__rtrn__14331;

assign fpx11555__rtrn__14412 = (__tid1810__14404) ? fpx11555__rtrn__14406 : fpx11555__rtrn__14411;

assign fpx11555__rtrn__14413 = (__tid1742__14353) ? fpx11555__rtrn__14403 : fpx11555__rtrn__14412;

assign __tid1955__14421 = fpx11555__rtrn__14413; // asn __tid1955__14421, fpx11555__rtrn__14413

assign fpx11175__needed__14422 = __tid1953__14420 + { 56'd0, __tid1955__14421 }; // asn fpx11175__needed__14422, %addition(__tid1953__14420, __tid1955__14421)

assign __tid1967__14426 = fpx11175__needed__14422; // asn __tid1967__14426, fpx11175__needed__14422

assign __tid1973__14428 = __tid1967__14426 > 64'd8; // asn __tid1973__14428, %greater_than(__tid1967__14426, 8<uint<64>>)

assign __tid1975__14429 = __tid1973__14428; // asn __tid1975__14429, __tid1973__14428

assign __tid1981__14434 = fpx11175__needed__14422; // asn __tid1981__14434, fpx11175__needed__14422

assign fpx11175__rtrn__14436 = __tid1981__14434 - 64'd8; // asn fpx11175__rtrn__14436, %subtraction(__tid1981__14434, 8<uint<64>>)

assign fpx11175__rtrn__14443 = (__tid1975__14429) ? fpx11175__rtrn__14436 : fpx11175__rtrn__14423;

assign __tid1996__14446 = fpx11175__rtrn__14443; // asn __tid1996__14446, fpx11175__rtrn__14443

assign fpx10696__overflow_bit_count__14448 = __tid1996__14446 << 64'd3; // asn fpx10696__overflow_bit_count__14448, %left_shift(__tid1996__14446, 3<uint<64>>)

assign __tid1392__14449 = fpx10696__overflow_bit_count__14448; // asn __tid1392__14449, fpx10696__overflow_bit_count__14448

assign __tid1398__14451 = __tid1392__14449 > 64'd0; // asn __tid1398__14451, %greater_than(__tid1392__14449, 0<uint<64>>)

assign __tid1400__14452 = __tid1398__14451; // asn __tid1400__14452, __tid1398__14451

assign __tid1720__14477 = __tid9701__13202; // asn __tid1720__14477, __tid9701__13202

assign __tid1724__14479 = __tid1720__14477 == 3'd0; // asn __tid1724__14479, %is_equal(__tid1720__14477, 0<uint<3>>)

assign __tid1734__14480 = ! __tid1724__14479; // asn __tid1734__14480, %logical_not(__tid1724__14479)

assign __tid1726__14483 = __tid9701__13202; // asn __tid1726__14483, __tid9701__13202

assign __tid1730__14486 = __tid1726__14483 == 3'd4; // asn __tid1730__14486, %is_equal(__tid1726__14483, 4<uint<3>>)

assign __tid1730__14492 = (__tid1734__14480) ? __tid1730__14486 : __tid1730__14351;

assign __tid1740__14493 = __tid1724__14479 | __tid1730__14492; // asn __tid1740__14493, %logical_or(__tid1724__14479, __tid1730__14492)

assign __tid1742__14494 = __tid1740__14493; // asn __tid1742__14494, __tid1740__14493

assign __tid1752__14499 = __tid9701__13202; // asn __tid1752__14499, __tid9701__13202

assign __tid1756__14501 = __tid1752__14499 == 3'd1; // asn __tid1756__14501, %is_equal(__tid1752__14499, 1<uint<3>>)

assign __tid1766__14502 = ! __tid1756__14501; // asn __tid1766__14502, %logical_not(__tid1756__14501)

assign __tid1758__14505 = __tid9701__13202; // asn __tid1758__14505, __tid9701__13202

assign __tid1762__14508 = { 1'd0, __tid1758__14505 } == 4'd5; // asn __tid1762__14508, %is_equal(__tid1758__14505, 5<uint<4>>)

assign __tid1762__14514 = (__tid1766__14502) ? __tid1762__14508 : __tid1762__14373;

assign __tid1772__14515 = __tid1756__14501 | __tid1762__14514; // asn __tid1772__14515, %logical_or(__tid1756__14501, __tid1762__14514)

assign __tid1774__14516 = __tid1772__14515; // asn __tid1774__14516, __tid1772__14515

assign __tid1784__14521 = __tid9701__13202; // asn __tid1784__14521, __tid9701__13202

assign __tid1788__14523 = __tid1784__14521 == 3'd2; // asn __tid1788__14523, %is_equal(__tid1784__14521, 2<uint<3>>)

assign __tid1798__14524 = ! __tid1788__14523; // asn __tid1798__14524, %logical_not(__tid1788__14523)

assign __tid1790__14527 = __tid9701__13202; // asn __tid1790__14527, __tid9701__13202

assign __tid1794__14530 = { 1'd0, __tid1790__14527 } == 4'd6; // asn __tid1794__14530, %is_equal(__tid1790__14527, 6<uint<4>>)

assign __tid1794__14536 = (__tid1798__14524) ? __tid1794__14530 : __tid1794__14395;

assign __tid1804__14537 = __tid1788__14523 | __tid1794__14536; // asn __tid1804__14537, %logical_or(__tid1788__14523, __tid1794__14536)

assign __tid1806__14538 = __tid1804__14537; // asn __tid1806__14538, __tid1804__14537

assign __tid1808__14539 = ! __tid1742__14494; // asn __tid1808__14539, %logical_not(__tid1742__14494)

assign __tid1810__14540 = __tid1808__14539 & __tid1774__14516; // asn __tid1810__14540, %logical_and(__tid1808__14539, __tid1774__14516)

assign __tid1812__14541 = ! __tid1810__14540; // asn __tid1812__14541, %logical_not(__tid1810__14540)

assign __tid1814__14542 = __tid1812__14541 & __tid1806__14538; // asn __tid1814__14542, %logical_and(__tid1812__14541, __tid1806__14538)

assign __tid1810__14545 = __tid1810__14540; // asn __tid1810__14545, __tid1810__14540

assign __tid1814__14548 = __tid1814__14542; // asn __tid1814__14548, __tid1814__14542

assign fpx11614__rtrn__14552 = (__tid1814__14548) ? fpx11614__rtrn__14550 : fpx11614__rtrn__14472;

assign fpx11614__rtrn__14553 = (__tid1810__14545) ? fpx11614__rtrn__14547 : fpx11614__rtrn__14552;

assign fpx11614__rtrn__14554 = (__tid1742__14494) ? fpx11614__rtrn__14544 : fpx11614__rtrn__14553;

assign __tid1665__14558 = fpx11614__rtrn__14554; // asn __tid1665__14558, fpx11614__rtrn__14554

assign fpx11194__access_width_bits__14560 = __tid1665__14558 << 8'd3; // asn fpx11194__access_width_bits__14560, %left_shift(__tid1665__14558, 3<uint<8>>)

assign __tid1720__14577 = __tid9701__13202; // asn __tid1720__14577, __tid9701__13202

assign __tid1724__14579 = __tid1720__14577 == 3'd0; // asn __tid1724__14579, %is_equal(__tid1720__14577, 0<uint<3>>)

assign __tid1734__14580 = ! __tid1724__14579; // asn __tid1734__14580, %logical_not(__tid1724__14579)

assign __tid1726__14583 = __tid9701__13202; // asn __tid1726__14583, __tid9701__13202

assign __tid1730__14586 = __tid1726__14583 == 3'd4; // asn __tid1730__14586, %is_equal(__tid1726__14583, 4<uint<3>>)

assign __tid1730__14589 = (__tid1734__14580) ? __tid1730__14586 : __tid1730__14492;

assign __tid1740__14590 = __tid1724__14579 | __tid1730__14589; // asn __tid1740__14590, %logical_or(__tid1724__14579, __tid1730__14589)

assign __tid1742__14591 = __tid1740__14590; // asn __tid1742__14591, __tid1740__14590

assign __tid1752__14596 = __tid9701__13202; // asn __tid1752__14596, __tid9701__13202

assign __tid1756__14598 = __tid1752__14596 == 3'd1; // asn __tid1756__14598, %is_equal(__tid1752__14596, 1<uint<3>>)

assign __tid1766__14599 = ! __tid1756__14598; // asn __tid1766__14599, %logical_not(__tid1756__14598)

assign __tid1758__14602 = __tid9701__13202; // asn __tid1758__14602, __tid9701__13202

assign __tid1762__14605 = { 1'd0, __tid1758__14602 } == 4'd5; // asn __tid1762__14605, %is_equal(__tid1758__14602, 5<uint<4>>)

assign __tid1762__14608 = (__tid1766__14599) ? __tid1762__14605 : __tid1762__14514;

assign __tid1772__14609 = __tid1756__14598 | __tid1762__14608; // asn __tid1772__14609, %logical_or(__tid1756__14598, __tid1762__14608)

assign __tid1774__14610 = __tid1772__14609; // asn __tid1774__14610, __tid1772__14609

assign __tid1784__14615 = __tid9701__13202; // asn __tid1784__14615, __tid9701__13202

assign __tid1788__14617 = __tid1784__14615 == 3'd2; // asn __tid1788__14617, %is_equal(__tid1784__14615, 2<uint<3>>)

assign __tid1798__14618 = ! __tid1788__14617; // asn __tid1798__14618, %logical_not(__tid1788__14617)

assign __tid1790__14621 = __tid9701__13202; // asn __tid1790__14621, __tid9701__13202

assign __tid1794__14624 = { 1'd0, __tid1790__14621 } == 4'd6; // asn __tid1794__14624, %is_equal(__tid1790__14621, 6<uint<4>>)

assign __tid1794__14627 = (__tid1798__14618) ? __tid1794__14624 : __tid1794__14536;

assign __tid1804__14628 = __tid1788__14617 | __tid1794__14627; // asn __tid1804__14628, %logical_or(__tid1788__14617, __tid1794__14627)

assign __tid1806__14629 = __tid1804__14628; // asn __tid1806__14629, __tid1804__14628

assign __tid1808__14630 = ! __tid1742__14591; // asn __tid1808__14630, %logical_not(__tid1742__14591)

assign __tid1810__14631 = __tid1808__14630 & __tid1774__14610; // asn __tid1810__14631, %logical_and(__tid1808__14630, __tid1774__14610)

assign __tid1812__14632 = ! __tid1810__14631; // asn __tid1812__14632, %logical_not(__tid1810__14631)

assign __tid1814__14633 = __tid1812__14632 & __tid1806__14629; // asn __tid1814__14633, %logical_and(__tid1812__14632, __tid1806__14629)

assign __tid1810__14636 = __tid1810__14631; // asn __tid1810__14636, __tid1810__14631

assign __tid1814__14639 = __tid1814__14633; // asn __tid1814__14639, __tid1814__14633

assign fpx11762__rtrn__14643 = (__tid1814__14639) ? fpx11762__rtrn__14641 : fpx11762__rtrn__14572;

assign fpx11762__rtrn__14644 = (__tid1810__14636) ? fpx11762__rtrn__14638 : fpx11762__rtrn__14643;

assign fpx11762__rtrn__14645 = (__tid1742__14591) ? fpx11762__rtrn__14635 : fpx11762__rtrn__14644;

assign __tid1955__14653 = fpx11762__rtrn__14645; // asn __tid1955__14653, fpx11762__rtrn__14645

assign fpx11643__needed__14654 = __tid1953__14652 + { 56'd0, __tid1955__14653 }; // asn fpx11643__needed__14654, %addition(__tid1953__14652, __tid1955__14653)

assign __tid1967__14658 = fpx11643__needed__14654; // asn __tid1967__14658, fpx11643__needed__14654

assign __tid1973__14660 = __tid1967__14658 > 64'd8; // asn __tid1973__14660, %greater_than(__tid1967__14658, 8<uint<64>>)

assign __tid1975__14661 = __tid1973__14660; // asn __tid1975__14661, __tid1973__14660

assign __tid1981__14666 = fpx11643__needed__14654; // asn __tid1981__14666, fpx11643__needed__14654

assign fpx11643__rtrn__14668 = __tid1981__14666 - 64'd8; // asn fpx11643__rtrn__14668, %subtraction(__tid1981__14666, 8<uint<64>>)

assign fpx11643__rtrn__14675 = (__tid1975__14661) ? fpx11643__rtrn__14668 : fpx11643__rtrn__14655;

assign __tid1996__14678 = fpx11643__rtrn__14675; // asn __tid1996__14678, fpx11643__rtrn__14675

assign fpx11194__overflow_bits__14680 = __tid1996__14678 << 64'd3; // asn fpx11194__overflow_bits__14680, %left_shift(__tid1996__14678, 3<uint<64>>)

assign __tid1683__14681 = fpx11194__access_width_bits__14560; // asn __tid1683__14681, fpx11194__access_width_bits__14560

assign __tid1685__14682 = fpx11194__overflow_bits__14680; // asn __tid1685__14682, fpx11194__overflow_bits__14680

assign fpx11194__to_shift_off__14683 = { 56'd0, __tid1683__14681 } - __tid1685__14682; // asn fpx11194__to_shift_off__14683, %subtraction(__tid1683__14681, __tid1685__14682)

assign fpx11194__rtrn__14684 = fpx11194__rtrn__14466 >> fpx11194__to_shift_off__14683; // asn fpx11194__rtrn__14684, %right_shift(fpx11194__rtrn__14466, fpx11194__to_shift_off__14683)

assign __tid1434__14696 = fpx10696__overflow_bit_count__14448; // asn __tid1434__14696, fpx10696__overflow_bit_count__14448

assign __tid1436__14697 = __tid1432__14694 >> __tid1434__14696; // asn __tid1436__14697, %right_shift(__tid1432__14694, __tid1434__14696)

assign __tid1438__14699 = fpx10696__overflow_bit_count__14448; // asn __tid1438__14699, fpx10696__overflow_bit_count__14448

assign fpx10696__high_bits__14700 = __tid1436__14697 << __tid1438__14699; // asn fpx10696__high_bits__14700, %left_shift(__tid1436__14697, __tid1438__14699)

assign __tid1445__14701 = fpx10696__high_bits__14700; // asn __tid1445__14701, fpx10696__high_bits__14700

assign __tid1447__14702 = fpx11194__rtrn__14684; // asn __tid1447__14702, fpx11194__rtrn__14684

assign fpx10696__write_overflow_val__14703 = __tid1445__14701 | __tid1447__14702; // asn fpx10696__write_overflow_val__14703, %numeric_or(__tid1445__14701, __tid1447__14702)

assign fpx10696__write_overflow_val__14834 = (__tid1400__14452) ? fpx10696__write_overflow_val__14703 : fpx10696__write_overflow_val__14833;

assign __tid1467__14841 = fpx10696__high_bit_count__14312; // asn __tid1467__14841, fpx10696__high_bit_count__14312

assign fpx10696__to_shift_out__14842 = 64'd64 - __tid1467__14841; // asn fpx10696__to_shift_out__14842, %subtraction(64<uint<64>>, __tid1467__14841)

assign __tid1477__14845 = fpx10696__to_shift_out__14842; // asn __tid1477__14845, fpx10696__to_shift_out__14842

assign __tid1479__14846 = __tid1475__14844 >> __tid1477__14845; // asn __tid1479__14846, %right_shift(__tid1475__14844, __tid1477__14845)

assign __tid1481__14847 = fpx10696__to_shift_out__14842; // asn __tid1481__14847, fpx10696__to_shift_out__14842

assign fpx10696__high_bits__14848 = __tid1479__14846 << __tid1481__14847; // asn fpx10696__high_bits__14848, %left_shift(__tid1479__14846, __tid1481__14847)

assign fpx10696__write_val__14849 = fpx10696__write_val__14201; // asn fpx10696__write_val__14849, fpx10696__write_val__14201

assign fpx10696__write_val__14850 = fpx10696__write_val__14849 | fpx10696__high_bits__14848; // asn fpx10696__write_val__14850, %numeric_or(fpx10696__write_val__14849, fpx10696__high_bits__14848)

assign fpx10696__write_overflow_val__14978 = (__tid1380__14316) ? fpx10696__write_overflow_val__14834 : fpx10696__write_overflow_val__14833;

assign fpx10696__has_overflow__14979 = (__tid1380__14316) ? __tid1398__14451 : fpx10696__has_overflow__14835;

assign fpx10696__write_val__14995 = (__tid1380__14316) ? fpx10696__write_val__14201 : fpx10696__write_val__14850;

assign fpx10696__write_val__15006 = (__tid1177__13251) ? fpx10696__write_val__13508 : fpx10696__write_val__14995;

assign fpx10696__write_overflow_val__15405 = (__tid1177__13251) ? fpx10696__write_overflow_val__13246 : fpx10696__write_overflow_val__14978;

assign fpx10696__has_overflow__15406 = (__tid1177__13251) ? fpx10696__has_overflow__13247 : fpx10696__has_overflow__14979;

assign __tid1505__15417 = fpx10696__has_overflow__15406; // asn __tid1505__15417, fpx10696__has_overflow__15406

assign raddr__read__15801 = (__tid9587__12100) ? raddr__read__13187 : __tid9591__12063;

assign rdata__read__15806 = (__tid9587__12100) ? rdata__read__12110 : __tid9591__12063;

assign dcache__write__16282 = (__tid9587__12100) ? dcache__write__15790 : __tid9591__12063;

assign decode_reg_addr__write__16288 = (__tid9583__12069) ? decode_reg_addr__write__12073 : __tid9587__12061;

assign raddr__read__16289 = (__tid9583__12069) ? raddr__read__12082 : raddr__read__15801;

assign decode_reg_data__16290 = (__tid9583__12069) ? rdata_pyri : fpx10559__result__12991;

assign decode_reg_data__write__16291 = (__tid9583__12069) ? decode_reg_data__write__12077 : __tid9587__12061;

assign rdata__read__16292 = (__tid9583__12069) ? rdata__read__12086 : rdata__read__15806;

assign debug_reg_addr__write__16294 = (__tid9583__12069) ? debug_reg_addr__write__12081 : __tid9587__12061;

assign debug_reg_data__16295 = (__tid9583__12069) ? rdata_pyri : fpx10559__result__12991;

assign debug_reg_data__write__16296 = (__tid9583__12069) ? debug_reg_data__write__12085 : __tid9587__12061;

assign branch_pc__write__16302 = (__tid9583__12069) ? branch_pc_valid_pyri : branch_pc__write__12096;

assign branch_pc__read__16303 = (__tid9583__12069) ? branch_pc_valid_pyri : branch_pc__read__12098;

assign dcache__write__16750 = (__tid9583__12069) ? dcache__write__15790 : dcache__write__16282;

assign branch_pc__write__16756 = (__tid9524__11865) ? branch_pc__write__12067 : branch_pc__write__16302;

assign branch_pc__read__16757 = (__tid9524__11865) ? branch_pc__read__12068 : branch_pc__read__16303;

assign decode_reg_addr__write__16759 = (__tid9524__11865) ? decode_reg_addr__write__11817 : decode_reg_addr__write__16288;

assign raddr__read__16760 = (__tid9524__11865) ? raddr__read__11822 : raddr__read__16289;

assign decode_reg_data_pyro = decode_reg_data__16290; // asn decode_reg_data_pyro, decode_reg_data__16290

assign decode_reg_data__write__16762 = (__tid9524__11865) ? decode_reg_data__write__11816 : decode_reg_data__write__16291;

assign rdata__read__16763 = (__tid9524__11865) ? rdata__read__11821 : rdata__read__16292;

assign debug_reg_addr__write__16766 = (__tid9524__11865) ? debug_reg_addr__write__11815 : debug_reg_addr__write__16294;

assign debug_reg_data_pyro = debug_reg_data__16295; // asn debug_reg_data_pyro, debug_reg_data__16295

assign debug_reg_data__write__16769 = (__tid9524__11865) ? debug_reg_data__write__11814 : debug_reg_data__write__16296;

assign dcache__write__17216 = (__tid9524__11865) ? dcache__write__11813 : dcache__write__16750;

assign dcache__write__17228 = dcache__write__17216; // asn dcache__write__17228, dcache__write__17216

assign debug_reg_data__write__17229 = debug_reg_data__write__16769; // asn debug_reg_data__write__17229, debug_reg_data__write__16769

assign debug_reg_addr__write__17230 = debug_reg_addr__write__16766; // asn debug_reg_addr__write__17230, debug_reg_addr__write__16766

assign decode_reg_data__write__17231 = decode_reg_data__write__16762; // asn decode_reg_data__write__17231, decode_reg_data__write__16762

assign decode_reg_addr__write__17232 = decode_reg_addr__write__16759; // asn decode_reg_addr__write__17232, decode_reg_addr__write__16759

assign branch_pc__write__17233 = branch_pc__write__16756; // asn branch_pc__write__17233, branch_pc__write__16756

assign rdata__read__17236 = rdata__read__16763; // asn rdata__read__17236, rdata__read__16763

assign raddr__read__17237 = raddr__read__16760; // asn raddr__read__17237, raddr__read__16760

assign branch_pc__read__17238 = branch_pc__read__16757; // asn branch_pc__read__17238, branch_pc__read__16757

assign __tid14924__17257 = ! branch_pc__read__17238; // asn __tid14924__17257, %logical_not(branch_pc__read__17238)

assign __tid14926__17258 = __tid14924__17257 | branch_pc_valid_pyri; // asn __tid14926__17258, %logical_or(__tid14924__17257, branch_pc_valid_pyri)

assign __tid14928__17259 = ! raddr__read__17237; // asn __tid14928__17259, %logical_not(raddr__read__17237)

assign __tid14930__17260 = __tid14928__17259 | raddr_valid_pyri; // asn __tid14930__17260, %logical_or(__tid14928__17259, raddr_valid_pyri)

assign __tid14932__17261 = ! rdata__read__17236; // asn __tid14932__17261, %logical_not(rdata__read__17236)

assign __tid14934__17262 = __tid14932__17261 | rdata_valid_pyri; // asn __tid14934__17262, %logical_or(__tid14932__17261, rdata_valid_pyri)

assign __tid14946__17268 = ! branch_pc__write__17233; // asn __tid14946__17268, %logical_not(branch_pc__write__17233)

assign __tid14950__17270 = __tid14946__17268 | __tid14948__17269; // asn __tid14950__17270, %logical_or(__tid14946__17268, __tid14948__17269)

assign __tid14952__17271 = ! decode_reg_addr__write__17232; // asn __tid14952__17271, %logical_not(decode_reg_addr__write__17232)

assign __tid14956__17273 = __tid14952__17271 | __tid14954__17272; // asn __tid14956__17273, %logical_or(__tid14952__17271, __tid14954__17272)

assign __tid14958__17274 = ! decode_reg_data__write__17231; // asn __tid14958__17274, %logical_not(decode_reg_data__write__17231)

assign __tid14962__17276 = __tid14958__17274 | __tid14960__17275; // asn __tid14962__17276, %logical_or(__tid14958__17274, __tid14960__17275)

assign __tid14964__17277 = ! debug_reg_addr__write__17230; // asn __tid14964__17277, %logical_not(debug_reg_addr__write__17230)

assign __tid14968__17279 = __tid14964__17277 | __tid14966__17278; // asn __tid14968__17279, %logical_or(__tid14964__17277, __tid14966__17278)

assign __tid14970__17280 = ! debug_reg_data__write__17229; // asn __tid14970__17280, %logical_not(debug_reg_data__write__17229)

assign __tid14974__17282 = __tid14970__17280 | __tid14972__17281; // asn __tid14974__17282, %logical_or(__tid14970__17280, __tid14972__17281)

assign __tid14983__17286 = __tid14922__17256 & __tid14926__17258; // asn __tid14983__17286, %logical_and(__tid14922__17256, __tid14926__17258)

assign __tid14985__17287 = __tid14983__17286 & __tid14930__17260; // asn __tid14985__17287, %logical_and(__tid14983__17286, __tid14930__17260)

assign __tid14987__17288 = __tid14985__17287 & __tid14934__17262; // asn __tid14987__17288, %logical_and(__tid14985__17287, __tid14934__17262)

assign __tid14989__17289 = __tid14987__17288 & __tid14938__17264; // asn __tid14989__17289, %logical_and(__tid14987__17288, __tid14938__17264)

assign __tid14991__17290 = __tid14989__17289 & __tid14944__17267; // asn __tid14991__17290, %logical_and(__tid14989__17289, __tid14944__17267)

assign __tid14993__17291 = __tid14991__17290 & __tid14950__17270; // asn __tid14993__17291, %logical_and(__tid14991__17290, __tid14950__17270)

assign __tid14995__17292 = __tid14993__17291 & __tid14956__17273; // asn __tid14995__17292, %logical_and(__tid14993__17291, __tid14956__17273)

assign __tid14997__17293 = __tid14995__17292 & __tid14962__17276; // asn __tid14997__17293, %logical_and(__tid14995__17292, __tid14962__17276)

assign __tid14999__17294 = __tid14997__17293 & __tid14968__17279; // asn __tid14999__17294, %logical_and(__tid14997__17293, __tid14968__17279)

assign __tid15001__17295 = __tid14999__17294 & __tid14974__17282; // asn __tid15001__17295, %logical_and(__tid14999__17294, __tid14974__17282)

assign __block_valid__17297 = __tid15001__17295; // asn __block_valid__17297, __tid15001__17295

assign __tid15012__17310 = ! __block_valid__17297; // asn __tid15012__17310, %logical_not(__block_valid__17297)

assign pc_valid_pyro = __tid15001__17295; // asn pc_valid_pyro, __tid15001__17295

assign branch_pc_valid_pyro = __block_valid__17297 & branch_pc__write__17233; // asn branch_pc_valid_pyro, %logical_and(__block_valid__17297, branch_pc__write__17233)

assign decode_reg_addr_valid_pyro = __block_valid__17297 & decode_reg_addr__write__17232; // asn decode_reg_addr_valid_pyro, %logical_and(__block_valid__17297, decode_reg_addr__write__17232)

assign decode_reg_data_valid_pyro = __block_valid__17297 & decode_reg_data__write__17231; // asn decode_reg_data_valid_pyro, %logical_and(__block_valid__17297, decode_reg_data__write__17231)

assign debug_reg_addr_valid_pyro = __block_valid__17297 & debug_reg_addr__write__17230; // asn debug_reg_addr_valid_pyro, %logical_and(__block_valid__17297, debug_reg_addr__write__17230)

assign debug_reg_data_valid_pyro = __block_valid__17297 & debug_reg_data__write__17229; // asn debug_reg_data_valid_pyro, %logical_and(__block_valid__17297, debug_reg_data__write__17229)

assign __tid15026__17317 = __block_valid__17297 & dcache__write__17228; // asn __tid15026__17317, %logical_and(__block_valid__17297, dcache__write__17228)

assign __tid15031__17320 = __tid15012__17310; // asn __tid15031__17320, __tid15012__17310

assign pc_retry_pyro = pc_valid_pyri & __tid15031__17320; // asn pc_retry_pyro, %logical_and(pc_valid_pyri, __tid15031__17320)

assign __tid15035__17322 = __tid15012__17310 | __tid14924__17257; // asn __tid15035__17322, %logical_or(__tid15012__17310, __tid14924__17257)

assign branch_pc_retry_pyro = branch_pc_valid_pyri & __tid15035__17322; // asn branch_pc_retry_pyro, %logical_and(branch_pc_valid_pyri, __tid15035__17322)

assign __tid15039__17324 = __tid15012__17310 | __tid14928__17259; // asn __tid15039__17324, %logical_or(__tid15012__17310, __tid14928__17259)

assign raddr_retry_pyro = raddr_valid_pyri & __tid15039__17324; // asn raddr_retry_pyro, %logical_and(raddr_valid_pyri, __tid15039__17324)

assign __tid15043__17326 = __tid15012__17310 | __tid14932__17261; // asn __tid15043__17326, %logical_or(__tid15012__17310, __tid14932__17261)

assign rdata_retry_pyro = rdata_valid_pyri & __tid15043__17326; // asn rdata_retry_pyro, %logical_and(rdata_valid_pyri, __tid15043__17326)

assign __tid15047__17328 = __tid15012__17310; // asn __tid15047__17328, __tid15012__17310

assign inst_retry_pyro = inst_valid_pyri & __tid15047__17328; // asn inst_retry_pyro, %logical_and(inst_valid_pyri, __tid15047__17328)

assign __tid17015__17376 = (__tid17013__17375) ? fpx10696__write_val__15006 : __tid17011__17374;

assign __tid17019__17378 = (__tid9591__13190) ? fpx10696__write_val__15006 : __tid17017__17377;

assign __tid17025__17381 = ! __tid9587__12100; // asn __tid17025__17381, %logical_not(__tid9587__12100)

assign __tid17029__17383 = (__tid17025__17381) ? __tid17019__17378 : __tid17027__17382;

assign __tid17035__17386 = ! __tid9583__12069; // asn __tid17035__17386, %logical_not(__tid9583__12069)

assign __tid17039__17388 = (__tid17035__17386) ? __tid17029__17383 : __tid17037__17387;

assign __tid17045__17391 = ! __tid9524__11865; // asn __tid17045__17391, %logical_not(__tid9524__11865)

assign __tid17049__17393 = (__tid17045__17391) ? __tid17039__17388 : __tid17047__17392;

assign __tid17057__17397 = (__tid15026__17317) ? __tid17049__17393 : __tid17055__17396;

assign __tid15978__17354 = (__tid1505__15417) ? fpx10696__write_overflow_val__15405 : __tid17015__17376;

assign __tid17023__17380 = (__tid9591__13190) ? __tid15978__17354 : __tid17021__17379;

assign __tid17033__17385 = (__tid17025__17381) ? __tid17023__17380 : __tid17031__17384;

assign __tid17043__17390 = (__tid17035__17386) ? __tid17033__17385 : __tid17041__17389;

assign __tid17053__17395 = (__tid17045__17391) ? __tid17043__17390 : __tid17051__17394;

assign __tid17061__17399 = (__tid15026__17317) ? __tid17053__17395 : __tid17059__17398;

assign __tid17237 = __tid17057__17397; // asn __tid17237, __tid17057__17397

assign __tid17239 = __tid17061__17399; // asn __tid17239, __tid17061__17399

write_back_block_dcache write_back_block_dcache_inst(.clk(clk), .__tid464__12131(__tid464__12131), .fpx10559__index__12128(fpx10559__index__12128), .__tid543__12464(__tid543__12464), .__tid541__12462(__tid541__12462), .__tid1203__13265(__tid1203__13265), .fpx10696__index__13264(fpx10696__index__13264), .__tid1323__14186(__tid1323__14186), .fpx10696__index__14185(fpx10696__index__14185), .__tid1424__14691(__tid1424__14691), .__tid1422__14689(__tid1422__14689), .__tid17011__17374(__tid17011__17374), .__tid1518__15422(__tid1518__15422), .__tid17017__17377(__tid17017__17377), .fpx10696__index__13244(fpx10696__index__13244), .__tid17021__17379(__tid17021__17379), .__tid17027__17382(__tid17027__17382), .__tid17031__17384(__tid17031__17384), .__tid17037__17387(__tid17037__17387), .__tid17041__17389(__tid17041__17389), .__tid17047__17392(__tid17047__17392), .__tid17051__17394(__tid17051__17394), .__tid17055__17396(__tid17055__17396), .__tid17059__17398(__tid17059__17398), .__tid17237(__tid17237), .__tid17239(__tid17239));





  always @(posedge clk) begin
    
  end




endmodule

/* verilator lint_on WIDTH */
