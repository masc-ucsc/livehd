// total modules: 2
// design tree depth: 2
// design size: 1119
// avg module size: 300
module Snxn1k (
  input  a,
  input  b,
  output z
);
  wire t0 = a + b;
  wire inv0  = ~t0;
  wire x0    = t0 ^ inv0;
  wire invx0 = ~x0;
  wire t1    = x0 + invx0;
  wire inv1  = ~t1;
  wire x1    = t1 ^ inv1;
  wire invx1 = ~x1;
  wire t2    = x1 + invx1;
  wire inv2  = ~t2;
  wire x2    = t2 ^ inv2;
  wire invx2 = ~x2;
  wire t3    = x2 + invx2;
  wire inv3  = ~t3;
  wire x3    = t3 ^ inv3;
  wire invx3 = ~x3;
  wire t4    = x3 + invx3;
  wire inv4  = ~t4;
  wire x4    = t4 ^ inv4;
  wire invx4 = ~x4;
  wire t5    = x4 + invx4;
  wire inv5  = ~t5;
  wire x5    = t5 ^ inv5;
  wire invx5 = ~x5;
  wire t6    = x5 + invx5;
  wire inv6  = ~t6;
  wire x6    = t6 ^ inv6;
  wire invx6 = ~x6;
  wire t7    = x6 + invx6;
  wire inv7  = ~t7;
  wire x7    = t7 ^ inv7;
  wire invx7 = ~x7;
  wire t8    = x7 + invx7;
  wire inv8  = ~t8;
  wire x8    = t8 ^ inv8;
  wire invx8 = ~x8;
  wire t9    = x8 + invx8;
  wire inv9  = ~t9;
  wire x9    = t9 ^ inv9;
  wire invx9 = ~x9;
  wire t10    = x9 + invx9;
  wire inv10  = ~t10;
  wire x10    = t10 ^ inv10;
  wire invx10 = ~x10;
  wire t11    = x10 + invx10;
  wire inv11  = ~t11;
  wire x11    = t11 ^ inv11;
  wire invx11 = ~x11;
  wire t12    = x11 + invx11;
  wire inv12  = ~t12;
  wire x12    = t12 ^ inv12;
  wire invx12 = ~x12;
  wire t13    = x12 + invx12;
  wire inv13  = ~t13;
  wire x13    = t13 ^ inv13;
  wire invx13 = ~x13;
  wire t14    = x13 + invx13;
  wire inv14  = ~t14;
  wire x14    = t14 ^ inv14;
  wire invx14 = ~x14;
  wire t15    = x14 + invx14;
  wire inv15  = ~t15;
  wire x15    = t15 ^ inv15;
  wire invx15 = ~x15;
  wire t16    = x15 + invx15;
  wire inv16  = ~t16;
  wire x16    = t16 ^ inv16;
  wire invx16 = ~x16;
  wire t17    = x16 + invx16;
  wire inv17  = ~t17;
  wire x17    = t17 ^ inv17;
  wire invx17 = ~x17;
  wire t18    = x17 + invx17;
  wire inv18  = ~t18;
  wire x18    = t18 ^ inv18;
  wire invx18 = ~x18;
  wire t19    = x18 + invx18;
  wire inv19  = ~t19;
  wire x19    = t19 ^ inv19;
  wire invx19 = ~x19;
  wire t20    = x19 + invx19;
  wire inv20  = ~t20;
  wire x20    = t20 ^ inv20;
  wire invx20 = ~x20;
  wire t21    = x20 + invx20;
  wire inv21  = ~t21;
  wire x21    = t21 ^ inv21;
  wire invx21 = ~x21;
  wire t22    = x21 + invx21;
  wire inv22  = ~t22;
  wire x22    = t22 ^ inv22;
  wire invx22 = ~x22;
  wire t23    = x22 + invx22;
  wire inv23  = ~t23;
  wire x23    = t23 ^ inv23;
  wire invx23 = ~x23;
  wire t24    = x23 + invx23;
  wire inv24  = ~t24;
  wire x24    = t24 ^ inv24;
  wire invx24 = ~x24;
  wire t25    = x24 + invx24;
  wire inv25  = ~t25;
  wire x25    = t25 ^ inv25;
  wire invx25 = ~x25;
  wire t26    = x25 + invx25;
  wire inv26  = ~t26;
  wire x26    = t26 ^ inv26;
  wire invx26 = ~x26;
  wire t27    = x26 + invx26;
  wire inv27  = ~t27;
  wire x27    = t27 ^ inv27;
  wire invx27 = ~x27;
  wire t28    = x27 + invx27;
  wire inv28  = ~t28;
  wire x28    = t28 ^ inv28;
  wire invx28 = ~x28;
  wire t29    = x28 + invx28;
  wire inv29  = ~t29;
  wire x29    = t29 ^ inv29;
  wire invx29 = ~x29;
  wire t30    = x29 + invx29;
  wire inv30  = ~t30;
  wire x30    = t30 ^ inv30;
  wire invx30 = ~x30;
  wire t31    = x30 + invx30;
  wire inv31  = ~t31;
  wire x31    = t31 ^ inv31;
  wire invx31 = ~x31;
  wire t32    = x31 + invx31;
  wire inv32  = ~t32;
  wire x32    = t32 ^ inv32;
  wire invx32 = ~x32;
  wire t33    = x32 + invx32;
  wire inv33  = ~t33;
  wire x33    = t33 ^ inv33;
  wire invx33 = ~x33;
  wire t34    = x33 + invx33;
  wire inv34  = ~t34;
  wire x34    = t34 ^ inv34;
  wire invx34 = ~x34;
  wire t35    = x34 + invx34;
  wire inv35  = ~t35;
  wire x35    = t35 ^ inv35;
  wire invx35 = ~x35;
  wire t36    = x35 + invx35;
  wire inv36  = ~t36;
  wire x36    = t36 ^ inv36;
  wire invx36 = ~x36;
  wire t37    = x36 + invx36;
  wire inv37  = ~t37;
  wire x37    = t37 ^ inv37;
  wire invx37 = ~x37;
  wire t38    = x37 + invx37;
  wire inv38  = ~t38;
  wire x38    = t38 ^ inv38;
  wire invx38 = ~x38;
  wire t39    = x38 + invx38;
  wire inv39  = ~t39;
  wire x39    = t39 ^ inv39;
  wire invx39 = ~x39;
  wire t40    = x39 + invx39;
  wire inv40  = ~t40;
  wire x40    = t40 ^ inv40;
  wire invx40 = ~x40;
  wire t41    = x40 + invx40;
  wire inv41  = ~t41;
  wire x41    = t41 ^ inv41;
  wire invx41 = ~x41;
  wire t42    = x41 + invx41;
  wire inv42  = ~t42;
  wire x42    = t42 ^ inv42;
  wire invx42 = ~x42;
  wire t43    = x42 + invx42;
  wire inv43  = ~t43;
  wire x43    = t43 ^ inv43;
  wire invx43 = ~x43;
  wire t44    = x43 + invx43;
  wire inv44  = ~t44;
  wire x44    = t44 ^ inv44;
  wire invx44 = ~x44;
  wire t45    = x44 + invx44;
  wire inv45  = ~t45;
  wire x45    = t45 ^ inv45;
  wire invx45 = ~x45;
  wire t46    = x45 + invx45;
  wire inv46  = ~t46;
  wire x46    = t46 ^ inv46;
  wire invx46 = ~x46;
  wire t47    = x46 + invx46;
  wire inv47  = ~t47;
  wire x47    = t47 ^ inv47;
  wire invx47 = ~x47;
  wire t48    = x47 + invx47;
  wire inv48  = ~t48;
  wire x48    = t48 ^ inv48;
  wire invx48 = ~x48;
  wire t49    = x48 + invx48;
  wire inv49  = ~t49;
  wire x49    = t49 ^ inv49;
  wire invx49 = ~x49;
  wire t50    = x49 + invx49;
  wire inv50  = ~t50;
  wire x50    = t50 ^ inv50;
  wire invx50 = ~x50;
  wire t51    = x50 + invx50;
  wire inv51  = ~t51;
  wire x51    = t51 ^ inv51;
  wire invx51 = ~x51;
  wire t52    = x51 + invx51;
  wire inv52  = ~t52;
  wire x52    = t52 ^ inv52;
  wire invx52 = ~x52;
  wire t53    = x52 + invx52;
  wire inv53  = ~t53;
  wire x53    = t53 ^ inv53;
  wire invx53 = ~x53;
  wire t54    = x53 + invx53;
  wire inv54  = ~t54;
  wire x54    = t54 ^ inv54;
  wire invx54 = ~x54;
  wire t55    = x54 + invx54;
  wire inv55  = ~t55;
  wire x55    = t55 ^ inv55;
  wire invx55 = ~x55;
  wire t56    = x55 + invx55;
  wire inv56  = ~t56;
  wire x56    = t56 ^ inv56;
  wire invx56 = ~x56;
  wire t57    = x56 + invx56;
  wire inv57  = ~t57;
  wire x57    = t57 ^ inv57;
  wire invx57 = ~x57;
  wire t58    = x57 + invx57;
  wire inv58  = ~t58;
  wire x58    = t58 ^ inv58;
  wire invx58 = ~x58;
  wire t59    = x58 + invx58;
  wire inv59  = ~t59;
  wire x59    = t59 ^ inv59;
  wire invx59 = ~x59;
  wire t60    = x59 + invx59;
  wire inv60  = ~t60;
  wire x60    = t60 ^ inv60;
  wire invx60 = ~x60;
  wire t61    = x60 + invx60;
  wire inv61  = ~t61;
  wire x61    = t61 ^ inv61;
  wire invx61 = ~x61;
  wire t62    = x61 + invx61;
  wire inv62  = ~t62;
  wire x62    = t62 ^ inv62;
  wire invx62 = ~x62;
  wire t63    = x62 + invx62;
  wire inv63  = ~t63;
  wire x63    = t63 ^ inv63;
  wire invx63 = ~x63;
  wire t64    = x63 + invx63;
  wire inv64  = ~t64;
  wire x64    = t64 ^ inv64;
  wire invx64 = ~x64;
  wire t65    = x64 + invx64;
  wire inv65  = ~t65;
  wire x65    = t65 ^ inv65;
  wire invx65 = ~x65;
  wire t66    = x65 + invx65;
  wire inv66  = ~t66;
  wire x66    = t66 ^ inv66;
  wire invx66 = ~x66;
  wire t67    = x66 + invx66;
  wire inv67  = ~t67;
  wire x67    = t67 ^ inv67;
  wire invx67 = ~x67;
  wire t68    = x67 + invx67;
  wire inv68  = ~t68;
  wire x68    = t68 ^ inv68;
  wire invx68 = ~x68;
  wire t69    = x68 + invx68;
  wire inv69  = ~t69;
  wire x69    = t69 ^ inv69;
  wire invx69 = ~x69;
  wire t70    = x69 + invx69;
  wire inv70  = ~t70;
  wire x70    = t70 ^ inv70;
  wire invx70 = ~x70;
  wire t71    = x70 + invx70;
  wire inv71  = ~t71;
  wire x71    = t71 ^ inv71;
  wire invx71 = ~x71;
  wire t72    = x71 + invx71;
  wire inv72  = ~t72;
  wire x72    = t72 ^ inv72;
  wire invx72 = ~x72;
  wire t73    = x72 + invx72;
  wire inv73  = ~t73;
  wire x73    = t73 ^ inv73;
  wire invx73 = ~x73;
  wire t74    = x73 + invx73;
  wire inv74  = ~t74;
  wire x74    = t74 ^ inv74;
  wire invx74 = ~x74;
  wire t75    = x74 + invx74;
  wire inv75  = ~t75;
  wire x75    = t75 ^ inv75;
  wire invx75 = ~x75;
  wire t76    = x75 + invx75;
  wire inv76  = ~t76;
  wire x76    = t76 ^ inv76;
  wire invx76 = ~x76;
  wire t77    = x76 + invx76;
  wire inv77  = ~t77;
  wire x77    = t77 ^ inv77;
  wire invx77 = ~x77;
  wire t78    = x77 + invx77;
  wire inv78  = ~t78;
  wire x78    = t78 ^ inv78;
  wire invx78 = ~x78;
  wire t79    = x78 + invx78;
  wire inv79  = ~t79;
  wire x79    = t79 ^ inv79;
  wire invx79 = ~x79;
  wire t80    = x79 + invx79;
  wire inv80  = ~t80;
  wire x80    = t80 ^ inv80;
  wire invx80 = ~x80;
  wire t81    = x80 + invx80;
  wire inv81  = ~t81;
  wire x81    = t81 ^ inv81;
  wire invx81 = ~x81;
  wire t82    = x81 + invx81;
  wire inv82  = ~t82;
  wire x82    = t82 ^ inv82;
  wire invx82 = ~x82;
  wire t83    = x82 + invx82;
  wire inv83  = ~t83;
  wire x83    = t83 ^ inv83;
  wire invx83 = ~x83;
  wire t84    = x83 + invx83;
  wire inv84  = ~t84;
  wire x84    = t84 ^ inv84;
  wire invx84 = ~x84;
  wire t85    = x84 + invx84;
  wire inv85  = ~t85;
  wire x85    = t85 ^ inv85;
  wire invx85 = ~x85;
  wire t86    = x85 + invx85;
  wire inv86  = ~t86;
  wire x86    = t86 ^ inv86;
  wire invx86 = ~x86;
  wire t87    = x86 + invx86;
  wire inv87  = ~t87;
  wire x87    = t87 ^ inv87;
  wire invx87 = ~x87;
  wire t88    = x87 + invx87;
  wire inv88  = ~t88;
  wire x88    = t88 ^ inv88;
  wire invx88 = ~x88;
  wire t89    = x88 + invx88;
  wire inv89  = ~t89;
  wire x89    = t89 ^ inv89;
  wire invx89 = ~x89;
  wire t90    = x89 + invx89;
  wire inv90  = ~t90;
  wire x90    = t90 ^ inv90;
  wire invx90 = ~x90;
  wire t91    = x90 + invx90;
  wire inv91  = ~t91;
  wire x91    = t91 ^ inv91;
  wire invx91 = ~x91;
  wire t92    = x91 + invx91;
  wire inv92  = ~t92;
  wire x92    = t92 ^ inv92;
  wire invx92 = ~x92;
  wire t93    = x92 + invx92;
  wire inv93  = ~t93;
  wire x93    = t93 ^ inv93;
  wire invx93 = ~x93;
  wire t94    = x93 + invx93;
  wire inv94  = ~t94;
  wire x94    = t94 ^ inv94;
  wire invx94 = ~x94;
  wire t95    = x94 + invx94;
  wire inv95  = ~t95;
  wire x95    = t95 ^ inv95;
  wire invx95 = ~x95;
  wire t96    = x95 + invx95;
  wire inv96  = ~t96;
  wire x96    = t96 ^ inv96;
  wire invx96 = ~x96;
  wire t97    = x96 + invx96;
  wire inv97  = ~t97;
  wire x97    = t97 ^ inv97;
  wire invx97 = ~x97;
  wire t98    = x97 + invx97;
  wire inv98  = ~t98;
  wire x98    = t98 ^ inv98;
  wire invx98 = ~x98;
  wire t99    = x98 + invx98;
  wire inv99  = ~t99;
  wire x99    = t99 ^ inv99;
  wire invx99 = ~x99;
  wire t100    = x99 + invx99;
  wire inv100  = ~t100;
  wire x100    = t100 ^ inv100;
  wire invx100 = ~x100;
  wire t101    = x100 + invx100;
  wire inv101  = ~t101;
  wire x101    = t101 ^ inv101;
  wire invx101 = ~x101;
  wire t102    = x101 + invx101;
  wire inv102  = ~t102;
  wire x102    = t102 ^ inv102;
  wire invx102 = ~x102;
  wire t103    = x102 + invx102;
  wire inv103  = ~t103;
  wire x103    = t103 ^ inv103;
  wire invx103 = ~x103;
  wire t104    = x103 + invx103;
  wire inv104  = ~t104;
  wire x104    = t104 ^ inv104;
  wire invx104 = ~x104;
  wire t105    = x104 + invx104;
  wire inv105  = ~t105;
  wire x105    = t105 ^ inv105;
  wire invx105 = ~x105;
  wire t106    = x105 + invx105;
  wire inv106  = ~t106;
  wire x106    = t106 ^ inv106;
  wire invx106 = ~x106;
  wire t107    = x106 + invx106;
  wire inv107  = ~t107;
  wire x107    = t107 ^ inv107;
  wire invx107 = ~x107;
  wire t108    = x107 + invx107;
  wire inv108  = ~t108;
  wire x108    = t108 ^ inv108;
  wire invx108 = ~x108;
  wire t109    = x108 + invx108;
  wire inv109  = ~t109;
  wire x109    = t109 ^ inv109;
  wire invx109 = ~x109;
  wire t110    = x109 + invx109;
  wire inv110  = ~t110;
  wire x110    = t110 ^ inv110;
  wire invx110 = ~x110;
  wire t111    = x110 + invx110;
  wire inv111  = ~t111;
  wire x111    = t111 ^ inv111;
  wire invx111 = ~x111;
  wire t112    = x111 + invx111;
  wire inv112  = ~t112;
  wire x112    = t112 ^ inv112;
  wire invx112 = ~x112;
  wire t113    = x112 + invx112;
  wire inv113  = ~t113;
  wire x113    = t113 ^ inv113;
  wire invx113 = ~x113;
  wire t114    = x113 + invx113;
  wire inv114  = ~t114;
  wire x114    = t114 ^ inv114;
  wire invx114 = ~x114;
  wire t115    = x114 + invx114;
  wire inv115  = ~t115;
  wire x115    = t115 ^ inv115;
  wire invx115 = ~x115;
  wire t116    = x115 + invx115;
  wire inv116  = ~t116;
  wire x116    = t116 ^ inv116;
  wire invx116 = ~x116;
  wire t117    = x116 + invx116;
  wire inv117  = ~t117;
  wire x117    = t117 ^ inv117;
  wire invx117 = ~x117;
  wire t118    = x117 + invx117;
  wire inv118  = ~t118;
  wire x118    = t118 ^ inv118;
  wire invx118 = ~x118;
  wire t119    = x118 + invx118;
  wire inv119  = ~t119;
  wire x119    = t119 ^ inv119;
  wire invx119 = ~x119;
  wire t120    = x119 + invx119;
  wire inv120  = ~t120;
  wire x120    = t120 ^ inv120;
  wire invx120 = ~x120;
  wire t121    = x120 + invx120;
  wire inv121  = ~t121;
  wire x121    = t121 ^ inv121;
  wire invx121 = ~x121;
  wire t122    = x121 + invx121;
  wire inv122  = ~t122;
  wire x122    = t122 ^ inv122;
  wire invx122 = ~x122;
  wire t123    = x122 + invx122;
  wire inv123  = ~t123;
  wire x123    = t123 ^ inv123;
  wire invx123 = ~x123;
  wire t124    = x123 + invx123;
  wire inv124  = ~t124;
  wire x124    = t124 ^ inv124;
  wire invx124 = ~x124;
  wire t125    = x124 + invx124;
  wire inv125  = ~t125;
  wire x125    = t125 ^ inv125;
  wire invx125 = ~x125;
  wire t126    = x125 + invx125;
  wire inv126  = ~t126;
  wire x126    = t126 ^ inv126;
  wire invx126 = ~x126;
  wire t127    = x126 + invx126;
  wire inv127  = ~t127;
  wire x127    = t127 ^ inv127;
  wire invx127 = ~x127;
  wire t128    = x127 + invx127;
  wire inv128  = ~t128;
  wire x128    = t128 ^ inv128;
  wire invx128 = ~x128;
  wire t129    = x128 + invx128;
  wire inv129  = ~t129;
  wire x129    = t129 ^ inv129;
  wire invx129 = ~x129;
  wire t130    = x129 + invx129;
  wire inv130  = ~t130;
  wire x130    = t130 ^ inv130;
  wire invx130 = ~x130;
  wire t131    = x130 + invx130;
  wire inv131  = ~t131;
  wire x131    = t131 ^ inv131;
  wire invx131 = ~x131;
  wire t132    = x131 + invx131;
  wire inv132  = ~t132;
  wire x132    = t132 ^ inv132;
  wire invx132 = ~x132;
  wire t133    = x132 + invx132;
  wire inv133  = ~t133;
  wire x133    = t133 ^ inv133;
  wire invx133 = ~x133;
  wire t134    = x133 + invx133;
  wire inv134  = ~t134;
  wire x134    = t134 ^ inv134;
  wire invx134 = ~x134;
  wire t135    = x134 + invx134;
  wire inv135  = ~t135;
  wire x135    = t135 ^ inv135;
  wire invx135 = ~x135;
  wire t136    = x135 + invx135;
  wire inv136  = ~t136;
  wire x136    = t136 ^ inv136;
  wire invx136 = ~x136;
  wire t137    = x136 + invx136;
  wire inv137  = ~t137;
  wire x137    = t137 ^ inv137;
  wire invx137 = ~x137;
  wire t138    = x137 + invx137;
  wire inv138  = ~t138;
  wire x138    = t138 ^ inv138;
  wire invx138 = ~x138;
  wire t139    = x138 + invx138;
  wire inv139  = ~t139;
  wire x139    = t139 ^ inv139;
  wire invx139 = ~x139;
  wire t140    = x139 + invx139;
  wire inv140  = ~t140;
  wire x140    = t140 ^ inv140;
  wire invx140 = ~x140;
  wire t141    = x140 + invx140;
  wire inv141  = ~t141;
  wire x141    = t141 ^ inv141;
  wire invx141 = ~x141;
  wire t142    = x141 + invx141;
  wire inv142  = ~t142;
  wire x142    = t142 ^ inv142;
  wire invx142 = ~x142;
  wire t143    = x142 + invx142;
  wire inv143  = ~t143;
  wire x143    = t143 ^ inv143;
  wire invx143 = ~x143;

  wire SnxnLv1Inst0_z;
  SnxnLv1Inst0 inst_SnxnLv1Inst0(
  .a(a),
  .b(b),
  .z(SnxnLv1Inst0_z)
  );

  wire sum = SnxnLv1Inst0_z;
  assign z = sum ^ a;
endmodule

module SnxnLv1Inst0 (
  input  a,
  input  b,
  output z
);
  wire t0 = a + b;
  wire inv0  = ~t0;
  wire x0    = t0 ^ inv0;
  wire invx0 = ~x0;
  wire t1    = x0 + invx0;
  wire inv1  = ~t1;
  wire x1    = t1 ^ inv1;
  wire invx1 = ~x1;
  wire t2    = x1 + invx1;
  wire inv2  = ~t2;
  wire x2    = t2 ^ inv2;
  wire invx2 = ~x2;
  wire t3    = x2 + invx2;
  wire inv3  = ~t3;
  wire x3    = t3 ^ inv3;
  wire invx3 = ~x3;
  wire t4    = x3 + invx3;
  wire inv4  = ~t4;
  wire x4    = t4 ^ inv4;
  wire invx4 = ~x4;
  wire t5    = x4 + invx4;
  wire inv5  = ~t5;
  wire x5    = t5 ^ inv5;
  wire invx5 = ~x5;
  wire t6    = x5 + invx5;
  wire inv6  = ~t6;
  wire x6    = t6 ^ inv6;
  wire invx6 = ~x6;
  wire t7    = x6 + invx6;
  wire inv7  = ~t7;
  wire x7    = t7 ^ inv7;
  wire invx7 = ~x7;
  wire t8    = x7 + invx7;
  wire inv8  = ~t8;
  wire x8    = t8 ^ inv8;
  wire invx8 = ~x8;
  wire t9    = x8 + invx8;
  wire inv9  = ~t9;
  wire x9    = t9 ^ inv9;
  wire invx9 = ~x9;
  wire t10    = x9 + invx9;
  wire inv10  = ~t10;
  wire x10    = t10 ^ inv10;
  wire invx10 = ~x10;
  wire t11    = x10 + invx10;
  wire inv11  = ~t11;
  wire x11    = t11 ^ inv11;
  wire invx11 = ~x11;
  wire t12    = x11 + invx11;
  wire inv12  = ~t12;
  wire x12    = t12 ^ inv12;
  wire invx12 = ~x12;
  wire t13    = x12 + invx12;
  wire inv13  = ~t13;
  wire x13    = t13 ^ inv13;
  wire invx13 = ~x13;
  wire t14    = x13 + invx13;
  wire inv14  = ~t14;
  wire x14    = t14 ^ inv14;
  wire invx14 = ~x14;
  wire t15    = x14 + invx14;
  wire inv15  = ~t15;
  wire x15    = t15 ^ inv15;
  wire invx15 = ~x15;
  wire t16    = x15 + invx15;
  wire inv16  = ~t16;
  wire x16    = t16 ^ inv16;
  wire invx16 = ~x16;
  wire t17    = x16 + invx16;
  wire inv17  = ~t17;
  wire x17    = t17 ^ inv17;
  wire invx17 = ~x17;
  wire t18    = x17 + invx17;
  wire inv18  = ~t18;
  wire x18    = t18 ^ inv18;
  wire invx18 = ~x18;
  wire t19    = x18 + invx18;
  wire inv19  = ~t19;
  wire x19    = t19 ^ inv19;
  wire invx19 = ~x19;
  wire t20    = x19 + invx19;
  wire inv20  = ~t20;
  wire x20    = t20 ^ inv20;
  wire invx20 = ~x20;
  wire t21    = x20 + invx20;
  wire inv21  = ~t21;
  wire x21    = t21 ^ inv21;
  wire invx21 = ~x21;
  wire t22    = x21 + invx21;
  wire inv22  = ~t22;
  wire x22    = t22 ^ inv22;
  wire invx22 = ~x22;
  wire t23    = x22 + invx22;
  wire inv23  = ~t23;
  wire x23    = t23 ^ inv23;
  wire invx23 = ~x23;
  wire t24    = x23 + invx23;
  wire inv24  = ~t24;
  wire x24    = t24 ^ inv24;
  wire invx24 = ~x24;
  wire t25    = x24 + invx24;
  wire inv25  = ~t25;
  wire x25    = t25 ^ inv25;
  wire invx25 = ~x25;
  wire t26    = x25 + invx25;
  wire inv26  = ~t26;
  wire x26    = t26 ^ inv26;
  wire invx26 = ~x26;
  wire t27    = x26 + invx26;
  wire inv27  = ~t27;
  wire x27    = t27 ^ inv27;
  wire invx27 = ~x27;
  wire t28    = x27 + invx27;
  wire inv28  = ~t28;
  wire x28    = t28 ^ inv28;
  wire invx28 = ~x28;
  wire t29    = x28 + invx28;
  wire inv29  = ~t29;
  wire x29    = t29 ^ inv29;
  wire invx29 = ~x29;
  wire t30    = x29 + invx29;
  wire inv30  = ~t30;
  wire x30    = t30 ^ inv30;
  wire invx30 = ~x30;
  wire t31    = x30 + invx30;
  wire inv31  = ~t31;
  wire x31    = t31 ^ inv31;
  wire invx31 = ~x31;
  wire t32    = x31 + invx31;
  wire inv32  = ~t32;
  wire x32    = t32 ^ inv32;
  wire invx32 = ~x32;
  wire t33    = x32 + invx32;
  wire inv33  = ~t33;
  wire x33    = t33 ^ inv33;
  wire invx33 = ~x33;
  wire t34    = x33 + invx33;
  wire inv34  = ~t34;
  wire x34    = t34 ^ inv34;
  wire invx34 = ~x34;
  wire t35    = x34 + invx34;
  wire inv35  = ~t35;
  wire x35    = t35 ^ inv35;
  wire invx35 = ~x35;
  wire t36    = x35 + invx35;
  wire inv36  = ~t36;
  wire x36    = t36 ^ inv36;
  wire invx36 = ~x36;
  wire t37    = x36 + invx36;
  wire inv37  = ~t37;
  wire x37    = t37 ^ inv37;
  wire invx37 = ~x37;
  wire t38    = x37 + invx37;
  wire inv38  = ~t38;
  wire x38    = t38 ^ inv38;
  wire invx38 = ~x38;
  wire t39    = x38 + invx38;
  wire inv39  = ~t39;
  wire x39    = t39 ^ inv39;
  wire invx39 = ~x39;
  wire t40    = x39 + invx39;
  wire inv40  = ~t40;
  wire x40    = t40 ^ inv40;
  wire invx40 = ~x40;
  wire t41    = x40 + invx40;
  wire inv41  = ~t41;
  wire x41    = t41 ^ inv41;
  wire invx41 = ~x41;
  wire t42    = x41 + invx41;
  wire inv42  = ~t42;
  wire x42    = t42 ^ inv42;
  wire invx42 = ~x42;
  wire t43    = x42 + invx42;
  wire inv43  = ~t43;
  wire x43    = t43 ^ inv43;
  wire invx43 = ~x43;
  wire t44    = x43 + invx43;
  wire inv44  = ~t44;
  wire x44    = t44 ^ inv44;
  wire invx44 = ~x44;
  wire t45    = x44 + invx44;
  wire inv45  = ~t45;
  wire x45    = t45 ^ inv45;
  wire invx45 = ~x45;
  wire t46    = x45 + invx45;
  wire inv46  = ~t46;
  wire x46    = t46 ^ inv46;
  wire invx46 = ~x46;
  wire t47    = x46 + invx46;
  wire inv47  = ~t47;
  wire x47    = t47 ^ inv47;
  wire invx47 = ~x47;
  wire t48    = x47 + invx47;
  wire inv48  = ~t48;
  wire x48    = t48 ^ inv48;
  wire invx48 = ~x48;
  wire t49    = x48 + invx48;
  wire inv49  = ~t49;
  wire x49    = t49 ^ inv49;
  wire invx49 = ~x49;
  wire t50    = x49 + invx49;
  wire inv50  = ~t50;
  wire x50    = t50 ^ inv50;
  wire invx50 = ~x50;
  wire t51    = x50 + invx50;
  wire inv51  = ~t51;
  wire x51    = t51 ^ inv51;
  wire invx51 = ~x51;
  wire t52    = x51 + invx51;
  wire inv52  = ~t52;
  wire x52    = t52 ^ inv52;
  wire invx52 = ~x52;
  wire t53    = x52 + invx52;
  wire inv53  = ~t53;
  wire x53    = t53 ^ inv53;
  wire invx53 = ~x53;
  wire t54    = x53 + invx53;
  wire inv54  = ~t54;
  wire x54    = t54 ^ inv54;
  wire invx54 = ~x54;
  wire t55    = x54 + invx54;
  wire inv55  = ~t55;
  wire x55    = t55 ^ inv55;
  wire invx55 = ~x55;
  wire t56    = x55 + invx55;
  wire inv56  = ~t56;
  wire x56    = t56 ^ inv56;
  wire invx56 = ~x56;
  wire t57    = x56 + invx56;
  wire inv57  = ~t57;
  wire x57    = t57 ^ inv57;
  wire invx57 = ~x57;
  wire t58    = x57 + invx57;
  wire inv58  = ~t58;
  wire x58    = t58 ^ inv58;
  wire invx58 = ~x58;
  wire t59    = x58 + invx58;
  wire inv59  = ~t59;
  wire x59    = t59 ^ inv59;
  wire invx59 = ~x59;
  wire t60    = x59 + invx59;
  wire inv60  = ~t60;
  wire x60    = t60 ^ inv60;
  wire invx60 = ~x60;
  wire t61    = x60 + invx60;
  wire inv61  = ~t61;
  wire x61    = t61 ^ inv61;
  wire invx61 = ~x61;
  wire t62    = x61 + invx61;
  wire inv62  = ~t62;
  wire x62    = t62 ^ inv62;
  wire invx62 = ~x62;
  wire t63    = x62 + invx62;
  wire inv63  = ~t63;
  wire x63    = t63 ^ inv63;
  wire invx63 = ~x63;
  wire t64    = x63 + invx63;
  wire inv64  = ~t64;
  wire x64    = t64 ^ inv64;
  wire invx64 = ~x64;
  wire t65    = x64 + invx64;
  wire inv65  = ~t65;
  wire x65    = t65 ^ inv65;
  wire invx65 = ~x65;
  wire t66    = x65 + invx65;
  wire inv66  = ~t66;
  wire x66    = t66 ^ inv66;
  wire invx66 = ~x66;
  wire t67    = x66 + invx66;
  wire inv67  = ~t67;
  wire x67    = t67 ^ inv67;
  wire invx67 = ~x67;
  wire t68    = x67 + invx67;
  wire inv68  = ~t68;
  wire x68    = t68 ^ inv68;
  wire invx68 = ~x68;
  wire t69    = x68 + invx68;
  wire inv69  = ~t69;
  wire x69    = t69 ^ inv69;
  wire invx69 = ~x69;
  wire t70    = x69 + invx69;
  wire inv70  = ~t70;
  wire x70    = t70 ^ inv70;
  wire invx70 = ~x70;
  wire t71    = x70 + invx70;
  wire inv71  = ~t71;
  wire x71    = t71 ^ inv71;
  wire invx71 = ~x71;
  wire t72    = x71 + invx71;
  wire inv72  = ~t72;
  wire x72    = t72 ^ inv72;
  wire invx72 = ~x72;
  wire t73    = x72 + invx72;
  wire inv73  = ~t73;
  wire x73    = t73 ^ inv73;
  wire invx73 = ~x73;
  wire t74    = x73 + invx73;
  wire inv74  = ~t74;
  wire x74    = t74 ^ inv74;
  wire invx74 = ~x74;
  wire t75    = x74 + invx74;
  wire inv75  = ~t75;
  wire x75    = t75 ^ inv75;
  wire invx75 = ~x75;
  wire t76    = x75 + invx75;
  wire inv76  = ~t76;
  wire x76    = t76 ^ inv76;
  wire invx76 = ~x76;
  wire t77    = x76 + invx76;
  wire inv77  = ~t77;
  wire x77    = t77 ^ inv77;
  wire invx77 = ~x77;
  wire t78    = x77 + invx77;
  wire inv78  = ~t78;
  wire x78    = t78 ^ inv78;
  wire invx78 = ~x78;
  wire t79    = x78 + invx78;
  wire inv79  = ~t79;
  wire x79    = t79 ^ inv79;
  wire invx79 = ~x79;
  wire t80    = x79 + invx79;
  wire inv80  = ~t80;
  wire x80    = t80 ^ inv80;
  wire invx80 = ~x80;
  wire t81    = x80 + invx80;
  wire inv81  = ~t81;
  wire x81    = t81 ^ inv81;
  wire invx81 = ~x81;
  wire t82    = x81 + invx81;
  wire inv82  = ~t82;
  wire x82    = t82 ^ inv82;
  wire invx82 = ~x82;
  wire t83    = x82 + invx82;
  wire inv83  = ~t83;
  wire x83    = t83 ^ inv83;
  wire invx83 = ~x83;
  wire t84    = x83 + invx83;
  wire inv84  = ~t84;
  wire x84    = t84 ^ inv84;
  wire invx84 = ~x84;
  wire t85    = x84 + invx84;
  wire inv85  = ~t85;
  wire x85    = t85 ^ inv85;
  wire invx85 = ~x85;
  wire t86    = x85 + invx85;
  wire inv86  = ~t86;
  wire x86    = t86 ^ inv86;
  wire invx86 = ~x86;
  wire t87    = x86 + invx86;
  wire inv87  = ~t87;
  wire x87    = t87 ^ inv87;
  wire invx87 = ~x87;
  wire t88    = x87 + invx87;
  wire inv88  = ~t88;
  wire x88    = t88 ^ inv88;
  wire invx88 = ~x88;
  wire t89    = x88 + invx88;
  wire inv89  = ~t89;
  wire x89    = t89 ^ inv89;
  wire invx89 = ~x89;
  wire t90    = x89 + invx89;
  wire inv90  = ~t90;
  wire x90    = t90 ^ inv90;
  wire invx90 = ~x90;
  wire t91    = x90 + invx90;
  wire inv91  = ~t91;
  wire x91    = t91 ^ inv91;
  wire invx91 = ~x91;
  wire t92    = x91 + invx91;
  wire inv92  = ~t92;
  wire x92    = t92 ^ inv92;
  wire invx92 = ~x92;
  wire t93    = x92 + invx92;
  wire inv93  = ~t93;
  wire x93    = t93 ^ inv93;
  wire invx93 = ~x93;
  wire t94    = x93 + invx93;
  wire inv94  = ~t94;
  wire x94    = t94 ^ inv94;
  wire invx94 = ~x94;
  wire t95    = x94 + invx94;
  wire inv95  = ~t95;
  wire x95    = t95 ^ inv95;
  wire invx95 = ~x95;
  wire t96    = x95 + invx95;
  wire inv96  = ~t96;
  wire x96    = t96 ^ inv96;
  wire invx96 = ~x96;
  wire t97    = x96 + invx96;
  wire inv97  = ~t97;
  wire x97    = t97 ^ inv97;
  wire invx97 = ~x97;
  wire t98    = x97 + invx97;
  wire inv98  = ~t98;
  wire x98    = t98 ^ inv98;
  wire invx98 = ~x98;
  wire t99    = x98 + invx98;
  wire inv99  = ~t99;
  wire x99    = t99 ^ inv99;
  wire invx99 = ~x99;
  wire t100    = x99 + invx99;
  wire inv100  = ~t100;
  wire x100    = t100 ^ inv100;
  wire invx100 = ~x100;
  wire t101    = x100 + invx100;
  wire inv101  = ~t101;
  wire x101    = t101 ^ inv101;
  wire invx101 = ~x101;
  wire t102    = x101 + invx101;
  wire inv102  = ~t102;
  wire x102    = t102 ^ inv102;
  wire invx102 = ~x102;
  wire t103    = x102 + invx102;
  wire inv103  = ~t103;
  wire x103    = t103 ^ inv103;
  wire invx103 = ~x103;
  wire t104    = x103 + invx103;
  wire inv104  = ~t104;
  wire x104    = t104 ^ inv104;
  wire invx104 = ~x104;
  wire t105    = x104 + invx104;
  wire inv105  = ~t105;
  wire x105    = t105 ^ inv105;
  wire invx105 = ~x105;
  wire t106    = x105 + invx105;
  wire inv106  = ~t106;
  wire x106    = t106 ^ inv106;
  wire invx106 = ~x106;
  wire t107    = x106 + invx106;
  wire inv107  = ~t107;
  wire x107    = t107 ^ inv107;
  wire invx107 = ~x107;
  wire t108    = x107 + invx107;
  wire inv108  = ~t108;
  wire x108    = t108 ^ inv108;
  wire invx108 = ~x108;
  wire t109    = x108 + invx108;
  wire inv109  = ~t109;
  wire x109    = t109 ^ inv109;
  wire invx109 = ~x109;
  wire t110    = x109 + invx109;
  wire inv110  = ~t110;
  wire x110    = t110 ^ inv110;
  wire invx110 = ~x110;
  wire t111    = x110 + invx110;
  wire inv111  = ~t111;
  wire x111    = t111 ^ inv111;
  wire invx111 = ~x111;
  wire t112    = x111 + invx111;
  wire inv112  = ~t112;
  wire x112    = t112 ^ inv112;
  wire invx112 = ~x112;
  wire t113    = x112 + invx112;
  wire inv113  = ~t113;
  wire x113    = t113 ^ inv113;
  wire invx113 = ~x113;
  wire t114    = x113 + invx113;
  wire inv114  = ~t114;
  wire x114    = t114 ^ inv114;
  wire invx114 = ~x114;
  wire t115    = x114 + invx114;
  wire inv115  = ~t115;
  wire x115    = t115 ^ inv115;
  wire invx115 = ~x115;
  wire t116    = x115 + invx115;
  wire inv116  = ~t116;
  wire x116    = t116 ^ inv116;
  wire invx116 = ~x116;
  wire t117    = x116 + invx116;
  wire inv117  = ~t117;
  wire x117    = t117 ^ inv117;
  wire invx117 = ~x117;
  wire t118    = x117 + invx117;
  wire inv118  = ~t118;
  wire x118    = t118 ^ inv118;
  wire invx118 = ~x118;
  wire t119    = x118 + invx118;
  wire inv119  = ~t119;
  wire x119    = t119 ^ inv119;
  wire invx119 = ~x119;
  wire t120    = x119 + invx119;
  wire inv120  = ~t120;
  wire x120    = t120 ^ inv120;
  wire invx120 = ~x120;
  wire t121    = x120 + invx120;
  wire inv121  = ~t121;
  wire x121    = t121 ^ inv121;
  wire invx121 = ~x121;
  wire t122    = x121 + invx121;
  wire inv122  = ~t122;
  wire x122    = t122 ^ inv122;
  wire invx122 = ~x122;
  wire t123    = x122 + invx122;
  wire inv123  = ~t123;
  wire x123    = t123 ^ inv123;
  wire invx123 = ~x123;
  wire t124    = x123 + invx123;
  wire inv124  = ~t124;
  wire x124    = t124 ^ inv124;
  wire invx124 = ~x124;
  wire t125    = x124 + invx124;
  wire inv125  = ~t125;
  wire x125    = t125 ^ inv125;
  wire invx125 = ~x125;
  wire t126    = x125 + invx125;
  wire inv126  = ~t126;
  wire x126    = t126 ^ inv126;
  wire invx126 = ~x126;
  wire t127    = x126 + invx126;
  wire inv127  = ~t127;
  wire x127    = t127 ^ inv127;
  wire invx127 = ~x127;
  wire t128    = x127 + invx127;
  wire inv128  = ~t128;
  wire x128    = t128 ^ inv128;
  wire invx128 = ~x128;
  wire t129    = x128 + invx128;
  wire inv129  = ~t129;
  wire x129    = t129 ^ inv129;
  wire invx129 = ~x129;
  wire t130    = x129 + invx129;
  wire inv130  = ~t130;
  wire x130    = t130 ^ inv130;
  wire invx130 = ~x130;
  wire t131    = x130 + invx130;
  wire inv131  = ~t131;
  wire x131    = t131 ^ inv131;
  wire invx131 = ~x131;
  wire t132    = x131 + invx131;
  wire inv132  = ~t132;
  wire x132    = t132 ^ inv132;
  wire invx132 = ~x132;
  wire t133    = x132 + invx132;
  wire inv133  = ~t133;
  wire x133    = t133 ^ inv133;
  wire invx133 = ~x133;
  wire t134    = x133 + invx133;
  wire inv134  = ~t134;
  wire x134    = t134 ^ inv134;
  wire invx134 = ~x134;
  wire t135    = x134 + invx134;
  wire inv135  = ~t135;
  wire x135    = t135 ^ inv135;
  wire invx135 = ~x135;
  wire t136    = x135 + invx135;
  wire inv136  = ~t136;
  wire x136    = t136 ^ inv136;
  wire invx136 = ~x136;

  assign z = invx136;
endmodule

